`define DEFINES_DONE
`define EXPONENT 5
`define MANTISSA 10
`define SIGN 1
`define DATAWIDTH (`SIGN+`EXPONENT+`MANTISSA)
`define IEEE_COMPLIANCE 1
`define NUM 8
`define ADDRSIZE 7
`define ADDRSIZE_FOR_TB 10
`define EXPONENT 5
`define MANTISSA 10
`define ACTUAL_MANTISSA 11
`define EXPONENT_LSB 10
`define EXPONENT_MSB 14
`define MANTISSA_LSB 0
`define MANTISSA_MSB 9
`define MANTISSA_MUL_SPLIT_LSB 3
`define MANTISSA_MUL_SPLIT_MSB 9
`define SIGN 1
`define SIGN_LOC 15
`define DWIDTH (`SIGN+`EXPONENT+`MANTISSA)
`define IEEE_COMPLIANCE 1
`define EXPONENT 5
`define MANTISSA 10
`define ACTUAL_MANTISSA 11
`define EXPONENT_LSB 10
`define EXPONENT_MSB 14
`define MANTISSA_LSB 0
`define MANTISSA_MSB 9
`define MANTISSA_MUL_SPLIT_LSB 3
`define MANTISSA_MUL_SPLIT_MSB 9
`define SIGN 1
`define SIGN_LOC 15
`define DWIDTH (`SIGN+`EXPONENT+`MANTISSA)
`define IEEE_COMPLIANCE 1
`define EXPONENT 5
`define MANTISSA 10
`define ACTUAL_MANTISSA 11
`define EXPONENT_LSB 10
`define EXPONENT_MSB 14
`define MANTISSA_LSB 0
`define MANTISSA_MSB 9
`define MANTISSA_MUL_SPLIT_LSB 3
`define MANTISSA_MUL_SPLIT_MSB 9
`define SIGN 1
`define SIGN_LOC 15
`define DWIDTH (`SIGN+`EXPONENT+`MANTISSA)
`define IEEE_COMPLIANCE 1

module LUT2(addr, log);
    input [5:0] addr;
    output reg [15:0] log;

    always @(addr) begin
        case (addr)
			6'b0 		: log = 16'b0000000000000000;
			6'b1 		: log = 16'b0010001111110000;
			6'b10 		: log = 16'b0010011111100001;
			6'b11 		: log = 16'b0010100111011101;
			6'b100 		: log = 16'b0010101111000011;
			6'b101 		: log = 16'b0010110011010000;
			6'b110 		: log = 16'b0010110110111100;
			6'b111 		: log = 16'b0010111010100101;
			6'b1000 		: log = 16'b0010111110001010;
			6'b1001 		: log = 16'b0011000000110110;
			6'b1010 		: log = 16'b0011000010100101;
			6'b1011 		: log = 16'b0011000100010011;
			6'b1100 		: log = 16'b0011000110000000;
			6'b1101 		: log = 16'b0011000111101011;
			6'b1110 		: log = 16'b0011001001010101;
			6'b1111 		: log = 16'b0011001010111101;
			6'b10000 		: log = 16'b0011001100100100;
			6'b10001 		: log = 16'b0011001110001010;
			6'b10010 		: log = 16'b0011001111101110;
			6'b10011 		: log = 16'b0011010000101001;
			6'b10100 		: log = 16'b0011010001011010;
			6'b10101 		: log = 16'b0011010010001010;
			6'b10110 		: log = 16'b0011010010111010;
			6'b10111 		: log = 16'b0011010011101010;
			6'b11000 		: log = 16'b0011010100011000;
			6'b11001 		: log = 16'b0011010101000111;
			6'b11010 		: log = 16'b0011010101110100;
			6'b11011 		: log = 16'b0011010110100010;
			6'b11100 		: log = 16'b0011010111001110;
			6'b11101 		: log = 16'b0011010111111011;
			6'b11110 		: log = 16'b0011011000100111;
			6'b11111 		: log = 16'b0011011001010010;
			6'b100000 		: log = 16'b0011011001111101;
			6'b100001 		: log = 16'b0011011010100111;
			6'b100010 		: log = 16'b0011011011010001;
			6'b100011 		: log = 16'b0011011011111011;
			6'b100100 		: log = 16'b0011011100100100;
			6'b100101 		: log = 16'b0011011101001101;
			6'b100110 		: log = 16'b0011011101110101;
			6'b100111 		: log = 16'b0011011110011101;
			6'b101000 		: log = 16'b0011011111000101;
			6'b101001 		: log = 16'b0011011111101100;
			6'b101010 		: log = 16'b0011100000001001;
			6'b101011 		: log = 16'b0011100000011101;
			6'b101100 		: log = 16'b0011100000110000;
			6'b101101 		: log = 16'b0011100001000010;
			6'b101110 		: log = 16'b0011100001010101;
			6'b101111 		: log = 16'b0011100001101000;
			6'b110000 		: log = 16'b0011100001111010;
			6'b110001 		: log = 16'b0011100010001100;
			6'b110010 		: log = 16'b0011100010011110;
			6'b110011 		: log = 16'b0011100010110000;
			6'b110100 		: log = 16'b0011100011000010;
			6'b110101 		: log = 16'b0011100011010100;
			6'b110110 		: log = 16'b0011100011100101;
			6'b110111 		: log = 16'b0011100011110110;
			6'b111000 		: log = 16'b0011100100000111;
			6'b111001 		: log = 16'b0011100100011000;
			6'b111010 		: log = 16'b0011100100101001;
			6'b111011 		: log = 16'b0011100100111010;
			6'b111100 		: log = 16'b0011100101001011;
			6'b111101 		: log = 16'b0011100101011011;
			6'b111110 		: log = 16'b0011100101101011;
			6'b111111 		: log = 16'b0011100101111100;
        endcase
    end
endmodule
