`define INPUT_WIDTH 32
`define INPUT_WIDTH 32
`define INPUT_WIDTH 32
`define INPUT_WIDTH 32
`define INPUT_WIDTH 32
`define INPUT_WIDTH 32
`define INPUT_WIDTH 32
`define INPUT_WIDTH 32

module cosine_lut (quad, enable, degrees, data, rst, clk);

input [1:0] quad;
input enable;
input rst;
input [`INPUT_WIDTH-1:0] degrees ;
input clk;

//////////////inputs/////////////////

output reg [63:0] data;

//////////////output/////////////////


always@(posedge clk )

//needs to be positive in first and fourth quadrants

 begin
        if (quad == 2'b01 || quad == 2'b10)
        begin
        data[63] <= 1'b1;
        end

        else
        begin
        data[63] <= 1'b0;
        end

	if(enable)
	case (degrees)

//look up table
 
`INPUT_WIDTH'd0  : data[62:0] <= 64'h3ff0000000000000;
`INPUT_WIDTH'd1  : data[62:0] <= 64'h3feffec097f5af8a;
`INPUT_WIDTH'd2  : data[62:0] <= 64'h3feffb0278bf0567;
`INPUT_WIDTH'd3  : data[62:0] <= 64'h3feff4c5ed12e61d;
`INPUT_WIDTH'd4  : data[62:0] <= 64'h3fefec0b7170fff6;
`INPUT_WIDTH'd5  : data[62:0] <= 64'h3fefe0d3b41815a2;
`INPUT_WIDTH'd6  : data[62:0] <= 64'h3fefd31f94f867c6;
`INPUT_WIDTH'd7  : data[62:0] <= 64'h3fefc2f025a23e8b;
`INPUT_WIDTH'd8  : data[62:0] <= 64'h3fefb046a930947a;
`INPUT_WIDTH'd9  : data[62:0] <= 64'h3fef9b24942fe45c;
`INPUT_WIDTH'd10 : data[62:0] <= 64'h3fef838b8c811c17;
`INPUT_WIDTH'd11 : data[62:0] <= 64'h3fef697d6938b6c2;
`INPUT_WIDTH'd12 : data[62:0] <= 64'h3fef4cfc327a0080;
`INPUT_WIDTH'd13 : data[62:0] <= 64'h3fef2e0a214e870f;
`INPUT_WIDTH'd14 : data[62:0] <= 64'h3fef0ca99f79ba25;
`INPUT_WIDTH'd15 : data[62:0] <= 64'h3feee8dd4748bf15;
`INPUT_WIDTH'd16 : data[62:0] <= 64'h3feec2a7e35e7b80;
`INPUT_WIDTH'd17 : data[62:0] <= 64'h3fee9a0c6e7bdb20;
`INPUT_WIDTH'd18 : data[62:0] <= 64'h3fee6f0e134454ff;
`INPUT_WIDTH'd19 : data[62:0] <= 64'h3fee41b02bfeb4cb;
`INPUT_WIDTH'd20 : data[62:0] <= 64'h3fee11f642522d1c;
`INPUT_WIDTH'd21 : data[62:0] <= 64'h3feddfe40effb805;
`INPUT_WIDTH'd22 : data[62:0] <= 64'h3fedab7d7997cb58;
`INPUT_WIDTH'd23 : data[62:0] <= 64'h3fed74c6982c666f;
`INPUT_WIDTH'd24 : data[62:0] <= 64'h3fed3bc3aeff7f95;
`INPUT_WIDTH'd25 : data[62:0] <= 64'h3fed0079302dd767;
`INPUT_WIDTH'd26 : data[62:0] <= 64'h3fecc2ebbb5638ca;
`INPUT_WIDTH'd27 : data[62:0] <= 64'h3fec83201d3d2c6d;
`INPUT_WIDTH'd28 : data[62:0] <= 64'h3fec411b4f6d2708;
`INPUT_WIDTH'd29 : data[62:0] <= 64'h3febfce277d339c6;
`INPUT_WIDTH'd30 : data[62:0] <= 64'h3febb67ae8584cab;
`INPUT_WIDTH'd31 : data[62:0] <= 64'h3feb6dea1e76eade;
`INPUT_WIDTH'd32 : data[62:0] <= 64'h3feb2335c2cda945;
`INPUT_WIDTH'd33 : data[62:0] <= 64'h3fead663a8ae2fdc;
`INPUT_WIDTH'd34 : data[62:0] <= 64'h3fea8779cda8eea5;
`INPUT_WIDTH'd35 : data[62:0] <= 64'h3fea367e59158747;
`INPUT_WIDTH'd36 : data[62:0] <= 64'h3fe9e3779b97f4a8;
`INPUT_WIDTH'd37 : data[62:0] <= 64'h3fe98e6c0ea27a14;
`INPUT_WIDTH'd38 : data[62:0] <= 64'h3fe9376253f463d1;
`INPUT_WIDTH'd39 : data[62:0] <= 64'h3fe8de613515a328;
`INPUT_WIDTH'd40 : data[62:0] <= 64'h3fe8836fa2cf5039;
`INPUT_WIDTH'd41 : data[62:0] <= 64'h3fe82694b4a11c37;
`INPUT_WIDTH'd42 : data[62:0] <= 64'h3fe7c7d7a833bec2;
`INPUT_WIDTH'd43 : data[62:0] <= 64'h3fe7673fe0c86982;
`INPUT_WIDTH'd44 : data[62:0] <= 64'h3fe704d4e6a54d39;
`INPUT_WIDTH'd45 : data[62:0] <= 64'h3fe6a09e667f3bcd;
`INPUT_WIDTH'd46 : data[62:0] <= 64'h3fe63aa430e07311;
`INPUT_WIDTH'd47 : data[62:0] <= 64'h3fe5d2ee398c9c2b;
`INPUT_WIDTH'd48 : data[62:0] <= 64'h3fe5698496e20bd8;
`INPUT_WIDTH'd49 : data[62:0] <= 64'h3fe4fe6f81384fd5;
`INPUT_WIDTH'd50 : data[62:0] <= 64'h3fe491b7523c161d;
`INPUT_WIDTH'd51 : data[62:0] <= 64'h3fe4236484487abe;
`INPUT_WIDTH'd52 : data[62:0] <= 64'h3fe3b37fb1bdc939;
`INPUT_WIDTH'd53 : data[62:0] <= 64'h3fe342119455beb7;
`INPUT_WIDTH'd54 : data[62:0] <= 64'h3fe2cf2304755a5e;
`INPUT_WIDTH'd55 : data[62:0] <= 64'h3fe25abcf87c4979;
`INPUT_WIDTH'd56 : data[62:0] <= 64'h3fe1e4e88411fd12;
`INPUT_WIDTH'd57 : data[62:0] <= 64'h3fe16daed770771e;
`INPUT_WIDTH'd58 : data[62:0] <= 64'h3fe0f5193eacdd2a;
`INPUT_WIDTH'd59 : data[62:0] <= 64'h3fe07b3120fddf15;
`INPUT_WIDTH'd60 : data[62:0] <= 64'h3fe0000000000001;
`INPUT_WIDTH'd61 : data[62:0] <= 64'h3fdf071eedefa0ee;
`INPUT_WIDTH'd62 : data[62:0] <= 64'h3fde0bd27424507a;
`INPUT_WIDTH'd63 : data[62:0] <= 64'h3fdd0e2e2b44de01;
`INPUT_WIDTH'd64 : data[62:0] <= 64'h3fdc0e45dabe05c9;
`INPUT_WIDTH'd65 : data[62:0] <= 64'h3fdb0c2d77379853;
`INPUT_WIDTH'd66 : data[62:0] <= 64'h3fda07f921061ad4;
`INPUT_WIDTH'd67 : data[62:0] <= 64'h3fd901bd2298ffaa;
`INPUT_WIDTH'd68 : data[62:0] <= 64'h3fd7f98deee59684;
`INPUT_WIDTH'd69 : data[62:0] <= 64'h3fd6ef801fced33a;
`INPUT_WIDTH'd70 : data[62:0] <= 64'h3fd5e3a8748a0bf7;
`INPUT_WIDTH'd71 : data[62:0] <= 64'h3fd4d61bd000cddd;
`INPUT_WIDTH'd72 : data[62:0] <= 64'h3fd3c6ef372fe950;
`INPUT_WIDTH'd73 : data[62:0] <= 64'h3fd2b637cf83d5c8;
`INPUT_WIDTH'd74 : data[62:0] <= 64'h3fd1a40add328e29;
`INPUT_WIDTH'd75 : data[62:0] <= 64'h3fd0907dc1930690;
`INPUT_WIDTH'd76 : data[62:0] <= 64'h3fcef74bf2e4b91b;
`INPUT_WIDTH'd77 : data[62:0] <= 64'h3fcccb3236cdc67a;
`INPUT_WIDTH'd78 : data[62:0] <= 64'h3fca9cd9ac4258f2;
`INPUT_WIDTH'd79 : data[62:0] <= 64'h3fc86c6ddd766253;
`INPUT_WIDTH'd80 : data[62:0] <= 64'h3fc63a1a7e0b738c;
`INPUT_WIDTH'd81 : data[62:0] <= 64'h3fc4060b67a85377;
`INPUT_WIDTH'd82 : data[62:0] <= 64'h3fc1d06c968d9e1a;
`INPUT_WIDTH'd83 : data[62:0] <= 64'h3fbf32d44c4f62d4;
`INPUT_WIDTH'd84 : data[62:0] <= 64'h3fbac2609b3c576b;
`INPUT_WIDTH'd85 : data[62:0] <= 64'h3fb64fd6b8c28110;
`INPUT_WIDTH'd86 : data[62:0] <= 64'h3fb1db8f6d6a5123;
`INPUT_WIDTH'd87 : data[62:0] <= 64'h3faacbc748efc921;
`INPUT_WIDTH'd88 : data[62:0] <= 64'h3fa1de58c9f7dc37;
`INPUT_WIDTH'd89 : data[62:0] <= 64'h3f91df0b2b89dd37;
`INPUT_WIDTH'd90 : data[62:0] <= 64'h0000000000000000;

default:data <= 64'h0;

endcase

else 
  data <= 64'hxxxxxxxxxxxxxxx;




end

endmodule
