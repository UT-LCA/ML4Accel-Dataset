`define M     593         // M is the degree of the irreducible polynomial
`define WIDTH (2*`M-1)    // width for a GF(3^M) element
`define WIDTH_D0 1187
`define M     593         // M is the degree of the irreducible polynomial
`define WIDTH (2*`M-1)    // width for a GF(3^M) element
`define WIDTH_D0 1187
`define M     593         // M is the degree of the irreducible polynomial
`define WIDTH (2*`M-1)    // width for a GF(3^M) element
`define WIDTH_D0 1187
`define M     593         // M is the degree of the irreducible polynomial
`define WIDTH (2*`M-1)    // width for a GF(3^M) element
`define WIDTH_D0 1187
`define M     593         // M is the degree of the irreducible polynomial
`define WIDTH (2*`M-1)    // width for a GF(3^M) element
`define WIDTH_D0 1187

module v2(a, c);
    input [1185:0] a;
    output [1185:0] c;
    assign c[1:0] = 0;
    assign c[3:2] = 0;
    assign c[5:4] = 0;
    assign c[7:6] = 0;
    assign c[9:8] = 0;
    assign c[11:10] = 0;
    assign c[13:12] = 0;
    assign c[15:14] = 0;
    assign c[17:16] = 0;
    assign c[19:18] = 0;
    assign c[21:20] = 0;
    assign c[23:22] = 0;
    assign c[25:24] = 0;
    assign c[27:26] = 0;
    assign c[29:28] = 0;
    assign c[31:30] = 0;
    assign c[33:32] = 0;
    assign c[35:34] = 0;
    assign c[37:36] = 0;
    assign c[39:38] = 0;
    assign c[41:40] = 0;
    assign c[43:42] = 0;
    assign c[45:44] = 0;
    assign c[47:46] = 0;
    assign c[49:48] = 0;
    assign c[51:50] = 0;
    assign c[53:52] = 0;
    assign c[55:54] = 0;
    assign c[57:56] = 0;
    assign c[59:58] = 0;
    assign c[61:60] = 0;
    assign c[63:62] = 0;
    assign c[65:64] = 0;
    assign c[67:66] = 0;
    assign c[69:68] = 0;
    assign c[71:70] = 0;
    assign c[73:72] = 0;
    assign c[75:74] = 0;
    assign c[77:76] = 0;
    assign c[79:78] = 0;
    assign c[81:80] = 0;
    assign c[83:82] = 0;
    assign c[85:84] = 0;
    assign c[87:86] = 0;
    assign c[89:88] = 0;
    assign c[91:90] = 0;
    assign c[93:92] = 0;
    assign c[95:94] = 0;
    assign c[97:96] = 0;
    assign c[99:98] = 0;
    assign c[101:100] = 0;
    assign c[103:102] = 0;
    assign c[105:104] = 0;
    assign c[107:106] = 0;
    assign c[109:108] = 0;
    assign c[111:110] = 0;
    assign c[113:112] = 0;
    assign c[115:114] = 0;
    assign c[117:116] = 0;
    assign c[119:118] = 0;
    assign c[121:120] = 0;
    assign c[123:122] = 0;
    assign c[125:124] = 0;
    assign c[127:126] = 0;
    assign c[129:128] = 0;
    assign c[131:130] = 0;
    assign c[133:132] = 0;
    assign c[135:134] = 0;
    assign c[137:136] = 0;
    assign c[139:138] = 0;
    assign c[141:140] = 0;
    assign c[143:142] = 0;
    assign c[145:144] = 0;
    assign c[147:146] = 0;
    assign c[149:148] = 0;
    assign c[151:150] = 0;
    assign c[153:152] = 0;
    assign c[155:154] = 0;
    assign c[157:156] = 0;
    assign c[159:158] = 0;
    assign c[161:160] = 0;
    assign c[163:162] = 0;
    assign c[165:164] = 0;
    assign c[167:166] = 0;
    assign c[169:168] = 0;
    assign c[171:170] = 0;
    assign c[173:172] = 0;
    assign c[175:174] = 0;
    assign c[177:176] = 0;
    assign c[179:178] = 0;
    assign c[181:180] = 0;
    assign c[183:182] = 0;
    assign c[185:184] = 0;
    assign c[187:186] = 0;
    assign c[189:188] = 0;
    assign c[191:190] = 0;
    assign c[193:192] = 0;
    assign c[195:194] = 0;
    assign c[197:196] = 0;
    assign c[199:198] = 0;
    assign c[201:200] = 0;
    assign c[203:202] = 0;
    assign c[205:204] = 0;
    assign c[207:206] = 0;
    assign c[209:208] = 0;
    assign c[211:210] = 0;
    assign c[213:212] = 0;
    assign c[215:214] = 0;
    assign c[217:216] = 0;
    assign c[219:218] = 0;
    assign c[221:220] = 0;
    assign c[223:222] = 0;
    assign c[225:224] = 0;
    assign c[227:226] = 0;
    assign c[229:228] = {a[1038], a[1039]};
    assign c[231:230] = 0;
    assign c[233:232] = 0;
    assign c[235:234] = a[79:78];
    assign c[237:236] = 0;
    assign c[239:238] = 0;
    assign c[241:240] = a[797:796];
    assign c[243:242] = 0;
    assign c[245:244] = 0;
    assign c[247:246] = a[799:798];
    assign c[249:248] = 0;
    assign c[251:250] = 0;
    assign c[253:252] = {a[1046], a[1047]};
    assign c[255:254] = 0;
    assign c[257:256] = 0;
    assign c[259:258] = {a[1048], a[1049]};
    assign c[261:260] = 0;
    assign c[263:262] = 0;
    assign c[265:264] = {a[1050], a[1051]};
    assign c[267:266] = 0;
    assign c[269:268] = 0;
    assign c[271:270] = {a[1052], a[1053]};
    assign c[273:272] = 0;
    assign c[275:274] = 0;
    assign c[277:276] = {a[1054], a[1055]};
    assign c[279:278] = 0;
    assign c[281:280] = 0;
    assign c[283:282] = a[95:94];
    assign c[285:284] = 0;
    assign c[287:286] = 0;
    assign c[289:288] = a[813:812];
    assign c[291:290] = 0;
    assign c[293:292] = 0;
    assign c[295:294] = a[815:814];
    assign c[297:296] = 0;
    assign c[299:298] = 0;
    assign c[301:300] = {a[1062], a[1063]};
    assign c[303:302] = 0;
    assign c[305:304] = 0;
    assign c[307:306] = {a[1064], a[1065]};
    assign c[309:308] = 0;
    assign c[311:310] = 0;
    assign c[313:312] = {a[1066], a[1067]};
    assign c[315:314] = 0;
    assign c[317:316] = 0;
    assign c[319:318] = {a[1068], a[1069]};
    assign c[321:320] = 0;
    assign c[323:322] = 0;
    assign c[325:324] = {a[1070], a[1071]};
    assign c[327:326] = 0;
    assign c[329:328] = 0;
    assign c[331:330] = a[111:110];
    assign c[333:332] = 0;
    assign c[335:334] = 0;
    assign c[337:336] = a[829:828];
    assign c[339:338] = 0;
    assign c[341:340] = 0;
    assign c[343:342] = a[831:830];
    assign c[345:344] = 0;
    assign c[347:346] = 0;
    assign c[349:348] = {a[1078], a[1079]};
    assign c[351:350] = 0;
    assign c[353:352] = 0;
    assign c[355:354] = {a[1080], a[1081]};
    assign c[357:356] = 0;
    assign c[359:358] = 0;
    assign c[361:360] = {a[1082], a[1083]};
    assign c[363:362] = 0;
    assign c[365:364] = 0;
    assign c[367:366] = {a[1084], a[1085]};
    assign c[369:368] = 0;
    assign c[371:370] = 0;
    assign c[373:372] = {a[1086], a[1087]};
    assign c[375:374] = 0;
    assign c[377:376] = 0;
    assign c[379:378] = a[127:126];
    assign c[381:380] = 0;
    assign c[383:382] = 0;
    assign c[385:384] = a[845:844];
    assign c[387:386] = 0;
    assign c[389:388] = 0;
    assign c[391:390] = a[847:846];
    assign c[393:392] = 0;
    assign c[395:394] = 0;
    assign c[397:396] = {a[1094], a[1095]};
    assign c[399:398] = 0;
    assign c[401:400] = 0;
    assign c[403:402] = {a[1096], a[1097]};
    assign c[405:404] = 0;
    assign c[407:406] = 0;
    assign c[409:408] = {a[1098], a[1099]};
    assign c[411:410] = 0;
    assign c[413:412] = 0;
    assign c[415:414] = {a[1100], a[1101]};
    assign c[417:416] = 0;
    assign c[419:418] = 0;
    assign c[421:420] = {a[1102], a[1103]};
    assign c[423:422] = 0;
    assign c[425:424] = 0;
    assign c[427:426] = a[143:142];
    assign c[429:428] = 0;
    assign c[431:430] = 0;
    assign c[433:432] = a[861:860];
    assign c[435:434] = 0;
    assign c[437:436] = 0;
    assign c[439:438] = a[863:862];
    assign c[441:440] = 0;
    assign c[443:442] = 0;
    assign c[445:444] = {a[1110], a[1111]};
    assign c[447:446] = 0;
    assign c[449:448] = 0;
    assign c[451:450] = {a[1112], a[1113]};
    assign c[453:452] = 0;
    assign c[455:454] = 0;
    assign c[457:456] = {a[1114], a[1115]};
    assign c[459:458] = 0;
    assign c[461:460] = 0;
    assign c[463:462] = {a[1116], a[1117]};
    assign c[465:464] = 0;
    assign c[467:466] = 0;
    assign c[469:468] = {a[1118], a[1119]};
    assign c[471:470] = 0;
    assign c[473:472] = 0;
    assign c[475:474] = a[159:158];
    assign c[477:476] = 0;
    assign c[479:478] = 0;
    assign c[481:480] = a[877:876];
    assign c[483:482] = 0;
    assign c[485:484] = 0;
    assign c[487:486] = a[879:878];
    assign c[489:488] = 0;
    assign c[491:490] = 0;
    assign c[493:492] = {a[1126], a[1127]};
    assign c[495:494] = 0;
    assign c[497:496] = 0;
    assign c[499:498] = {a[1128], a[1129]};
    assign c[501:500] = 0;
    assign c[503:502] = 0;
    assign c[505:504] = {a[1130], a[1131]};
    assign c[507:506] = 0;
    assign c[509:508] = 0;
    assign c[511:510] = {a[1132], a[1133]};
    assign c[513:512] = 0;
    assign c[515:514] = 0;
    assign c[517:516] = {a[1134], a[1135]};
    assign c[519:518] = 0;
    assign c[521:520] = 0;
    assign c[523:522] = a[175:174];
    assign c[525:524] = 0;
    assign c[527:526] = 0;
    assign c[529:528] = a[893:892];
    assign c[531:530] = 0;
    assign c[533:532] = 0;
    assign c[535:534] = a[895:894];
    assign c[537:536] = 0;
    assign c[539:538] = 0;
    assign c[541:540] = {a[1142], a[1143]};
    assign c[543:542] = 0;
    assign c[545:544] = 0;
    assign c[547:546] = {a[1144], a[1145]};
    assign c[549:548] = 0;
    assign c[551:550] = 0;
    assign c[553:552] = {a[1146], a[1147]};
    assign c[555:554] = 0;
    assign c[557:556] = 0;
    assign c[559:558] = {a[1148], a[1149]};
    assign c[561:560] = 0;
    assign c[563:562] = 0;
    assign c[565:564] = {a[1150], a[1151]};
    assign c[567:566] = 0;
    assign c[569:568] = 0;
    assign c[571:570] = a[191:190];
    assign c[573:572] = 0;
    assign c[575:574] = 0;
    assign c[577:576] = a[909:908];
    assign c[579:578] = 0;
    assign c[581:580] = 0;
    assign c[583:582] = a[911:910];
    assign c[585:584] = 0;
    assign c[587:586] = 0;
    assign c[589:588] = {a[1158], a[1159]};
    assign c[591:590] = 0;
    assign c[593:592] = 0;
    assign c[595:594] = {a[1160], a[1161]};
    assign c[597:596] = 0;
    assign c[599:598] = 0;
    assign c[601:600] = {a[1162], a[1163]};
    assign c[603:602] = 0;
    assign c[605:604] = 0;
    assign c[607:606] = {a[1164], a[1165]};
    assign c[609:608] = 0;
    assign c[611:610] = 0;
    assign c[613:612] = {a[1166], a[1167]};
    assign c[615:614] = 0;
    assign c[617:616] = 0;
    assign c[619:618] = a[207:206];
    assign c[621:620] = 0;
    assign c[623:622] = 0;
    assign c[625:624] = a[925:924];
    assign c[627:626] = 0;
    assign c[629:628] = 0;
    assign c[631:630] = a[927:926];
    assign c[633:632] = 0;
    assign c[635:634] = 0;
    assign c[637:636] = {a[1174], a[1175]};
    assign c[639:638] = 0;
    assign c[641:640] = 0;
    assign c[643:642] = {a[1176], a[1177]};
    assign c[645:644] = 0;
    assign c[647:646] = 0;
    assign c[649:648] = {a[1178], a[1179]};
    assign c[651:650] = 0;
    assign c[653:652] = 0;
    assign c[655:654] = {a[1180], a[1181]};
    assign c[657:656] = 0;
    assign c[659:658] = 0;
    assign c[661:660] = {a[1182], a[1183]};
    assign c[663:662] = 0;
    assign c[665:664] = 0;
    assign c[667:666] = a[223:222];
    assign c[669:668] = 0;
    assign c[671:670] = 0;
    assign c[673:672] = 0;
    assign c[675:674] = 0;
    assign c[677:676] = 0;
    assign c[679:678] = 0;
    assign c[681:680] = 0;
    assign c[683:682] = 0;
    assign c[685:684] = 0;
    assign c[687:686] = 0;
    assign c[689:688] = 0;
    assign c[691:690] = 0;
    assign c[693:692] = 0;
    assign c[695:694] = 0;
    assign c[697:696] = 0;
    assign c[699:698] = 0;
    assign c[701:700] = 0;
    assign c[703:702] = 0;
    assign c[705:704] = 0;
    assign c[707:706] = 0;
    assign c[709:708] = 0;
    assign c[711:710] = 0;
    assign c[713:712] = 0;
    assign c[715:714] = 0;
    assign c[717:716] = 0;
    assign c[719:718] = 0;
    assign c[721:720] = 0;
    assign c[723:722] = 0;
    assign c[725:724] = 0;
    assign c[727:726] = 0;
    assign c[729:728] = 0;
    assign c[731:730] = 0;
    assign c[733:732] = 0;
    assign c[735:734] = 0;
    assign c[737:736] = 0;
    assign c[739:738] = 0;
    assign c[741:740] = 0;
    assign c[743:742] = 0;
    assign c[745:744] = 0;
    assign c[747:746] = 0;
    assign c[749:748] = 0;
    assign c[751:750] = 0;
    assign c[753:752] = 0;
    assign c[755:754] = 0;
    assign c[757:756] = 0;
    assign c[759:758] = 0;
    assign c[761:760] = 0;
    assign c[763:762] = 0;
    assign c[765:764] = 0;
    assign c[767:766] = 0;
    assign c[769:768] = 0;
    assign c[771:770] = 0;
    assign c[773:772] = 0;
    assign c[775:774] = 0;
    assign c[777:776] = 0;
    assign c[779:778] = 0;
    assign c[781:780] = 0;
    assign c[783:782] = 0;
    assign c[785:784] = 0;
    assign c[787:786] = 0;
    assign c[789:788] = 0;
    assign c[791:790] = 0;
    assign c[793:792] = 0;
    assign c[795:794] = 0;
    assign c[797:796] = 0;
    assign c[799:798] = 0;
    assign c[801:800] = 0;
    assign c[803:802] = 0;
    assign c[805:804] = 0;
    assign c[807:806] = 0;
    assign c[809:808] = 0;
    assign c[811:810] = 0;
    assign c[813:812] = 0;
    assign c[815:814] = 0;
    assign c[817:816] = 0;
    assign c[819:818] = 0;
    assign c[821:820] = 0;
    assign c[823:822] = 0;
    assign c[825:824] = 0;
    assign c[827:826] = 0;
    assign c[829:828] = 0;
    assign c[831:830] = 0;
    assign c[833:832] = 0;
    assign c[835:834] = 0;
    assign c[837:836] = 0;
    assign c[839:838] = 0;
    assign c[841:840] = 0;
    assign c[843:842] = 0;
    assign c[845:844] = 0;
    assign c[847:846] = 0;
    assign c[849:848] = 0;
    assign c[851:850] = 0;
    assign c[853:852] = 0;
    assign c[855:854] = 0;
    assign c[857:856] = 0;
    assign c[859:858] = 0;
    assign c[861:860] = 0;
    assign c[863:862] = 0;
    assign c[865:864] = 0;
    assign c[867:866] = 0;
    assign c[869:868] = 0;
    assign c[871:870] = 0;
    assign c[873:872] = 0;
    assign c[875:874] = 0;
    assign c[877:876] = 0;
    assign c[879:878] = 0;
    assign c[881:880] = 0;
    assign c[883:882] = 0;
    assign c[885:884] = 0;
    assign c[887:886] = 0;
    assign c[889:888] = 0;
    assign c[891:890] = 0;
    assign c[893:892] = 0;
    assign c[895:894] = 0;
    assign c[897:896] = 0;
    assign c[899:898] = 0;
    assign c[901:900] = 0;
    assign c[903:902] = 0;
    assign c[905:904] = 0;
    assign c[907:906] = 0;
    assign c[909:908] = 0;
    assign c[911:910] = 0;
    assign c[913:912] = 0;
    assign c[915:914] = 0;
    assign c[917:916] = 0;
    assign c[919:918] = 0;
    assign c[921:920] = 0;
    assign c[923:922] = 0;
    assign c[925:924] = 0;
    assign c[927:926] = 0;
    assign c[929:928] = 0;
    assign c[931:930] = 0;
    assign c[933:932] = 0;
    assign c[935:934] = 0;
    assign c[937:936] = 0;
    assign c[939:938] = 0;
    assign c[941:940] = 0;
    assign c[943:942] = 0;
    assign c[945:944] = 0;
    assign c[947:946] = 0;
    assign c[949:948] = 0;
    assign c[951:950] = 0;
    assign c[953:952] = 0;
    assign c[955:954] = 0;
    assign c[957:956] = 0;
    assign c[959:958] = 0;
    assign c[961:960] = 0;
    assign c[963:962] = 0;
    assign c[965:964] = 0;
    assign c[967:966] = 0;
    assign c[969:968] = 0;
    assign c[971:970] = 0;
    assign c[973:972] = 0;
    assign c[975:974] = 0;
    assign c[977:976] = 0;
    assign c[979:978] = 0;
    assign c[981:980] = 0;
    assign c[983:982] = 0;
    assign c[985:984] = 0;
    assign c[987:986] = 0;
    assign c[989:988] = 0;
    assign c[991:990] = 0;
    assign c[993:992] = 0;
    assign c[995:994] = 0;
    assign c[997:996] = 0;
    assign c[999:998] = 0;
    assign c[1001:1000] = 0;
    assign c[1003:1002] = 0;
    assign c[1005:1004] = 0;
    assign c[1007:1006] = 0;
    assign c[1009:1008] = 0;
    assign c[1011:1010] = 0;
    assign c[1013:1012] = 0;
    assign c[1015:1014] = 0;
    assign c[1017:1016] = 0;
    assign c[1019:1018] = 0;
    assign c[1021:1020] = 0;
    assign c[1023:1022] = 0;
    assign c[1025:1024] = 0;
    assign c[1027:1026] = 0;
    assign c[1029:1028] = 0;
    assign c[1031:1030] = 0;
    assign c[1033:1032] = 0;
    assign c[1035:1034] = 0;
    assign c[1037:1036] = 0;
    assign c[1039:1038] = 0;
    assign c[1041:1040] = 0;
    assign c[1043:1042] = 0;
    assign c[1045:1044] = 0;
    assign c[1047:1046] = 0;
    assign c[1049:1048] = 0;
    assign c[1051:1050] = 0;
    assign c[1053:1052] = 0;
    assign c[1055:1054] = 0;
    assign c[1057:1056] = 0;
    assign c[1059:1058] = 0;
    assign c[1061:1060] = 0;
    assign c[1063:1062] = 0;
    assign c[1065:1064] = 0;
    assign c[1067:1066] = 0;
    assign c[1069:1068] = 0;
    assign c[1071:1070] = 0;
    assign c[1073:1072] = 0;
    assign c[1075:1074] = 0;
    assign c[1077:1076] = 0;
    assign c[1079:1078] = 0;
    assign c[1081:1080] = 0;
    assign c[1083:1082] = 0;
    assign c[1085:1084] = 0;
    assign c[1087:1086] = 0;
    assign c[1089:1088] = 0;
    assign c[1091:1090] = 0;
    assign c[1093:1092] = 0;
    assign c[1095:1094] = 0;
    assign c[1097:1096] = 0;
    assign c[1099:1098] = 0;
    assign c[1101:1100] = 0;
    assign c[1103:1102] = 0;
    assign c[1105:1104] = 0;
    assign c[1107:1106] = 0;
    assign c[1109:1108] = 0;
    assign c[1111:1110] = 0;
    assign c[1113:1112] = 0;
    assign c[1115:1114] = 0;
    assign c[1117:1116] = 0;
    assign c[1119:1118] = 0;
    assign c[1121:1120] = 0;
    assign c[1123:1122] = 0;
    assign c[1125:1124] = 0;
    assign c[1127:1126] = 0;
    assign c[1129:1128] = 0;
    assign c[1131:1130] = 0;
    assign c[1133:1132] = 0;
    assign c[1135:1134] = 0;
    assign c[1137:1136] = 0;
    assign c[1139:1138] = 0;
    assign c[1141:1140] = 0;
    assign c[1143:1142] = 0;
    assign c[1145:1144] = 0;
    assign c[1147:1146] = 0;
    assign c[1149:1148] = 0;
    assign c[1151:1150] = 0;
    assign c[1153:1152] = 0;
    assign c[1155:1154] = 0;
    assign c[1157:1156] = 0;
    assign c[1159:1158] = 0;
    assign c[1161:1160] = 0;
    assign c[1163:1162] = 0;
    assign c[1165:1164] = 0;
    assign c[1167:1166] = 0;
    assign c[1169:1168] = 0;
    assign c[1171:1170] = 0;
    assign c[1173:1172] = 0;
    assign c[1175:1174] = 0;
    assign c[1177:1176] = 0;
    assign c[1179:1178] = 0;
    assign c[1181:1180] = 0;
    assign c[1183:1182] = 0;
    assign c[1185:1184] = 0;
endmodule
