`define SIMULATION_MEMORY

module shift_register_group_18_32_3 (
	input clk,
	input enable,
	input [17:0] in_0,
	output [17:0] out_0,
	input [17:0] in_1,
	output [17:0] out_1,
	input [17:0] in_2,
	output [17:0] out_2,
	input [17:0] in_3,
	output [17:0] out_3,
	input [17:0] in_4,
	output [17:0] out_4,
	input [17:0] in_5,
	output [17:0] out_5,
	input [17:0] in_6,
	output [17:0] out_6,
	input [17:0] in_7,
	output [17:0] out_7,
	input [17:0] in_8,
	output [17:0] out_8,
	input [17:0] in_9,
	output [17:0] out_9,
	input [17:0] in_10,
	output [17:0] out_10,
	input [17:0] in_11,
	output [17:0] out_11,
	input [17:0] in_12,
	output [17:0] out_12,
	input [17:0] in_13,
	output [17:0] out_13,
	input [17:0] in_14,
	output [17:0] out_14,
	input [17:0] in_15,
	output [17:0] out_15,
	input [17:0] in_16,
	output [17:0] out_16,
	input [17:0] in_17,
	output [17:0] out_17,
	input [17:0] in_18,
	output [17:0] out_18,
	input [17:0] in_19,
	output [17:0] out_19,
	input [17:0] in_20,
	output [17:0] out_20,
	input [17:0] in_21,
	output [17:0] out_21,
	input [17:0] in_22,
	output [17:0] out_22,
	input [17:0] in_23,
	output [17:0] out_23,
	input [17:0] in_24,
	output [17:0] out_24,
	input [17:0] in_25,
	output [17:0] out_25,
	input [17:0] in_26,
	output [17:0] out_26,
	input [17:0] in_27,
	output [17:0] out_27,
	input [17:0] in_28,
	output [17:0] out_28,
	input [17:0] in_29,
	output [17:0] out_29,
	input [17:0] in_30,
	output [17:0] out_30,
	input [17:0] in_31,
	output [17:0] out_31,
	input reset
);

shift_register_unit_18_3 shift_register_unit_18_3_inst_0 (
	.clk(clk),
	.reset(reset),
	.enable(enable),
	.in(in_0),
	.out(out_0)
);

shift_register_unit_18_3 shift_register_unit_18_3_inst_1 (
	.clk(clk),
	.reset(reset),
	.enable(enable),
	.in(in_1),
	.out(out_1)
);

shift_register_unit_18_3 shift_register_unit_18_3_inst_2 (
	.clk(clk),
	.reset(reset),
	.enable(enable),
	.in(in_2),
	.out(out_2)
);

shift_register_unit_18_3 shift_register_unit_18_3_inst_3 (
	.clk(clk),
	.reset(reset),
	.enable(enable),
	.in(in_3),
	.out(out_3)
);

shift_register_unit_18_3 shift_register_unit_18_3_inst_4 (
	.clk(clk),
	.reset(reset),
	.enable(enable),
	.in(in_4),
	.out(out_4)
);

shift_register_unit_18_3 shift_register_unit_18_3_inst_5 (
	.clk(clk),
	.reset(reset),
	.enable(enable),
	.in(in_5),
	.out(out_5)
);

shift_register_unit_18_3 shift_register_unit_18_3_inst_6 (
	.clk(clk),
	.reset(reset),
	.enable(enable),
	.in(in_6),
	.out(out_6)
);

shift_register_unit_18_3 shift_register_unit_18_3_inst_7 (
	.clk(clk),
	.reset(reset),
	.enable(enable),
	.in(in_7),
	.out(out_7)
);

shift_register_unit_18_3 shift_register_unit_18_3_inst_8 (
	.clk(clk),
	.reset(reset),
	.enable(enable),
	.in(in_8),
	.out(out_8)
);

shift_register_unit_18_3 shift_register_unit_18_3_inst_9 (
	.clk(clk),
	.reset(reset),
	.enable(enable),
	.in(in_9),
	.out(out_9)
);

shift_register_unit_18_3 shift_register_unit_18_3_inst_10 (
	.clk(clk),
	.reset(reset),
	.enable(enable),
	.in(in_10),
	.out(out_10)
);

shift_register_unit_18_3 shift_register_unit_18_3_inst_11 (
	.clk(clk),
	.reset(reset),
	.enable(enable),
	.in(in_11),
	.out(out_11)
);

shift_register_unit_18_3 shift_register_unit_18_3_inst_12 (
	.clk(clk),
	.reset(reset),
	.enable(enable),
	.in(in_12),
	.out(out_12)
);

shift_register_unit_18_3 shift_register_unit_18_3_inst_13 (
	.clk(clk),
	.reset(reset),
	.enable(enable),
	.in(in_13),
	.out(out_13)
);

shift_register_unit_18_3 shift_register_unit_18_3_inst_14 (
	.clk(clk),
	.reset(reset),
	.enable(enable),
	.in(in_14),
	.out(out_14)
);

shift_register_unit_18_3 shift_register_unit_18_3_inst_15 (
	.clk(clk),
	.reset(reset),
	.enable(enable),
	.in(in_15),
	.out(out_15)
);

shift_register_unit_18_3 shift_register_unit_18_3_inst_16 (
	.clk(clk),
	.reset(reset),
	.enable(enable),
	.in(in_16),
	.out(out_16)
);

shift_register_unit_18_3 shift_register_unit_18_3_inst_17 (
	.clk(clk),
	.reset(reset),
	.enable(enable),
	.in(in_17),
	.out(out_17)
);

shift_register_unit_18_3 shift_register_unit_18_3_inst_18 (
	.clk(clk),
	.reset(reset),
	.enable(enable),
	.in(in_18),
	.out(out_18)
);

shift_register_unit_18_3 shift_register_unit_18_3_inst_19 (
	.clk(clk),
	.reset(reset),
	.enable(enable),
	.in(in_19),
	.out(out_19)
);

shift_register_unit_18_3 shift_register_unit_18_3_inst_20 (
	.clk(clk),
	.reset(reset),
	.enable(enable),
	.in(in_20),
	.out(out_20)
);

shift_register_unit_18_3 shift_register_unit_18_3_inst_21 (
	.clk(clk),
	.reset(reset),
	.enable(enable),
	.in(in_21),
	.out(out_21)
);

shift_register_unit_18_3 shift_register_unit_18_3_inst_22 (
	.clk(clk),
	.reset(reset),
	.enable(enable),
	.in(in_22),
	.out(out_22)
);

shift_register_unit_18_3 shift_register_unit_18_3_inst_23 (
	.clk(clk),
	.reset(reset),
	.enable(enable),
	.in(in_23),
	.out(out_23)
);

shift_register_unit_18_3 shift_register_unit_18_3_inst_24 (
	.clk(clk),
	.reset(reset),
	.enable(enable),
	.in(in_24),
	.out(out_24)
);

shift_register_unit_18_3 shift_register_unit_18_3_inst_25 (
	.clk(clk),
	.reset(reset),
	.enable(enable),
	.in(in_25),
	.out(out_25)
);

shift_register_unit_18_3 shift_register_unit_18_3_inst_26 (
	.clk(clk),
	.reset(reset),
	.enable(enable),
	.in(in_26),
	.out(out_26)
);

shift_register_unit_18_3 shift_register_unit_18_3_inst_27 (
	.clk(clk),
	.reset(reset),
	.enable(enable),
	.in(in_27),
	.out(out_27)
);

shift_register_unit_18_3 shift_register_unit_18_3_inst_28 (
	.clk(clk),
	.reset(reset),
	.enable(enable),
	.in(in_28),
	.out(out_28)
);

shift_register_unit_18_3 shift_register_unit_18_3_inst_29 (
	.clk(clk),
	.reset(reset),
	.enable(enable),
	.in(in_29),
	.out(out_29)
);

shift_register_unit_18_3 shift_register_unit_18_3_inst_30 (
	.clk(clk),
	.reset(reset),
	.enable(enable),
	.in(in_30),
	.out(out_30)
);

shift_register_unit_18_3 shift_register_unit_18_3_inst_31 (
	.clk(clk),
	.reset(reset),
	.enable(enable),
	.in(in_31),
	.out(out_31)
);

endmodule

module shift_register_unit_18_3 (
	input clk,
	input reset,
	input enable,
	input [17:0] in,
	output [17:0] out
);

reg [17:0] shift_registers_0;
reg [17:0] shift_registers_1;
reg [17:0] shift_registers_2;
always @ (posedge clk) begin
	if (reset) begin
		shift_registers_0 <= 18'd0;
		shift_registers_1 <= 18'd0;
		shift_registers_2 <= 18'd0;
	end else if (enable) begin
		shift_registers_0 <= in;
		shift_registers_1 <= shift_registers_0;
		shift_registers_2 <= shift_registers_1;
	end
end

assign out = shift_registers_2;

endmodule



