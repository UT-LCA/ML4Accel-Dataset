
module myproject_mul_16s_8ns_24_2_0(
    clk,
    reset,
    ce,
    din0,
    din1,
    dout);

parameter ID = 32'd1;
parameter NUM_STAGE = 32'd1;
parameter din0_WIDTH = 32'd1;
parameter din1_WIDTH = 32'd1;
parameter dout_WIDTH = 32'd1;
input clk;
input reset;
input ce;
input[din0_WIDTH - 1:0] din0;
input[din1_WIDTH - 1:0] din1;
output[dout_WIDTH - 1:0] dout;



myproject_mul_16s_8ns_24_2_0_MulnS_5 myproject_mul_16s_8ns_24_2_0_MulnS_5_U(
    .clk( clk ),
    .ce( ce ),
    .a( din0 ),
    .b( din1 ),
    .p( dout ));

endmodule
module myproject_mul_16s_8ns_24_2_0_MulnS_5(clk, ce, a, b, p);
input clk;
input ce;
input  [16 - 1 : 0] a;
input [8 - 1 : 0] b;
output[24 - 1 : 0] p;
reg  [24 - 1 : 0] p;
wire  [24 - 1 : 0] tmp_product;

assign tmp_product = (a) * ({1'b0, b});
always @ (posedge clk) begin
    if (ce) begin
        p <= tmp_product;
    end
end
endmodule
