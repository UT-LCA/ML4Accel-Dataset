
module dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s (
        ap_clk,
        ap_rst,
        data_0_V_read,
        data_1_V_read,
        data_2_V_read,
        data_3_V_read,
        data_4_V_read,
        data_5_V_read,
        data_6_V_read,
        data_7_V_read,
        data_8_V_read,
        data_9_V_read,
        data_10_V_read,
        data_11_V_read,
        data_12_V_read,
        data_13_V_read,
        data_14_V_read,
        data_15_V_read,
        data_16_V_read,
        data_17_V_read,
        data_18_V_read,
        data_19_V_read,
        data_20_V_read,
        data_21_V_read,
        data_22_V_read,
        data_23_V_read,
        data_24_V_read,
        data_25_V_read,
        data_26_V_read,
        data_27_V_read,
        data_28_V_read,
        data_29_V_read,
        data_30_V_read,
        data_31_V_read,
        data_32_V_read,
        data_33_V_read,
        data_34_V_read,
        data_35_V_read,
        data_36_V_read,
        data_37_V_read,
        data_38_V_read,
        data_39_V_read,
        data_40_V_read,
        data_41_V_read,
        data_42_V_read,
        data_43_V_read,
        data_44_V_read,
        data_45_V_read,
        data_46_V_read,
        data_47_V_read,
        data_48_V_read,
        data_49_V_read,
        data_50_V_read,
        data_51_V_read,
        data_52_V_read,
        data_53_V_read,
        data_54_V_read,
        data_55_V_read,
        data_56_V_read,
        data_57_V_read,
        data_58_V_read,
        data_59_V_read,
        data_60_V_read,
        data_61_V_read,
        data_62_V_read,
        data_63_V_read,
        ap_return_0,
        ap_return_1,
        ap_return_2,
        ap_return_3,
        ap_return_4,
        ap_return_5,
        ap_return_6,
        ap_return_7,
        ap_return_8,
        ap_return_9,
        ap_return_10,
        ap_return_11,
        ap_return_12,
        ap_return_13,
        ap_return_14,
        ap_return_15,
        ap_return_16,
        ap_return_17,
        ap_return_18,
        ap_return_19,
        ap_return_20,
        ap_return_21,
        ap_return_22,
        ap_return_23,
        ap_return_24,
        ap_return_25,
        ap_return_26,
        ap_return_27,
        ap_return_28,
        ap_return_29,
        ap_return_30,
        ap_return_31,
        ap_ce
);


input   ap_clk;
input   ap_rst;
input  [15:0] data_0_V_read;
input  [15:0] data_1_V_read;
input  [15:0] data_2_V_read;
input  [15:0] data_3_V_read;
input  [15:0] data_4_V_read;
input  [15:0] data_5_V_read;
input  [15:0] data_6_V_read;
input  [15:0] data_7_V_read;
input  [15:0] data_8_V_read;
input  [15:0] data_9_V_read;
input  [15:0] data_10_V_read;
input  [15:0] data_11_V_read;
input  [15:0] data_12_V_read;
input  [15:0] data_13_V_read;
input  [15:0] data_14_V_read;
input  [15:0] data_15_V_read;
input  [15:0] data_16_V_read;
input  [15:0] data_17_V_read;
input  [15:0] data_18_V_read;
input  [15:0] data_19_V_read;
input  [15:0] data_20_V_read;
input  [15:0] data_21_V_read;
input  [15:0] data_22_V_read;
input  [15:0] data_23_V_read;
input  [15:0] data_24_V_read;
input  [15:0] data_25_V_read;
input  [15:0] data_26_V_read;
input  [15:0] data_27_V_read;
input  [15:0] data_28_V_read;
input  [15:0] data_29_V_read;
input  [15:0] data_30_V_read;
input  [15:0] data_31_V_read;
input  [15:0] data_32_V_read;
input  [15:0] data_33_V_read;
input  [15:0] data_34_V_read;
input  [15:0] data_35_V_read;
input  [15:0] data_36_V_read;
input  [15:0] data_37_V_read;
input  [15:0] data_38_V_read;
input  [15:0] data_39_V_read;
input  [15:0] data_40_V_read;
input  [15:0] data_41_V_read;
input  [15:0] data_42_V_read;
input  [15:0] data_43_V_read;
input  [15:0] data_44_V_read;
input  [15:0] data_45_V_read;
input  [15:0] data_46_V_read;
input  [15:0] data_47_V_read;
input  [15:0] data_48_V_read;
input  [15:0] data_49_V_read;
input  [15:0] data_50_V_read;
input  [15:0] data_51_V_read;
input  [15:0] data_52_V_read;
input  [15:0] data_53_V_read;
input  [15:0] data_54_V_read;
input  [15:0] data_55_V_read;
input  [15:0] data_56_V_read;
input  [15:0] data_57_V_read;
input  [15:0] data_58_V_read;
input  [15:0] data_59_V_read;
input  [15:0] data_60_V_read;
input  [15:0] data_61_V_read;
input  [15:0] data_62_V_read;
input  [15:0] data_63_V_read;
output  [15:0] ap_return_0;
output  [15:0] ap_return_1;
output  [15:0] ap_return_2;
output  [15:0] ap_return_3;
output  [15:0] ap_return_4;
output  [15:0] ap_return_5;
output  [15:0] ap_return_6;
output  [15:0] ap_return_7;
output  [15:0] ap_return_8;
output  [15:0] ap_return_9;
output  [15:0] ap_return_10;
output  [15:0] ap_return_11;
output  [15:0] ap_return_12;
output  [15:0] ap_return_13;
output  [15:0] ap_return_14;
output  [15:0] ap_return_15;
output  [15:0] ap_return_16;
output  [15:0] ap_return_17;
output  [15:0] ap_return_18;
output  [15:0] ap_return_19;
output  [15:0] ap_return_20;
output  [15:0] ap_return_21;
output  [15:0] ap_return_22;
output  [15:0] ap_return_23;
output  [15:0] ap_return_24;
output  [15:0] ap_return_25;
output  [15:0] ap_return_26;
output  [15:0] ap_return_27;
output  [15:0] ap_return_28;
output  [15:0] ap_return_29;
output  [15:0] ap_return_30;
output  [15:0] ap_return_31;
input   ap_ce;

reg[15:0] ap_return_0;
reg[15:0] ap_return_1;
reg[15:0] ap_return_2;
reg[15:0] ap_return_3;
reg[15:0] ap_return_4;
reg[15:0] ap_return_5;
reg[15:0] ap_return_6;
reg[15:0] ap_return_7;
reg[15:0] ap_return_8;
reg[15:0] ap_return_9;
reg[15:0] ap_return_10;
reg[15:0] ap_return_11;
reg[15:0] ap_return_12;
reg[15:0] ap_return_13;
reg[15:0] ap_return_14;
reg[15:0] ap_return_15;
reg[15:0] ap_return_16;
reg[15:0] ap_return_17;
reg[15:0] ap_return_18;
reg[15:0] ap_return_19;
reg[15:0] ap_return_20;
reg[15:0] ap_return_21;
reg[15:0] ap_return_22;
reg[15:0] ap_return_23;
reg[15:0] ap_return_24;
reg[15:0] ap_return_25;
reg[15:0] ap_return_26;
reg[15:0] ap_return_27;
reg[15:0] ap_return_28;
reg[15:0] ap_return_29;
reg[15:0] ap_return_30;
reg[15:0] ap_return_31;

reg   [15:0] data_63_V_read_3_reg_8620;
wire    ap_block_state1_pp0_stage0_iter0;
wire    ap_block_state2_pp0_stage0_iter1;
wire    ap_block_state3_pp0_stage0_iter2;
wire    ap_block_state4_pp0_stage0_iter3;
wire    ap_block_state5_pp0_stage0_iter4;
wire    ap_block_state6_pp0_stage0_iter5;
wire    ap_block_state7_pp0_stage0_iter6;
wire    ap_block_state8_pp0_stage0_iter7;
wire    ap_block_state9_pp0_stage0_iter8;
wire    ap_block_state10_pp0_stage0_iter9;
wire    ap_block_state11_pp0_stage0_iter10;
wire    ap_block_state12_pp0_stage0_iter11;
wire    ap_block_state13_pp0_stage0_iter12;
wire    ap_block_state14_pp0_stage0_iter13;
wire    ap_block_state15_pp0_stage0_iter14;
wire    ap_block_state16_pp0_stage0_iter15;
wire    ap_block_state17_pp0_stage0_iter16;
wire    ap_block_state18_pp0_stage0_iter17;
wire    ap_block_pp0_stage0_11001;
reg   [15:0] data_63_V_read_3_reg_8620_pp0_iter1_reg;
reg   [15:0] data_63_V_read_3_reg_8620_pp0_iter2_reg;
reg   [15:0] data_63_V_read_3_reg_8620_pp0_iter3_reg;
reg   [15:0] data_63_V_read_3_reg_8620_pp0_iter4_reg;
reg   [15:0] data_63_V_read_3_reg_8620_pp0_iter5_reg;
reg   [15:0] data_63_V_read_3_reg_8620_pp0_iter6_reg;
reg   [15:0] data_63_V_read_3_reg_8620_pp0_iter7_reg;
reg   [15:0] data_63_V_read_3_reg_8620_pp0_iter8_reg;
reg   [15:0] data_63_V_read_3_reg_8620_pp0_iter9_reg;
reg   [15:0] data_63_V_read_3_reg_8620_pp0_iter10_reg;
reg   [15:0] data_63_V_read_3_reg_8620_pp0_iter11_reg;
reg   [15:0] data_63_V_read_3_reg_8620_pp0_iter12_reg;
reg   [15:0] data_63_V_read_3_reg_8620_pp0_iter13_reg;
reg   [15:0] data_63_V_read_3_reg_8620_pp0_iter14_reg;
reg   [15:0] data_63_V_read_3_reg_8620_pp0_iter15_reg;
reg   [15:0] data_63_V_read_3_reg_8620_pp0_iter16_reg;
reg   [15:0] data_62_V_read_3_reg_8645;
reg   [15:0] data_62_V_read_3_reg_8645_pp0_iter1_reg;
reg   [15:0] data_62_V_read_3_reg_8645_pp0_iter2_reg;
reg   [15:0] data_62_V_read_3_reg_8645_pp0_iter3_reg;
reg   [15:0] data_62_V_read_3_reg_8645_pp0_iter4_reg;
reg   [15:0] data_62_V_read_3_reg_8645_pp0_iter5_reg;
reg   [15:0] data_62_V_read_3_reg_8645_pp0_iter6_reg;
reg   [15:0] data_62_V_read_3_reg_8645_pp0_iter7_reg;
reg   [15:0] data_62_V_read_3_reg_8645_pp0_iter8_reg;
reg   [15:0] data_62_V_read_3_reg_8645_pp0_iter9_reg;
reg   [15:0] data_62_V_read_3_reg_8645_pp0_iter10_reg;
reg   [15:0] data_62_V_read_3_reg_8645_pp0_iter11_reg;
reg   [15:0] data_62_V_read_3_reg_8645_pp0_iter12_reg;
reg   [15:0] data_62_V_read_3_reg_8645_pp0_iter13_reg;
reg   [15:0] data_62_V_read_3_reg_8645_pp0_iter14_reg;
reg   [15:0] data_62_V_read_3_reg_8645_pp0_iter15_reg;
reg   [15:0] data_62_V_read_3_reg_8645_pp0_iter16_reg;
reg   [15:0] data_61_V_read62_reg_8663;
reg   [15:0] data_61_V_read62_reg_8663_pp0_iter1_reg;
reg   [15:0] data_61_V_read62_reg_8663_pp0_iter2_reg;
reg   [15:0] data_61_V_read62_reg_8663_pp0_iter3_reg;
reg   [15:0] data_61_V_read62_reg_8663_pp0_iter4_reg;
reg   [15:0] data_61_V_read62_reg_8663_pp0_iter5_reg;
reg   [15:0] data_61_V_read62_reg_8663_pp0_iter6_reg;
reg   [15:0] data_61_V_read62_reg_8663_pp0_iter7_reg;
reg   [15:0] data_61_V_read62_reg_8663_pp0_iter8_reg;
reg   [15:0] data_61_V_read62_reg_8663_pp0_iter9_reg;
reg   [15:0] data_61_V_read62_reg_8663_pp0_iter10_reg;
reg   [15:0] data_61_V_read62_reg_8663_pp0_iter11_reg;
reg   [15:0] data_61_V_read62_reg_8663_pp0_iter12_reg;
reg   [15:0] data_61_V_read62_reg_8663_pp0_iter13_reg;
reg   [15:0] data_61_V_read62_reg_8663_pp0_iter14_reg;
reg   [15:0] data_61_V_read62_reg_8663_pp0_iter15_reg;
reg   [15:0] data_61_V_read62_reg_8663_pp0_iter16_reg;
reg   [15:0] data_60_V_read61_reg_8691;
reg   [15:0] data_60_V_read61_reg_8691_pp0_iter1_reg;
reg   [15:0] data_60_V_read61_reg_8691_pp0_iter2_reg;
reg   [15:0] data_60_V_read61_reg_8691_pp0_iter3_reg;
reg   [15:0] data_60_V_read61_reg_8691_pp0_iter4_reg;
reg   [15:0] data_60_V_read61_reg_8691_pp0_iter5_reg;
reg   [15:0] data_60_V_read61_reg_8691_pp0_iter6_reg;
reg   [15:0] data_60_V_read61_reg_8691_pp0_iter7_reg;
reg   [15:0] data_60_V_read61_reg_8691_pp0_iter8_reg;
reg   [15:0] data_60_V_read61_reg_8691_pp0_iter9_reg;
reg   [15:0] data_60_V_read61_reg_8691_pp0_iter10_reg;
reg   [15:0] data_60_V_read61_reg_8691_pp0_iter11_reg;
reg   [15:0] data_60_V_read61_reg_8691_pp0_iter12_reg;
reg   [15:0] data_60_V_read61_reg_8691_pp0_iter13_reg;
reg   [15:0] data_60_V_read61_reg_8691_pp0_iter14_reg;
reg   [15:0] data_60_V_read61_reg_8691_pp0_iter15_reg;
reg   [15:0] data_60_V_read61_reg_8691_pp0_iter16_reg;
reg   [15:0] data_59_V_read_3_reg_8724;
reg   [15:0] data_59_V_read_3_reg_8724_pp0_iter1_reg;
reg   [15:0] data_59_V_read_3_reg_8724_pp0_iter2_reg;
reg   [15:0] data_59_V_read_3_reg_8724_pp0_iter3_reg;
reg   [15:0] data_59_V_read_3_reg_8724_pp0_iter4_reg;
reg   [15:0] data_59_V_read_3_reg_8724_pp0_iter5_reg;
reg   [15:0] data_59_V_read_3_reg_8724_pp0_iter6_reg;
reg   [15:0] data_59_V_read_3_reg_8724_pp0_iter7_reg;
reg   [15:0] data_59_V_read_3_reg_8724_pp0_iter8_reg;
reg   [15:0] data_59_V_read_3_reg_8724_pp0_iter9_reg;
reg   [15:0] data_59_V_read_3_reg_8724_pp0_iter10_reg;
reg   [15:0] data_59_V_read_3_reg_8724_pp0_iter11_reg;
reg   [15:0] data_59_V_read_3_reg_8724_pp0_iter12_reg;
reg   [15:0] data_59_V_read_3_reg_8724_pp0_iter13_reg;
reg   [15:0] data_59_V_read_3_reg_8724_pp0_iter14_reg;
reg   [15:0] data_59_V_read_3_reg_8724_pp0_iter15_reg;
reg   [15:0] data_59_V_read_3_reg_8724_pp0_iter16_reg;
reg   [15:0] data_58_V_read_3_reg_8756;
reg   [15:0] data_58_V_read_3_reg_8756_pp0_iter1_reg;
reg   [15:0] data_58_V_read_3_reg_8756_pp0_iter2_reg;
reg   [15:0] data_58_V_read_3_reg_8756_pp0_iter3_reg;
reg   [15:0] data_58_V_read_3_reg_8756_pp0_iter4_reg;
reg   [15:0] data_58_V_read_3_reg_8756_pp0_iter5_reg;
reg   [15:0] data_58_V_read_3_reg_8756_pp0_iter6_reg;
reg   [15:0] data_58_V_read_3_reg_8756_pp0_iter7_reg;
reg   [15:0] data_58_V_read_3_reg_8756_pp0_iter8_reg;
reg   [15:0] data_58_V_read_3_reg_8756_pp0_iter9_reg;
reg   [15:0] data_58_V_read_3_reg_8756_pp0_iter10_reg;
reg   [15:0] data_58_V_read_3_reg_8756_pp0_iter11_reg;
reg   [15:0] data_58_V_read_3_reg_8756_pp0_iter12_reg;
reg   [15:0] data_58_V_read_3_reg_8756_pp0_iter13_reg;
reg   [15:0] data_58_V_read_3_reg_8756_pp0_iter14_reg;
reg   [15:0] data_58_V_read_3_reg_8756_pp0_iter15_reg;
reg   [15:0] data_57_V_read_3_reg_8786;
reg   [15:0] data_57_V_read_3_reg_8786_pp0_iter1_reg;
reg   [15:0] data_57_V_read_3_reg_8786_pp0_iter2_reg;
reg   [15:0] data_57_V_read_3_reg_8786_pp0_iter3_reg;
reg   [15:0] data_57_V_read_3_reg_8786_pp0_iter4_reg;
reg   [15:0] data_57_V_read_3_reg_8786_pp0_iter5_reg;
reg   [15:0] data_57_V_read_3_reg_8786_pp0_iter6_reg;
reg   [15:0] data_57_V_read_3_reg_8786_pp0_iter7_reg;
reg   [15:0] data_57_V_read_3_reg_8786_pp0_iter8_reg;
reg   [15:0] data_57_V_read_3_reg_8786_pp0_iter9_reg;
reg   [15:0] data_57_V_read_3_reg_8786_pp0_iter10_reg;
reg   [15:0] data_57_V_read_3_reg_8786_pp0_iter11_reg;
reg   [15:0] data_57_V_read_3_reg_8786_pp0_iter12_reg;
reg   [15:0] data_57_V_read_3_reg_8786_pp0_iter13_reg;
reg   [15:0] data_57_V_read_3_reg_8786_pp0_iter14_reg;
reg   [15:0] data_57_V_read_3_reg_8786_pp0_iter15_reg;
reg   [15:0] data_56_V_read_3_reg_8814;
reg   [15:0] data_56_V_read_3_reg_8814_pp0_iter1_reg;
reg   [15:0] data_56_V_read_3_reg_8814_pp0_iter2_reg;
reg   [15:0] data_56_V_read_3_reg_8814_pp0_iter3_reg;
reg   [15:0] data_56_V_read_3_reg_8814_pp0_iter4_reg;
reg   [15:0] data_56_V_read_3_reg_8814_pp0_iter5_reg;
reg   [15:0] data_56_V_read_3_reg_8814_pp0_iter6_reg;
reg   [15:0] data_56_V_read_3_reg_8814_pp0_iter7_reg;
reg   [15:0] data_56_V_read_3_reg_8814_pp0_iter8_reg;
reg   [15:0] data_56_V_read_3_reg_8814_pp0_iter9_reg;
reg   [15:0] data_56_V_read_3_reg_8814_pp0_iter10_reg;
reg   [15:0] data_56_V_read_3_reg_8814_pp0_iter11_reg;
reg   [15:0] data_56_V_read_3_reg_8814_pp0_iter12_reg;
reg   [15:0] data_56_V_read_3_reg_8814_pp0_iter13_reg;
reg   [15:0] data_56_V_read_3_reg_8814_pp0_iter14_reg;
reg   [15:0] data_56_V_read_3_reg_8814_pp0_iter15_reg;
reg   [15:0] data_55_V_read_3_reg_8844;
reg   [15:0] data_55_V_read_3_reg_8844_pp0_iter1_reg;
reg   [15:0] data_55_V_read_3_reg_8844_pp0_iter2_reg;
reg   [15:0] data_55_V_read_3_reg_8844_pp0_iter3_reg;
reg   [15:0] data_55_V_read_3_reg_8844_pp0_iter4_reg;
reg   [15:0] data_55_V_read_3_reg_8844_pp0_iter5_reg;
reg   [15:0] data_55_V_read_3_reg_8844_pp0_iter6_reg;
reg   [15:0] data_55_V_read_3_reg_8844_pp0_iter7_reg;
reg   [15:0] data_55_V_read_3_reg_8844_pp0_iter8_reg;
reg   [15:0] data_55_V_read_3_reg_8844_pp0_iter9_reg;
reg   [15:0] data_55_V_read_3_reg_8844_pp0_iter10_reg;
reg   [15:0] data_55_V_read_3_reg_8844_pp0_iter11_reg;
reg   [15:0] data_55_V_read_3_reg_8844_pp0_iter12_reg;
reg   [15:0] data_55_V_read_3_reg_8844_pp0_iter13_reg;
reg   [15:0] data_55_V_read_3_reg_8844_pp0_iter14_reg;
reg   [15:0] data_55_V_read_3_reg_8844_pp0_iter15_reg;
reg   [15:0] data_54_V_read_3_reg_8873;
reg   [15:0] data_54_V_read_3_reg_8873_pp0_iter1_reg;
reg   [15:0] data_54_V_read_3_reg_8873_pp0_iter2_reg;
reg   [15:0] data_54_V_read_3_reg_8873_pp0_iter3_reg;
reg   [15:0] data_54_V_read_3_reg_8873_pp0_iter4_reg;
reg   [15:0] data_54_V_read_3_reg_8873_pp0_iter5_reg;
reg   [15:0] data_54_V_read_3_reg_8873_pp0_iter6_reg;
reg   [15:0] data_54_V_read_3_reg_8873_pp0_iter7_reg;
reg   [15:0] data_54_V_read_3_reg_8873_pp0_iter8_reg;
reg   [15:0] data_54_V_read_3_reg_8873_pp0_iter9_reg;
reg   [15:0] data_54_V_read_3_reg_8873_pp0_iter10_reg;
reg   [15:0] data_54_V_read_3_reg_8873_pp0_iter11_reg;
reg   [15:0] data_54_V_read_3_reg_8873_pp0_iter12_reg;
reg   [15:0] data_54_V_read_3_reg_8873_pp0_iter13_reg;
reg   [15:0] data_54_V_read_3_reg_8873_pp0_iter14_reg;
reg   [15:0] data_53_V_read_3_reg_8899;
reg   [15:0] data_53_V_read_3_reg_8899_pp0_iter1_reg;
reg   [15:0] data_53_V_read_3_reg_8899_pp0_iter2_reg;
reg   [15:0] data_53_V_read_3_reg_8899_pp0_iter3_reg;
reg   [15:0] data_53_V_read_3_reg_8899_pp0_iter4_reg;
reg   [15:0] data_53_V_read_3_reg_8899_pp0_iter5_reg;
reg   [15:0] data_53_V_read_3_reg_8899_pp0_iter6_reg;
reg   [15:0] data_53_V_read_3_reg_8899_pp0_iter7_reg;
reg   [15:0] data_53_V_read_3_reg_8899_pp0_iter8_reg;
reg   [15:0] data_53_V_read_3_reg_8899_pp0_iter9_reg;
reg   [15:0] data_53_V_read_3_reg_8899_pp0_iter10_reg;
reg   [15:0] data_53_V_read_3_reg_8899_pp0_iter11_reg;
reg   [15:0] data_53_V_read_3_reg_8899_pp0_iter12_reg;
reg   [15:0] data_53_V_read_3_reg_8899_pp0_iter13_reg;
reg   [15:0] data_53_V_read_3_reg_8899_pp0_iter14_reg;
reg   [15:0] data_52_V_read_3_reg_8928;
reg   [15:0] data_52_V_read_3_reg_8928_pp0_iter1_reg;
reg   [15:0] data_52_V_read_3_reg_8928_pp0_iter2_reg;
reg   [15:0] data_52_V_read_3_reg_8928_pp0_iter3_reg;
reg   [15:0] data_52_V_read_3_reg_8928_pp0_iter4_reg;
reg   [15:0] data_52_V_read_3_reg_8928_pp0_iter5_reg;
reg   [15:0] data_52_V_read_3_reg_8928_pp0_iter6_reg;
reg   [15:0] data_52_V_read_3_reg_8928_pp0_iter7_reg;
reg   [15:0] data_52_V_read_3_reg_8928_pp0_iter8_reg;
reg   [15:0] data_52_V_read_3_reg_8928_pp0_iter9_reg;
reg   [15:0] data_52_V_read_3_reg_8928_pp0_iter10_reg;
reg   [15:0] data_52_V_read_3_reg_8928_pp0_iter11_reg;
reg   [15:0] data_52_V_read_3_reg_8928_pp0_iter12_reg;
reg   [15:0] data_52_V_read_3_reg_8928_pp0_iter13_reg;
reg   [15:0] data_52_V_read_3_reg_8928_pp0_iter14_reg;
reg   [15:0] data_51_V_read52_reg_8956;
reg   [15:0] data_51_V_read52_reg_8956_pp0_iter1_reg;
reg   [15:0] data_51_V_read52_reg_8956_pp0_iter2_reg;
reg   [15:0] data_51_V_read52_reg_8956_pp0_iter3_reg;
reg   [15:0] data_51_V_read52_reg_8956_pp0_iter4_reg;
reg   [15:0] data_51_V_read52_reg_8956_pp0_iter5_reg;
reg   [15:0] data_51_V_read52_reg_8956_pp0_iter6_reg;
reg   [15:0] data_51_V_read52_reg_8956_pp0_iter7_reg;
reg   [15:0] data_51_V_read52_reg_8956_pp0_iter8_reg;
reg   [15:0] data_51_V_read52_reg_8956_pp0_iter9_reg;
reg   [15:0] data_51_V_read52_reg_8956_pp0_iter10_reg;
reg   [15:0] data_51_V_read52_reg_8956_pp0_iter11_reg;
reg   [15:0] data_51_V_read52_reg_8956_pp0_iter12_reg;
reg   [15:0] data_51_V_read52_reg_8956_pp0_iter13_reg;
reg   [15:0] data_51_V_read52_reg_8956_pp0_iter14_reg;
reg   [15:0] data_50_V_read51_reg_8984;
reg   [15:0] data_50_V_read51_reg_8984_pp0_iter1_reg;
reg   [15:0] data_50_V_read51_reg_8984_pp0_iter2_reg;
reg   [15:0] data_50_V_read51_reg_8984_pp0_iter3_reg;
reg   [15:0] data_50_V_read51_reg_8984_pp0_iter4_reg;
reg   [15:0] data_50_V_read51_reg_8984_pp0_iter5_reg;
reg   [15:0] data_50_V_read51_reg_8984_pp0_iter6_reg;
reg   [15:0] data_50_V_read51_reg_8984_pp0_iter7_reg;
reg   [15:0] data_50_V_read51_reg_8984_pp0_iter8_reg;
reg   [15:0] data_50_V_read51_reg_8984_pp0_iter9_reg;
reg   [15:0] data_50_V_read51_reg_8984_pp0_iter10_reg;
reg   [15:0] data_50_V_read51_reg_8984_pp0_iter11_reg;
reg   [15:0] data_50_V_read51_reg_8984_pp0_iter12_reg;
reg   [15:0] data_50_V_read51_reg_8984_pp0_iter13_reg;
reg   [15:0] data_50_V_read51_reg_8984_pp0_iter14_reg;
reg   [15:0] data_49_V_read_3_reg_9012;
reg   [15:0] data_49_V_read_3_reg_9012_pp0_iter1_reg;
reg   [15:0] data_49_V_read_3_reg_9012_pp0_iter2_reg;
reg   [15:0] data_49_V_read_3_reg_9012_pp0_iter3_reg;
reg   [15:0] data_49_V_read_3_reg_9012_pp0_iter4_reg;
reg   [15:0] data_49_V_read_3_reg_9012_pp0_iter5_reg;
reg   [15:0] data_49_V_read_3_reg_9012_pp0_iter6_reg;
reg   [15:0] data_49_V_read_3_reg_9012_pp0_iter7_reg;
reg   [15:0] data_49_V_read_3_reg_9012_pp0_iter8_reg;
reg   [15:0] data_49_V_read_3_reg_9012_pp0_iter9_reg;
reg   [15:0] data_49_V_read_3_reg_9012_pp0_iter10_reg;
reg   [15:0] data_49_V_read_3_reg_9012_pp0_iter11_reg;
reg   [15:0] data_49_V_read_3_reg_9012_pp0_iter12_reg;
reg   [15:0] data_49_V_read_3_reg_9012_pp0_iter13_reg;
reg   [15:0] data_48_V_read_3_reg_9040;
reg   [15:0] data_48_V_read_3_reg_9040_pp0_iter1_reg;
reg   [15:0] data_48_V_read_3_reg_9040_pp0_iter2_reg;
reg   [15:0] data_48_V_read_3_reg_9040_pp0_iter3_reg;
reg   [15:0] data_48_V_read_3_reg_9040_pp0_iter4_reg;
reg   [15:0] data_48_V_read_3_reg_9040_pp0_iter5_reg;
reg   [15:0] data_48_V_read_3_reg_9040_pp0_iter6_reg;
reg   [15:0] data_48_V_read_3_reg_9040_pp0_iter7_reg;
reg   [15:0] data_48_V_read_3_reg_9040_pp0_iter8_reg;
reg   [15:0] data_48_V_read_3_reg_9040_pp0_iter9_reg;
reg   [15:0] data_48_V_read_3_reg_9040_pp0_iter10_reg;
reg   [15:0] data_48_V_read_3_reg_9040_pp0_iter11_reg;
reg   [15:0] data_48_V_read_3_reg_9040_pp0_iter12_reg;
reg   [15:0] data_48_V_read_3_reg_9040_pp0_iter13_reg;
reg   [15:0] data_47_V_read_3_reg_9066;
reg   [15:0] data_47_V_read_3_reg_9066_pp0_iter1_reg;
reg   [15:0] data_47_V_read_3_reg_9066_pp0_iter2_reg;
reg   [15:0] data_47_V_read_3_reg_9066_pp0_iter3_reg;
reg   [15:0] data_47_V_read_3_reg_9066_pp0_iter4_reg;
reg   [15:0] data_47_V_read_3_reg_9066_pp0_iter5_reg;
reg   [15:0] data_47_V_read_3_reg_9066_pp0_iter6_reg;
reg   [15:0] data_47_V_read_3_reg_9066_pp0_iter7_reg;
reg   [15:0] data_47_V_read_3_reg_9066_pp0_iter8_reg;
reg   [15:0] data_47_V_read_3_reg_9066_pp0_iter9_reg;
reg   [15:0] data_47_V_read_3_reg_9066_pp0_iter10_reg;
reg   [15:0] data_47_V_read_3_reg_9066_pp0_iter11_reg;
reg   [15:0] data_47_V_read_3_reg_9066_pp0_iter12_reg;
reg   [15:0] data_47_V_read_3_reg_9066_pp0_iter13_reg;
reg   [15:0] data_46_V_read_3_reg_9094;
reg   [15:0] data_46_V_read_3_reg_9094_pp0_iter1_reg;
reg   [15:0] data_46_V_read_3_reg_9094_pp0_iter2_reg;
reg   [15:0] data_46_V_read_3_reg_9094_pp0_iter3_reg;
reg   [15:0] data_46_V_read_3_reg_9094_pp0_iter4_reg;
reg   [15:0] data_46_V_read_3_reg_9094_pp0_iter5_reg;
reg   [15:0] data_46_V_read_3_reg_9094_pp0_iter6_reg;
reg   [15:0] data_46_V_read_3_reg_9094_pp0_iter7_reg;
reg   [15:0] data_46_V_read_3_reg_9094_pp0_iter8_reg;
reg   [15:0] data_46_V_read_3_reg_9094_pp0_iter9_reg;
reg   [15:0] data_46_V_read_3_reg_9094_pp0_iter10_reg;
reg   [15:0] data_46_V_read_3_reg_9094_pp0_iter11_reg;
reg   [15:0] data_46_V_read_3_reg_9094_pp0_iter12_reg;
reg   [15:0] data_46_V_read_3_reg_9094_pp0_iter13_reg;
reg   [15:0] data_45_V_read_3_reg_9125;
reg   [15:0] data_45_V_read_3_reg_9125_pp0_iter1_reg;
reg   [15:0] data_45_V_read_3_reg_9125_pp0_iter2_reg;
reg   [15:0] data_45_V_read_3_reg_9125_pp0_iter3_reg;
reg   [15:0] data_45_V_read_3_reg_9125_pp0_iter4_reg;
reg   [15:0] data_45_V_read_3_reg_9125_pp0_iter5_reg;
reg   [15:0] data_45_V_read_3_reg_9125_pp0_iter6_reg;
reg   [15:0] data_45_V_read_3_reg_9125_pp0_iter7_reg;
reg   [15:0] data_45_V_read_3_reg_9125_pp0_iter8_reg;
reg   [15:0] data_45_V_read_3_reg_9125_pp0_iter9_reg;
reg   [15:0] data_45_V_read_3_reg_9125_pp0_iter10_reg;
reg   [15:0] data_45_V_read_3_reg_9125_pp0_iter11_reg;
reg   [15:0] data_45_V_read_3_reg_9125_pp0_iter12_reg;
reg   [15:0] data_44_V_read_3_reg_9154;
reg   [15:0] data_44_V_read_3_reg_9154_pp0_iter1_reg;
reg   [15:0] data_44_V_read_3_reg_9154_pp0_iter2_reg;
reg   [15:0] data_44_V_read_3_reg_9154_pp0_iter3_reg;
reg   [15:0] data_44_V_read_3_reg_9154_pp0_iter4_reg;
reg   [15:0] data_44_V_read_3_reg_9154_pp0_iter5_reg;
reg   [15:0] data_44_V_read_3_reg_9154_pp0_iter6_reg;
reg   [15:0] data_44_V_read_3_reg_9154_pp0_iter7_reg;
reg   [15:0] data_44_V_read_3_reg_9154_pp0_iter8_reg;
reg   [15:0] data_44_V_read_3_reg_9154_pp0_iter9_reg;
reg   [15:0] data_44_V_read_3_reg_9154_pp0_iter10_reg;
reg   [15:0] data_44_V_read_3_reg_9154_pp0_iter11_reg;
reg   [15:0] data_44_V_read_3_reg_9154_pp0_iter12_reg;
reg   [15:0] data_43_V_read_3_reg_9184;
reg   [15:0] data_43_V_read_3_reg_9184_pp0_iter1_reg;
reg   [15:0] data_43_V_read_3_reg_9184_pp0_iter2_reg;
reg   [15:0] data_43_V_read_3_reg_9184_pp0_iter3_reg;
reg   [15:0] data_43_V_read_3_reg_9184_pp0_iter4_reg;
reg   [15:0] data_43_V_read_3_reg_9184_pp0_iter5_reg;
reg   [15:0] data_43_V_read_3_reg_9184_pp0_iter6_reg;
reg   [15:0] data_43_V_read_3_reg_9184_pp0_iter7_reg;
reg   [15:0] data_43_V_read_3_reg_9184_pp0_iter8_reg;
reg   [15:0] data_43_V_read_3_reg_9184_pp0_iter9_reg;
reg   [15:0] data_43_V_read_3_reg_9184_pp0_iter10_reg;
reg   [15:0] data_43_V_read_3_reg_9184_pp0_iter11_reg;
reg   [15:0] data_43_V_read_3_reg_9184_pp0_iter12_reg;
reg   [15:0] data_42_V_read_3_reg_9212;
reg   [15:0] data_42_V_read_3_reg_9212_pp0_iter1_reg;
reg   [15:0] data_42_V_read_3_reg_9212_pp0_iter2_reg;
reg   [15:0] data_42_V_read_3_reg_9212_pp0_iter3_reg;
reg   [15:0] data_42_V_read_3_reg_9212_pp0_iter4_reg;
reg   [15:0] data_42_V_read_3_reg_9212_pp0_iter5_reg;
reg   [15:0] data_42_V_read_3_reg_9212_pp0_iter6_reg;
reg   [15:0] data_42_V_read_3_reg_9212_pp0_iter7_reg;
reg   [15:0] data_42_V_read_3_reg_9212_pp0_iter8_reg;
reg   [15:0] data_42_V_read_3_reg_9212_pp0_iter9_reg;
reg   [15:0] data_42_V_read_3_reg_9212_pp0_iter10_reg;
reg   [15:0] data_42_V_read_3_reg_9212_pp0_iter11_reg;
reg   [15:0] data_42_V_read_3_reg_9212_pp0_iter12_reg;
reg   [15:0] data_41_V_read42_reg_9242;
reg   [15:0] data_41_V_read42_reg_9242_pp0_iter1_reg;
reg   [15:0] data_41_V_read42_reg_9242_pp0_iter2_reg;
reg   [15:0] data_41_V_read42_reg_9242_pp0_iter3_reg;
reg   [15:0] data_41_V_read42_reg_9242_pp0_iter4_reg;
reg   [15:0] data_41_V_read42_reg_9242_pp0_iter5_reg;
reg   [15:0] data_41_V_read42_reg_9242_pp0_iter6_reg;
reg   [15:0] data_41_V_read42_reg_9242_pp0_iter7_reg;
reg   [15:0] data_41_V_read42_reg_9242_pp0_iter8_reg;
reg   [15:0] data_41_V_read42_reg_9242_pp0_iter9_reg;
reg   [15:0] data_41_V_read42_reg_9242_pp0_iter10_reg;
reg   [15:0] data_41_V_read42_reg_9242_pp0_iter11_reg;
reg   [15:0] data_40_V_read41_reg_9272;
reg   [15:0] data_40_V_read41_reg_9272_pp0_iter1_reg;
reg   [15:0] data_40_V_read41_reg_9272_pp0_iter2_reg;
reg   [15:0] data_40_V_read41_reg_9272_pp0_iter3_reg;
reg   [15:0] data_40_V_read41_reg_9272_pp0_iter4_reg;
reg   [15:0] data_40_V_read41_reg_9272_pp0_iter5_reg;
reg   [15:0] data_40_V_read41_reg_9272_pp0_iter6_reg;
reg   [15:0] data_40_V_read41_reg_9272_pp0_iter7_reg;
reg   [15:0] data_40_V_read41_reg_9272_pp0_iter8_reg;
reg   [15:0] data_40_V_read41_reg_9272_pp0_iter9_reg;
reg   [15:0] data_40_V_read41_reg_9272_pp0_iter10_reg;
reg   [15:0] data_40_V_read41_reg_9272_pp0_iter11_reg;
reg   [15:0] data_39_V_read_3_reg_9301;
reg   [15:0] data_39_V_read_3_reg_9301_pp0_iter1_reg;
reg   [15:0] data_39_V_read_3_reg_9301_pp0_iter2_reg;
reg   [15:0] data_39_V_read_3_reg_9301_pp0_iter3_reg;
reg   [15:0] data_39_V_read_3_reg_9301_pp0_iter4_reg;
reg   [15:0] data_39_V_read_3_reg_9301_pp0_iter5_reg;
reg   [15:0] data_39_V_read_3_reg_9301_pp0_iter6_reg;
reg   [15:0] data_39_V_read_3_reg_9301_pp0_iter7_reg;
reg   [15:0] data_39_V_read_3_reg_9301_pp0_iter8_reg;
reg   [15:0] data_39_V_read_3_reg_9301_pp0_iter9_reg;
reg   [15:0] data_39_V_read_3_reg_9301_pp0_iter10_reg;
reg   [15:0] data_39_V_read_3_reg_9301_pp0_iter11_reg;
reg   [15:0] data_38_V_read_3_reg_9328;
reg   [15:0] data_38_V_read_3_reg_9328_pp0_iter1_reg;
reg   [15:0] data_38_V_read_3_reg_9328_pp0_iter2_reg;
reg   [15:0] data_38_V_read_3_reg_9328_pp0_iter3_reg;
reg   [15:0] data_38_V_read_3_reg_9328_pp0_iter4_reg;
reg   [15:0] data_38_V_read_3_reg_9328_pp0_iter5_reg;
reg   [15:0] data_38_V_read_3_reg_9328_pp0_iter6_reg;
reg   [15:0] data_38_V_read_3_reg_9328_pp0_iter7_reg;
reg   [15:0] data_38_V_read_3_reg_9328_pp0_iter8_reg;
reg   [15:0] data_38_V_read_3_reg_9328_pp0_iter9_reg;
reg   [15:0] data_38_V_read_3_reg_9328_pp0_iter10_reg;
reg   [15:0] data_38_V_read_3_reg_9328_pp0_iter11_reg;
reg   [15:0] data_37_V_read_3_reg_9353;
reg   [15:0] data_37_V_read_3_reg_9353_pp0_iter1_reg;
reg   [15:0] data_37_V_read_3_reg_9353_pp0_iter2_reg;
reg   [15:0] data_37_V_read_3_reg_9353_pp0_iter3_reg;
reg   [15:0] data_37_V_read_3_reg_9353_pp0_iter4_reg;
reg   [15:0] data_37_V_read_3_reg_9353_pp0_iter5_reg;
reg   [15:0] data_37_V_read_3_reg_9353_pp0_iter6_reg;
reg   [15:0] data_37_V_read_3_reg_9353_pp0_iter7_reg;
reg   [15:0] data_37_V_read_3_reg_9353_pp0_iter8_reg;
reg   [15:0] data_37_V_read_3_reg_9353_pp0_iter9_reg;
reg   [15:0] data_37_V_read_3_reg_9353_pp0_iter10_reg;
reg   [15:0] data_36_V_read_3_reg_9383;
reg   [15:0] data_36_V_read_3_reg_9383_pp0_iter1_reg;
reg   [15:0] data_36_V_read_3_reg_9383_pp0_iter2_reg;
reg   [15:0] data_36_V_read_3_reg_9383_pp0_iter3_reg;
reg   [15:0] data_36_V_read_3_reg_9383_pp0_iter4_reg;
reg   [15:0] data_36_V_read_3_reg_9383_pp0_iter5_reg;
reg   [15:0] data_36_V_read_3_reg_9383_pp0_iter6_reg;
reg   [15:0] data_36_V_read_3_reg_9383_pp0_iter7_reg;
reg   [15:0] data_36_V_read_3_reg_9383_pp0_iter8_reg;
reg   [15:0] data_36_V_read_3_reg_9383_pp0_iter9_reg;
reg   [15:0] data_36_V_read_3_reg_9383_pp0_iter10_reg;
reg   [15:0] data_35_V_read_3_reg_9410;
reg   [15:0] data_35_V_read_3_reg_9410_pp0_iter1_reg;
reg   [15:0] data_35_V_read_3_reg_9410_pp0_iter2_reg;
reg   [15:0] data_35_V_read_3_reg_9410_pp0_iter3_reg;
reg   [15:0] data_35_V_read_3_reg_9410_pp0_iter4_reg;
reg   [15:0] data_35_V_read_3_reg_9410_pp0_iter5_reg;
reg   [15:0] data_35_V_read_3_reg_9410_pp0_iter6_reg;
reg   [15:0] data_35_V_read_3_reg_9410_pp0_iter7_reg;
reg   [15:0] data_35_V_read_3_reg_9410_pp0_iter8_reg;
reg   [15:0] data_35_V_read_3_reg_9410_pp0_iter9_reg;
reg   [15:0] data_35_V_read_3_reg_9410_pp0_iter10_reg;
reg   [15:0] data_34_V_read_3_reg_9434;
reg   [15:0] data_34_V_read_3_reg_9434_pp0_iter1_reg;
reg   [15:0] data_34_V_read_3_reg_9434_pp0_iter2_reg;
reg   [15:0] data_34_V_read_3_reg_9434_pp0_iter3_reg;
reg   [15:0] data_34_V_read_3_reg_9434_pp0_iter4_reg;
reg   [15:0] data_34_V_read_3_reg_9434_pp0_iter5_reg;
reg   [15:0] data_34_V_read_3_reg_9434_pp0_iter6_reg;
reg   [15:0] data_34_V_read_3_reg_9434_pp0_iter7_reg;
reg   [15:0] data_34_V_read_3_reg_9434_pp0_iter8_reg;
reg   [15:0] data_34_V_read_3_reg_9434_pp0_iter9_reg;
reg   [15:0] data_34_V_read_3_reg_9434_pp0_iter10_reg;
reg   [15:0] data_33_V_read_3_reg_9463;
reg   [15:0] data_33_V_read_3_reg_9463_pp0_iter1_reg;
reg   [15:0] data_33_V_read_3_reg_9463_pp0_iter2_reg;
reg   [15:0] data_33_V_read_3_reg_9463_pp0_iter3_reg;
reg   [15:0] data_33_V_read_3_reg_9463_pp0_iter4_reg;
reg   [15:0] data_33_V_read_3_reg_9463_pp0_iter5_reg;
reg   [15:0] data_33_V_read_3_reg_9463_pp0_iter6_reg;
reg   [15:0] data_33_V_read_3_reg_9463_pp0_iter7_reg;
reg   [15:0] data_33_V_read_3_reg_9463_pp0_iter8_reg;
reg   [15:0] data_33_V_read_3_reg_9463_pp0_iter9_reg;
reg   [15:0] data_33_V_read_3_reg_9463_pp0_iter10_reg;
reg   [15:0] data_32_V_read_3_reg_9492;
reg   [15:0] data_32_V_read_3_reg_9492_pp0_iter1_reg;
reg   [15:0] data_32_V_read_3_reg_9492_pp0_iter2_reg;
reg   [15:0] data_32_V_read_3_reg_9492_pp0_iter3_reg;
reg   [15:0] data_32_V_read_3_reg_9492_pp0_iter4_reg;
reg   [15:0] data_32_V_read_3_reg_9492_pp0_iter5_reg;
reg   [15:0] data_32_V_read_3_reg_9492_pp0_iter6_reg;
reg   [15:0] data_32_V_read_3_reg_9492_pp0_iter7_reg;
reg   [15:0] data_32_V_read_3_reg_9492_pp0_iter8_reg;
reg   [15:0] data_32_V_read_3_reg_9492_pp0_iter9_reg;
reg   [15:0] data_31_V_read32_reg_9521;
reg   [15:0] data_31_V_read32_reg_9521_pp0_iter1_reg;
reg   [15:0] data_31_V_read32_reg_9521_pp0_iter2_reg;
reg   [15:0] data_31_V_read32_reg_9521_pp0_iter3_reg;
reg   [15:0] data_31_V_read32_reg_9521_pp0_iter4_reg;
reg   [15:0] data_31_V_read32_reg_9521_pp0_iter5_reg;
reg   [15:0] data_31_V_read32_reg_9521_pp0_iter6_reg;
reg   [15:0] data_31_V_read32_reg_9521_pp0_iter7_reg;
reg   [15:0] data_31_V_read32_reg_9521_pp0_iter8_reg;
reg   [15:0] data_31_V_read32_reg_9521_pp0_iter9_reg;
reg   [15:0] data_30_V_read31_reg_9549;
reg   [15:0] data_30_V_read31_reg_9549_pp0_iter1_reg;
reg   [15:0] data_30_V_read31_reg_9549_pp0_iter2_reg;
reg   [15:0] data_30_V_read31_reg_9549_pp0_iter3_reg;
reg   [15:0] data_30_V_read31_reg_9549_pp0_iter4_reg;
reg   [15:0] data_30_V_read31_reg_9549_pp0_iter5_reg;
reg   [15:0] data_30_V_read31_reg_9549_pp0_iter6_reg;
reg   [15:0] data_30_V_read31_reg_9549_pp0_iter7_reg;
reg   [15:0] data_30_V_read31_reg_9549_pp0_iter8_reg;
reg   [15:0] data_30_V_read31_reg_9549_pp0_iter9_reg;
reg   [15:0] data_29_V_read_8_reg_9573;
reg   [15:0] data_29_V_read_8_reg_9573_pp0_iter1_reg;
reg   [15:0] data_29_V_read_8_reg_9573_pp0_iter2_reg;
reg   [15:0] data_29_V_read_8_reg_9573_pp0_iter3_reg;
reg   [15:0] data_29_V_read_8_reg_9573_pp0_iter4_reg;
reg   [15:0] data_29_V_read_8_reg_9573_pp0_iter5_reg;
reg   [15:0] data_29_V_read_8_reg_9573_pp0_iter6_reg;
reg   [15:0] data_29_V_read_8_reg_9573_pp0_iter7_reg;
reg   [15:0] data_29_V_read_8_reg_9573_pp0_iter8_reg;
reg   [15:0] data_29_V_read_8_reg_9573_pp0_iter9_reg;
reg   [15:0] data_28_V_read_8_reg_9598;
reg   [15:0] data_28_V_read_8_reg_9598_pp0_iter1_reg;
reg   [15:0] data_28_V_read_8_reg_9598_pp0_iter2_reg;
reg   [15:0] data_28_V_read_8_reg_9598_pp0_iter3_reg;
reg   [15:0] data_28_V_read_8_reg_9598_pp0_iter4_reg;
reg   [15:0] data_28_V_read_8_reg_9598_pp0_iter5_reg;
reg   [15:0] data_28_V_read_8_reg_9598_pp0_iter6_reg;
reg   [15:0] data_28_V_read_8_reg_9598_pp0_iter7_reg;
reg   [15:0] data_28_V_read_8_reg_9598_pp0_iter8_reg;
reg   [15:0] data_27_V_read28_reg_9625;
reg   [15:0] data_27_V_read28_reg_9625_pp0_iter1_reg;
reg   [15:0] data_27_V_read28_reg_9625_pp0_iter2_reg;
reg   [15:0] data_27_V_read28_reg_9625_pp0_iter3_reg;
reg   [15:0] data_27_V_read28_reg_9625_pp0_iter4_reg;
reg   [15:0] data_27_V_read28_reg_9625_pp0_iter5_reg;
reg   [15:0] data_27_V_read28_reg_9625_pp0_iter6_reg;
reg   [15:0] data_27_V_read28_reg_9625_pp0_iter7_reg;
reg   [15:0] data_27_V_read28_reg_9625_pp0_iter8_reg;
reg   [15:0] data_26_V_read27_reg_9652;
reg   [15:0] data_26_V_read27_reg_9652_pp0_iter1_reg;
reg   [15:0] data_26_V_read27_reg_9652_pp0_iter2_reg;
reg   [15:0] data_26_V_read27_reg_9652_pp0_iter3_reg;
reg   [15:0] data_26_V_read27_reg_9652_pp0_iter4_reg;
reg   [15:0] data_26_V_read27_reg_9652_pp0_iter5_reg;
reg   [15:0] data_26_V_read27_reg_9652_pp0_iter6_reg;
reg   [15:0] data_26_V_read27_reg_9652_pp0_iter7_reg;
reg   [15:0] data_26_V_read27_reg_9652_pp0_iter8_reg;
reg   [15:0] data_25_V_read26_reg_9677;
reg   [15:0] data_25_V_read26_reg_9677_pp0_iter1_reg;
reg   [15:0] data_25_V_read26_reg_9677_pp0_iter2_reg;
reg   [15:0] data_25_V_read26_reg_9677_pp0_iter3_reg;
reg   [15:0] data_25_V_read26_reg_9677_pp0_iter4_reg;
reg   [15:0] data_25_V_read26_reg_9677_pp0_iter5_reg;
reg   [15:0] data_25_V_read26_reg_9677_pp0_iter6_reg;
reg   [15:0] data_25_V_read26_reg_9677_pp0_iter7_reg;
reg   [15:0] data_25_V_read26_reg_9677_pp0_iter8_reg;
reg   [15:0] data_24_V_read25_reg_9704;
reg   [15:0] data_24_V_read25_reg_9704_pp0_iter1_reg;
reg   [15:0] data_24_V_read25_reg_9704_pp0_iter2_reg;
reg   [15:0] data_24_V_read25_reg_9704_pp0_iter3_reg;
reg   [15:0] data_24_V_read25_reg_9704_pp0_iter4_reg;
reg   [15:0] data_24_V_read25_reg_9704_pp0_iter5_reg;
reg   [15:0] data_24_V_read25_reg_9704_pp0_iter6_reg;
reg   [15:0] data_24_V_read25_reg_9704_pp0_iter7_reg;
reg   [15:0] data_24_V_read25_reg_9704_pp0_iter8_reg;
reg   [15:0] data_23_V_read24_reg_9730;
reg   [15:0] data_23_V_read24_reg_9730_pp0_iter1_reg;
reg   [15:0] data_23_V_read24_reg_9730_pp0_iter2_reg;
reg   [15:0] data_23_V_read24_reg_9730_pp0_iter3_reg;
reg   [15:0] data_23_V_read24_reg_9730_pp0_iter4_reg;
reg   [15:0] data_23_V_read24_reg_9730_pp0_iter5_reg;
reg   [15:0] data_23_V_read24_reg_9730_pp0_iter6_reg;
reg   [15:0] data_23_V_read24_reg_9730_pp0_iter7_reg;
reg   [15:0] data_22_V_read23_reg_9756;
reg   [15:0] data_22_V_read23_reg_9756_pp0_iter1_reg;
reg   [15:0] data_22_V_read23_reg_9756_pp0_iter2_reg;
reg   [15:0] data_22_V_read23_reg_9756_pp0_iter3_reg;
reg   [15:0] data_22_V_read23_reg_9756_pp0_iter4_reg;
reg   [15:0] data_22_V_read23_reg_9756_pp0_iter5_reg;
reg   [15:0] data_22_V_read23_reg_9756_pp0_iter6_reg;
reg   [15:0] data_22_V_read23_reg_9756_pp0_iter7_reg;
reg   [15:0] data_22_V_read23_reg_9756_pp0_iter8_reg;
reg   [15:0] data_21_V_read22_reg_9784;
reg   [15:0] data_21_V_read22_reg_9784_pp0_iter1_reg;
reg   [15:0] data_21_V_read22_reg_9784_pp0_iter2_reg;
reg   [15:0] data_21_V_read22_reg_9784_pp0_iter3_reg;
reg   [15:0] data_21_V_read22_reg_9784_pp0_iter4_reg;
reg   [15:0] data_21_V_read22_reg_9784_pp0_iter5_reg;
reg   [15:0] data_21_V_read22_reg_9784_pp0_iter6_reg;
reg   [15:0] data_21_V_read22_reg_9784_pp0_iter7_reg;
reg   [15:0] data_20_V_read21_reg_9814;
reg   [15:0] data_20_V_read21_reg_9814_pp0_iter1_reg;
reg   [15:0] data_20_V_read21_reg_9814_pp0_iter2_reg;
reg   [15:0] data_20_V_read21_reg_9814_pp0_iter3_reg;
reg   [15:0] data_20_V_read21_reg_9814_pp0_iter4_reg;
reg   [15:0] data_20_V_read21_reg_9814_pp0_iter5_reg;
reg   [15:0] data_20_V_read21_reg_9814_pp0_iter6_reg;
reg   [15:0] data_20_V_read21_reg_9814_pp0_iter7_reg;
reg   [15:0] data_19_V_read_8_reg_9845;
reg   [15:0] data_19_V_read_8_reg_9845_pp0_iter1_reg;
reg   [15:0] data_19_V_read_8_reg_9845_pp0_iter2_reg;
reg   [15:0] data_19_V_read_8_reg_9845_pp0_iter3_reg;
reg   [15:0] data_19_V_read_8_reg_9845_pp0_iter4_reg;
reg   [15:0] data_19_V_read_8_reg_9845_pp0_iter5_reg;
reg   [15:0] data_19_V_read_8_reg_9845_pp0_iter6_reg;
reg   [15:0] data_18_V_read_8_reg_9874;
reg   [15:0] data_18_V_read_8_reg_9874_pp0_iter1_reg;
reg   [15:0] data_18_V_read_8_reg_9874_pp0_iter2_reg;
reg   [15:0] data_18_V_read_8_reg_9874_pp0_iter3_reg;
reg   [15:0] data_18_V_read_8_reg_9874_pp0_iter4_reg;
reg   [15:0] data_18_V_read_8_reg_9874_pp0_iter5_reg;
reg   [15:0] data_18_V_read_8_reg_9874_pp0_iter6_reg;
reg   [15:0] data_17_V_read18_reg_9904;
reg   [15:0] data_17_V_read18_reg_9904_pp0_iter1_reg;
reg   [15:0] data_17_V_read18_reg_9904_pp0_iter2_reg;
reg   [15:0] data_17_V_read18_reg_9904_pp0_iter3_reg;
reg   [15:0] data_17_V_read18_reg_9904_pp0_iter4_reg;
reg   [15:0] data_17_V_read18_reg_9904_pp0_iter5_reg;
reg   [15:0] data_17_V_read18_reg_9904_pp0_iter6_reg;
reg   [15:0] data_16_V_read17_reg_9935;
reg   [15:0] data_16_V_read17_reg_9935_pp0_iter1_reg;
reg   [15:0] data_16_V_read17_reg_9935_pp0_iter2_reg;
reg   [15:0] data_16_V_read17_reg_9935_pp0_iter3_reg;
reg   [15:0] data_16_V_read17_reg_9935_pp0_iter4_reg;
reg   [15:0] data_16_V_read17_reg_9935_pp0_iter5_reg;
reg   [15:0] data_16_V_read17_reg_9935_pp0_iter6_reg;
reg   [15:0] data_15_V_read16_reg_9962;
reg   [15:0] data_15_V_read16_reg_9962_pp0_iter1_reg;
reg   [15:0] data_15_V_read16_reg_9962_pp0_iter2_reg;
reg   [15:0] data_15_V_read16_reg_9962_pp0_iter3_reg;
reg   [15:0] data_15_V_read16_reg_9962_pp0_iter4_reg;
reg   [15:0] data_15_V_read16_reg_9962_pp0_iter5_reg;
reg   [15:0] data_14_V_read15_reg_9987;
reg   [15:0] data_14_V_read15_reg_9987_pp0_iter1_reg;
reg   [15:0] data_14_V_read15_reg_9987_pp0_iter2_reg;
reg   [15:0] data_14_V_read15_reg_9987_pp0_iter3_reg;
reg   [15:0] data_14_V_read15_reg_9987_pp0_iter4_reg;
reg   [15:0] data_14_V_read15_reg_9987_pp0_iter5_reg;
reg   [15:0] data_13_V_read14_reg_10015;
reg   [15:0] data_13_V_read14_reg_10015_pp0_iter1_reg;
reg   [15:0] data_13_V_read14_reg_10015_pp0_iter2_reg;
reg   [15:0] data_13_V_read14_reg_10015_pp0_iter3_reg;
reg   [15:0] data_13_V_read14_reg_10015_pp0_iter4_reg;
reg   [15:0] data_13_V_read14_reg_10015_pp0_iter5_reg;
reg   [15:0] data_12_V_read13_reg_10045;
reg   [15:0] data_12_V_read13_reg_10045_pp0_iter1_reg;
reg   [15:0] data_12_V_read13_reg_10045_pp0_iter2_reg;
reg   [15:0] data_12_V_read13_reg_10045_pp0_iter3_reg;
reg   [15:0] data_12_V_read13_reg_10045_pp0_iter4_reg;
reg   [15:0] data_12_V_read13_reg_10045_pp0_iter5_reg;
reg   [15:0] data_11_V_read12_reg_10075;
reg   [15:0] data_11_V_read12_reg_10075_pp0_iter1_reg;
reg   [15:0] data_11_V_read12_reg_10075_pp0_iter2_reg;
reg   [15:0] data_11_V_read12_reg_10075_pp0_iter3_reg;
reg   [15:0] data_11_V_read12_reg_10075_pp0_iter4_reg;
reg   [15:0] data_11_V_read12_reg_10075_pp0_iter5_reg;
reg   [15:0] data_10_V_read11_reg_10105;
reg   [15:0] data_10_V_read11_reg_10105_pp0_iter1_reg;
reg   [15:0] data_10_V_read11_reg_10105_pp0_iter2_reg;
reg   [15:0] data_10_V_read11_reg_10105_pp0_iter3_reg;
reg   [15:0] data_10_V_read11_reg_10105_pp0_iter4_reg;
reg   [15:0] data_9_V_read_8_reg_10136;
reg   [15:0] data_9_V_read_8_reg_10136_pp0_iter1_reg;
reg   [15:0] data_9_V_read_8_reg_10136_pp0_iter2_reg;
reg   [15:0] data_9_V_read_8_reg_10136_pp0_iter3_reg;
reg   [15:0] data_9_V_read_8_reg_10136_pp0_iter4_reg;
reg   [15:0] data_8_V_read_8_reg_10164;
reg   [15:0] data_8_V_read_8_reg_10164_pp0_iter1_reg;
reg   [15:0] data_8_V_read_8_reg_10164_pp0_iter2_reg;
reg   [15:0] data_8_V_read_8_reg_10164_pp0_iter3_reg;
reg   [15:0] data_8_V_read_8_reg_10164_pp0_iter4_reg;
reg   [15:0] data_7_V_read_9_reg_10191;
reg   [15:0] data_7_V_read_9_reg_10191_pp0_iter1_reg;
reg   [15:0] data_7_V_read_9_reg_10191_pp0_iter2_reg;
reg   [15:0] data_7_V_read_9_reg_10191_pp0_iter3_reg;
reg   [15:0] data_7_V_read_9_reg_10191_pp0_iter4_reg;
reg   [15:0] data_6_V_read_9_reg_10218;
reg   [15:0] data_6_V_read_9_reg_10218_pp0_iter1_reg;
reg   [15:0] data_6_V_read_9_reg_10218_pp0_iter2_reg;
reg   [15:0] data_6_V_read_9_reg_10218_pp0_iter3_reg;
reg   [15:0] data_5_V_read_9_reg_10245;
reg   [15:0] data_5_V_read_9_reg_10245_pp0_iter1_reg;
reg   [15:0] data_5_V_read_9_reg_10245_pp0_iter2_reg;
reg   [15:0] data_5_V_read_9_reg_10245_pp0_iter3_reg;
reg   [15:0] data_4_V_read_10_reg_10273;
reg   [15:0] data_4_V_read_10_reg_10273_pp0_iter1_reg;
reg   [15:0] data_4_V_read_10_reg_10273_pp0_iter2_reg;
reg   [15:0] data_4_V_read_10_reg_10273_pp0_iter3_reg;
reg   [15:0] data_3_V_read_10_reg_10295;
reg   [15:0] data_3_V_read_10_reg_10295_pp0_iter1_reg;
reg   [15:0] data_3_V_read_10_reg_10295_pp0_iter2_reg;
reg   [15:0] data_2_V_read_10_reg_10312;
reg   [15:0] data_2_V_read_10_reg_10312_pp0_iter1_reg;
reg   [15:0] data_1_V_read_10_reg_10323;
reg   [15:0] data_0_V_read_10_reg_10329;
wire   [15:0] add_ln703_fu_530_p2;
reg   [15:0] add_ln703_reg_10335;
reg   [15:0] add_ln703_reg_10335_pp0_iter1_reg;
wire   [15:0] sub_ln703_fu_536_p2;
reg   [15:0] sub_ln703_reg_10342;
wire   [15:0] sub_ln703_1_fu_540_p2;
reg   [15:0] sub_ln703_1_reg_10348;
wire   [15:0] add_ln703_131_fu_544_p2;
reg   [15:0] add_ln703_131_reg_10354;
reg   [15:0] add_ln703_131_reg_10354_pp0_iter2_reg;
wire   [15:0] sub_ln703_4_fu_548_p2;
reg   [15:0] sub_ln703_4_reg_10361;
reg   [15:0] sub_ln703_4_reg_10361_pp0_iter2_reg;
wire   [15:0] sub_ln703_2_fu_552_p2;
reg   [15:0] sub_ln703_2_reg_10367;
wire   [15:0] add_ln703_130_fu_556_p2;
reg   [15:0] add_ln703_130_reg_10373;
wire   [15:0] sub_ln703_3_fu_560_p2;
reg   [15:0] sub_ln703_3_reg_10379;
wire   [15:0] add_ln703_134_fu_568_p2;
reg   [15:0] add_ln703_134_reg_10385;
wire   [15:0] sub_ln703_8_fu_572_p2;
reg   [15:0] sub_ln703_8_reg_10392;
wire   [15:0] sub_ln703_11_fu_576_p2;
reg   [15:0] sub_ln703_11_reg_10398;
reg   [15:0] sub_ln703_11_reg_10398_pp0_iter3_reg;
wire   [15:0] add_ln703_144_fu_589_p2;
reg   [15:0] add_ln703_144_reg_10403;
reg   [15:0] add_ln703_144_reg_10403_pp0_iter3_reg;
wire   [15:0] sub_ln703_6_fu_595_p2;
reg   [15:0] sub_ln703_6_reg_10408;
wire   [15:0] add_ln703_132_fu_599_p2;
reg   [15:0] add_ln703_132_reg_10414;
wire   [15:0] sub_ln703_10_fu_615_p2;
reg   [15:0] sub_ln703_10_reg_10420;
wire   [15:0] add_ln703_135_fu_619_p2;
reg   [15:0] add_ln703_135_reg_10425;
wire   [15:0] sub_ln703_15_fu_631_p2;
reg   [15:0] sub_ln703_15_reg_10430;
wire   [15:0] sub_ln703_16_fu_640_p2;
reg   [15:0] sub_ln703_16_reg_10436;
wire   [15:0] add_ln703_140_fu_644_p2;
reg   [15:0] add_ln703_140_reg_10442;
wire   [15:0] add_ln703_141_fu_649_p2;
reg   [15:0] add_ln703_141_reg_10447;
wire   [15:0] sub_ln703_17_fu_653_p2;
reg   [15:0] sub_ln703_17_reg_10453;
wire   [15:0] sub_ln703_18_fu_658_p2;
reg   [15:0] sub_ln703_18_reg_10459;
wire   [15:0] sub_ln703_20_fu_662_p2;
reg   [15:0] sub_ln703_20_reg_10465;
wire   [15:0] sub_ln703_23_fu_666_p2;
reg   [15:0] sub_ln703_23_reg_10471;
wire   [15:0] sub_ln703_28_fu_671_p2;
reg   [15:0] sub_ln703_28_reg_10476;
wire   [15:0] add_ln703_158_fu_676_p2;
reg   [15:0] add_ln703_158_reg_10482;
wire   [15:0] add_ln703_161_fu_681_p2;
reg   [15:0] add_ln703_161_reg_10487;
wire   [15:0] add_ln703_179_fu_685_p2;
reg   [15:0] add_ln703_179_reg_10495;
wire   [15:0] add_ln703_153_fu_809_p2;
reg   [15:0] add_ln703_153_reg_10503;
wire   [15:0] sub_ln703_38_fu_814_p2;
reg   [15:0] sub_ln703_38_reg_10508;
wire   [15:0] sub_ln703_39_fu_819_p2;
reg   [15:0] sub_ln703_39_reg_10513;
wire   [15:0] sub_ln703_40_fu_824_p2;
reg   [15:0] sub_ln703_40_reg_10519;
wire   [15:0] sub_ln703_43_fu_838_p2;
reg   [15:0] sub_ln703_43_reg_10524;
wire   [15:0] add_ln703_157_fu_892_p2;
reg   [15:0] add_ln703_157_reg_10529;
wire   [15:0] sub_ln703_53_fu_912_p2;
reg   [15:0] sub_ln703_53_reg_10534;
wire   [15:0] add_ln703_162_fu_917_p2;
reg   [15:0] add_ln703_162_reg_10539;
wire   [15:0] sub_ln703_58_fu_922_p2;
reg   [15:0] sub_ln703_58_reg_10545;
wire   [15:0] sub_ln703_62_fu_942_p2;
reg   [15:0] sub_ln703_62_reg_10550;
wire   [15:0] sub_ln703_63_fu_947_p2;
reg   [15:0] sub_ln703_63_reg_10555;
wire   [15:0] sub_ln703_64_fu_957_p2;
reg   [15:0] sub_ln703_64_reg_10560;
wire   [15:0] add_ln703_170_fu_972_p2;
reg   [15:0] add_ln703_170_reg_10566;
wire   [15:0] add_ln703_171_fu_977_p2;
reg   [15:0] add_ln703_171_reg_10571;
wire   [15:0] add_ln703_173_fu_982_p2;
reg   [15:0] add_ln703_173_reg_10576;
wire   [15:0] sub_ln703_66_fu_987_p2;
reg   [15:0] sub_ln703_66_reg_10581;
wire   [15:0] sub_ln703_70_fu_992_p2;
reg   [15:0] sub_ln703_70_reg_10586;
wire   [15:0] add_ln703_177_fu_997_p2;
reg   [15:0] add_ln703_177_reg_10591;
wire   [15:0] sub_ln703_71_fu_1002_p2;
reg   [15:0] sub_ln703_71_reg_10596;
wire   [15:0] add_ln703_181_fu_1015_p2;
reg   [15:0] add_ln703_181_reg_10601;
wire   [15:0] add_ln703_183_fu_1021_p2;
reg   [15:0] add_ln703_183_reg_10606;
wire   [15:0] sub_ln703_73_fu_1026_p2;
reg   [15:0] sub_ln703_73_reg_10611;
wire   [15:0] sub_ln703_75_fu_1031_p2;
reg   [15:0] sub_ln703_75_reg_10616;
wire   [15:0] add_ln703_186_fu_1036_p2;
reg   [15:0] add_ln703_186_reg_10621;
wire   [15:0] add_ln703_192_fu_1050_p2;
reg   [15:0] add_ln703_192_reg_10626;
wire   [15:0] sub_ln703_92_fu_1054_p2;
reg   [15:0] sub_ln703_92_reg_10636;
wire   [15:0] add_ln703_204_fu_1059_p2;
reg   [15:0] add_ln703_204_reg_10641;
wire   [15:0] add_ln703_209_fu_1064_p2;
reg   [15:0] add_ln703_209_reg_10646;
wire   [15:0] add_ln703_213_fu_1068_p2;
reg   [15:0] add_ln703_213_reg_10653;
wire   [15:0] add_ln703_223_fu_1073_p2;
reg   [15:0] add_ln703_223_reg_10658;
wire   [15:0] add_ln703_252_fu_1077_p2;
reg   [15:0] add_ln703_252_reg_10665;
reg   [15:0] add_ln703_252_reg_10665_pp0_iter5_reg;
wire   [15:0] add_ln703_254_fu_1081_p2;
reg   [15:0] add_ln703_254_reg_10672;
wire   [15:0] sub_ln703_96_fu_1294_p2;
reg   [15:0] sub_ln703_96_reg_10677;
wire   [15:0] add_ln703_207_fu_1299_p2;
reg   [15:0] add_ln703_207_reg_10682;
wire   [15:0] add_ln703_208_fu_1309_p2;
reg   [15:0] add_ln703_208_reg_10687;
wire   [15:0] add_ln703_210_fu_1314_p2;
reg   [15:0] add_ln703_210_reg_10692;
wire   [15:0] sub_ln703_98_fu_1319_p2;
reg   [15:0] sub_ln703_98_reg_10697;
wire   [15:0] add_ln703_216_fu_1358_p2;
reg   [15:0] add_ln703_216_reg_10702;
wire   [15:0] sub_ln703_106_fu_1378_p2;
reg   [15:0] sub_ln703_106_reg_10707;
wire   [15:0] sub_ln703_107_fu_1383_p2;
reg   [15:0] sub_ln703_107_reg_10712;
wire   [15:0] sub_ln703_108_fu_1388_p2;
reg   [15:0] sub_ln703_108_reg_10717;
wire   [15:0] sub_ln703_109_fu_1407_p2;
reg   [15:0] sub_ln703_109_reg_10722;
wire   [15:0] sub_ln703_115_fu_1432_p2;
reg   [15:0] sub_ln703_115_reg_10727;
wire   [15:0] add_ln703_224_fu_1437_p2;
reg   [15:0] add_ln703_224_reg_10732;
wire   [15:0] add_ln703_226_fu_1457_p2;
reg   [15:0] add_ln703_226_reg_10737;
wire   [15:0] sub_ln703_122_fu_1462_p2;
reg   [15:0] sub_ln703_122_reg_10742;
wire   [15:0] sub_ln703_123_fu_1467_p2;
reg   [15:0] sub_ln703_123_reg_10747;
wire   [15:0] add_ln703_227_fu_1472_p2;
reg   [15:0] add_ln703_227_reg_10752;
wire   [15:0] sub_ln703_125_fu_1482_p2;
reg   [15:0] sub_ln703_125_reg_10757;
wire   [15:0] sub_ln703_128_fu_1496_p2;
reg   [15:0] sub_ln703_128_reg_10762;
wire   [15:0] add_ln703_233_fu_1501_p2;
reg   [15:0] add_ln703_233_reg_10767;
wire   [15:0] add_ln703_236_fu_1511_p2;
reg   [15:0] add_ln703_236_reg_10772;
wire   [15:0] add_ln703_238_fu_1520_p2;
reg   [15:0] add_ln703_238_reg_10777;
wire   [15:0] sub_ln703_133_fu_1532_p2;
reg   [15:0] sub_ln703_133_reg_10782;
wire   [15:0] sub_ln703_137_fu_1548_p2;
reg   [15:0] sub_ln703_137_reg_10787;
wire   [15:0] sub_ln703_141_fu_1553_p2;
reg   [15:0] sub_ln703_141_reg_10792;
wire   [15:0] sub_ln703_142_fu_1558_p2;
reg   [15:0] sub_ln703_142_reg_10797;
wire   [15:0] add_ln703_247_fu_1563_p2;
reg   [15:0] add_ln703_247_reg_10802;
wire   [15:0] add_ln703_250_fu_1574_p2;
reg   [15:0] add_ln703_250_reg_10807;
wire   [15:0] sub_ln703_146_fu_1580_p2;
reg   [15:0] sub_ln703_146_reg_10812;
wire   [15:0] add_ln703_260_fu_1593_p2;
reg   [15:0] add_ln703_260_reg_10817;
wire   [15:0] sub_ln703_152_fu_1599_p2;
reg   [15:0] sub_ln703_152_reg_10822;
wire   [15:0] add_ln703_262_fu_1604_p2;
reg   [15:0] add_ln703_262_reg_10827;
wire   [15:0] sub_ln703_154_fu_1609_p2;
reg   [15:0] sub_ln703_154_reg_10832;
wire   [15:0] add_ln703_265_fu_1614_p2;
reg   [15:0] add_ln703_265_reg_10837;
wire   [15:0] add_ln703_280_fu_1618_p2;
reg   [15:0] add_ln703_280_reg_10846;
wire   [15:0] add_ln703_326_fu_1622_p2;
reg   [15:0] add_ln703_326_reg_10855;
reg   [15:0] add_ln703_326_reg_10855_pp0_iter6_reg;
wire   [15:0] sub_ln703_166_fu_1834_p2;
reg   [15:0] sub_ln703_166_reg_10863;
wire   [15:0] sub_ln703_183_fu_1959_p2;
reg   [15:0] sub_ln703_183_reg_10868;
wire   [15:0] add_ln703_283_fu_1979_p2;
reg   [15:0] add_ln703_283_reg_10873;
wire   [15:0] sub_ln703_184_fu_1984_p2;
reg   [15:0] sub_ln703_184_reg_10878;
wire   [15:0] sub_ln703_186_fu_1994_p2;
reg   [15:0] sub_ln703_186_reg_10883;
wire   [15:0] add_ln703_285_fu_2009_p2;
reg   [15:0] add_ln703_285_reg_10888;
wire   [15:0] sub_ln703_191_fu_2029_p2;
reg   [15:0] sub_ln703_191_reg_10893;
wire   [15:0] add_ln703_289_fu_2034_p2;
reg   [15:0] add_ln703_289_reg_10898;
wire   [15:0] add_ln703_290_fu_2039_p2;
reg   [15:0] add_ln703_290_reg_10903;
wire   [15:0] sub_ln703_194_fu_2054_p2;
reg   [15:0] sub_ln703_194_reg_10908;
wire   [15:0] sub_ln703_196_fu_2074_p2;
reg   [15:0] sub_ln703_196_reg_10913;
wire   [15:0] add_ln703_294_fu_2084_p2;
reg   [15:0] add_ln703_294_reg_10918;
wire   [15:0] add_ln703_295_fu_2089_p2;
reg   [15:0] add_ln703_295_reg_10923;
wire   [15:0] add_ln703_300_fu_2093_p2;
reg   [15:0] add_ln703_300_reg_10930;
wire   [15:0] sub_ln703_198_fu_2099_p2;
reg   [15:0] sub_ln703_198_reg_10935;
wire   [15:0] add_ln703_303_fu_2104_p2;
reg   [15:0] add_ln703_303_reg_10940;
wire   [15:0] add_ln703_304_fu_2110_p2;
reg   [15:0] add_ln703_304_reg_10945;
wire   [15:0] sub_ln703_200_fu_2115_p2;
reg   [15:0] sub_ln703_200_reg_10950;
wire   [15:0] sub_ln703_202_fu_2120_p2;
reg   [15:0] sub_ln703_202_reg_10955;
wire   [15:0] add_ln703_307_fu_2125_p2;
reg   [15:0] add_ln703_307_reg_10960;
wire   [15:0] sub_ln703_203_fu_2131_p2;
reg   [15:0] sub_ln703_203_reg_10965;
wire   [15:0] add_ln703_309_fu_2136_p2;
reg   [15:0] add_ln703_309_reg_10970;
wire   [15:0] sub_ln703_204_fu_2142_p2;
reg   [15:0] sub_ln703_204_reg_10975;
wire   [15:0] add_ln703_310_fu_2147_p2;
reg   [15:0] add_ln703_310_reg_10980;
wire   [15:0] sub_ln703_208_fu_2152_p2;
reg   [15:0] sub_ln703_208_reg_10985;
wire   [15:0] sub_ln703_209_fu_2157_p2;
reg   [15:0] sub_ln703_209_reg_10990;
wire   [15:0] sub_ln703_210_fu_2162_p2;
reg   [15:0] sub_ln703_210_reg_10995;
wire   [15:0] sub_ln703_212_fu_2173_p2;
reg   [15:0] sub_ln703_212_reg_11000;
wire   [15:0] add_ln703_323_fu_2188_p2;
reg   [15:0] add_ln703_323_reg_11005;
wire   [15:0] sub_ln703_230_fu_2194_p2;
reg   [15:0] sub_ln703_230_reg_11010;
wire   [15:0] add_ln703_328_fu_2208_p2;
reg   [15:0] add_ln703_328_reg_11015;
wire   [15:0] sub_ln703_237_fu_2214_p2;
reg   [15:0] sub_ln703_237_reg_11020;
wire   [15:0] add_ln703_333_fu_2224_p2;
reg   [15:0] add_ln703_333_reg_11025;
wire   [15:0] add_ln703_341_fu_2230_p2;
reg   [15:0] add_ln703_341_reg_11030;
wire   [15:0] add_ln703_369_fu_2234_p2;
reg   [15:0] add_ln703_369_reg_11037;
reg   [15:0] add_ln703_369_reg_11037_pp0_iter7_reg;
wire   [15:0] sub_ln703_234_fu_2395_p2;
reg   [15:0] sub_ln703_234_reg_11046;
wire   [15:0] sub_ln703_246_fu_2477_p2;
reg   [15:0] sub_ln703_246_reg_11051;
wire   [15:0] sub_ln703_249_fu_2496_p2;
reg   [15:0] sub_ln703_249_reg_11056;
wire   [15:0] sub_ln703_250_fu_2501_p2;
reg   [15:0] sub_ln703_250_reg_11061;
wire   [15:0] sub_ln703_251_fu_2506_p2;
reg   [15:0] sub_ln703_251_reg_11066;
wire   [15:0] add_ln703_342_fu_2520_p2;
reg   [15:0] add_ln703_342_reg_11071;
wire   [15:0] sub_ln703_254_fu_2525_p2;
reg   [15:0] sub_ln703_254_reg_11076;
wire   [15:0] sub_ln703_256_fu_2534_p2;
reg   [15:0] sub_ln703_256_reg_11081;
wire   [15:0] sub_ln703_257_fu_2539_p2;
reg   [15:0] sub_ln703_257_reg_11086;
wire   [15:0] sub_ln703_261_fu_2569_p2;
reg   [15:0] sub_ln703_261_reg_11091;
wire   [15:0] sub_ln703_262_fu_2574_p2;
reg   [15:0] sub_ln703_262_reg_11096;
wire   [15:0] sub_ln703_263_fu_2579_p2;
reg   [15:0] sub_ln703_263_reg_11101;
wire   [15:0] add_ln703_346_fu_2589_p2;
reg   [15:0] add_ln703_346_reg_11106;
wire   [15:0] add_ln703_350_fu_2602_p2;
reg   [15:0] add_ln703_350_reg_11111;
wire   [15:0] sub_ln703_265_fu_2613_p2;
reg   [15:0] sub_ln703_265_reg_11116;
wire   [15:0] sub_ln703_270_fu_2628_p2;
reg   [15:0] sub_ln703_270_reg_11121;
wire   [15:0] add_ln703_352_fu_2633_p2;
reg   [15:0] add_ln703_352_reg_11126;
wire   [15:0] add_ln703_354_fu_2638_p2;
reg   [15:0] add_ln703_354_reg_11131;
wire   [15:0] sub_ln703_272_fu_2647_p2;
reg   [15:0] sub_ln703_272_reg_11138;
wire   [15:0] sub_ln703_274_fu_2652_p2;
reg   [15:0] sub_ln703_274_reg_11143;
wire   [15:0] add_ln703_356_fu_2657_p2;
reg   [15:0] add_ln703_356_reg_11148;
wire   [15:0] sub_ln703_275_fu_2662_p2;
reg   [15:0] sub_ln703_275_reg_11153;
wire   [15:0] add_ln703_360_fu_2677_p2;
reg   [15:0] add_ln703_360_reg_11158;
wire   [15:0] sub_ln703_281_fu_2688_p2;
reg   [15:0] sub_ln703_281_reg_11163;
wire   [15:0] sub_ln703_284_fu_2698_p2;
reg   [15:0] sub_ln703_284_reg_11168;
wire   [15:0] sub_ln703_289_fu_2703_p2;
reg   [15:0] sub_ln703_289_reg_11173;
wire   [15:0] sub_ln703_293_fu_2708_p2;
reg   [15:0] sub_ln703_293_reg_11178;
wire   [15:0] sub_ln703_296_fu_2713_p2;
reg   [15:0] sub_ln703_296_reg_11183;
wire   [15:0] sub_ln703_301_fu_2718_p2;
reg   [15:0] sub_ln703_301_reg_11188;
wire   [15:0] add_ln703_371_fu_2732_p2;
reg   [15:0] add_ln703_371_reg_11193;
wire   [15:0] add_ln703_375_fu_2738_p2;
reg   [15:0] add_ln703_375_reg_11198;
wire   [15:0] add_ln703_384_fu_2743_p2;
reg   [15:0] add_ln703_384_reg_11203;
wire   [15:0] add_ln703_400_fu_2752_p2;
reg   [15:0] add_ln703_400_reg_11210;
wire   [15:0] add_ln703_402_fu_2758_p2;
reg   [15:0] add_ln703_402_reg_11215;
reg   [15:0] add_ln703_402_reg_11215_pp0_iter8_reg;
wire   [15:0] add_ln703_424_fu_2762_p2;
reg   [15:0] add_ln703_424_reg_11225;
wire   [15:0] add_ln703_439_fu_2766_p2;
reg   [15:0] add_ln703_439_reg_11233;
reg   [15:0] add_ln703_439_reg_11233_pp0_iter8_reg;
wire   [15:0] add_ln703_525_fu_2774_p2;
reg   [15:0] add_ln703_525_reg_11243;
reg   [15:0] add_ln703_525_reg_11243_pp0_iter8_reg;
reg   [15:0] add_ln703_525_reg_11243_pp0_iter9_reg;
wire   [15:0] add_ln703_534_fu_2779_p2;
reg   [15:0] add_ln703_534_reg_11248;
reg   [15:0] add_ln703_534_reg_11248_pp0_iter8_reg;
reg   [15:0] add_ln703_534_reg_11248_pp0_iter9_reg;
wire   [15:0] sub_ln703_313_fu_2998_p2;
reg   [15:0] sub_ln703_313_reg_11257;
wire   [15:0] add_ln703_386_fu_3015_p2;
reg   [15:0] add_ln703_386_reg_11262;
wire   [15:0] sub_ln703_315_fu_3021_p2;
reg   [15:0] sub_ln703_315_reg_11267;
wire   [15:0] add_ln703_390_fu_3050_p2;
reg   [15:0] add_ln703_390_reg_11272;
wire   [15:0] sub_ln703_326_fu_3101_p2;
reg   [15:0] sub_ln703_326_reg_11277;
wire   [15:0] sub_ln703_328_fu_3111_p2;
reg   [15:0] sub_ln703_328_reg_11282;
wire   [15:0] add_ln703_410_fu_3149_p2;
reg   [15:0] add_ln703_410_reg_11287;
wire   [15:0] sub_ln703_333_fu_3155_p2;
reg   [15:0] sub_ln703_333_reg_11292;
wire   [15:0] add_ln703_416_fu_3170_p2;
reg   [15:0] add_ln703_416_reg_11297;
wire   [15:0] sub_ln703_334_fu_3175_p2;
reg   [15:0] sub_ln703_334_reg_11302;
wire   [15:0] sub_ln703_336_fu_3180_p2;
reg   [15:0] sub_ln703_336_reg_11307;
wire   [15:0] add_ln703_417_fu_3185_p2;
reg   [15:0] add_ln703_417_reg_11312;
wire   [15:0] sub_ln703_339_fu_3200_p2;
reg   [15:0] sub_ln703_339_reg_11317;
wire   [15:0] sub_ln703_340_fu_3205_p2;
reg   [15:0] sub_ln703_340_reg_11322;
wire   [15:0] sub_ln703_342_fu_3215_p2;
reg   [15:0] sub_ln703_342_reg_11327;
wire   [15:0] sub_ln703_344_fu_3220_p2;
reg   [15:0] sub_ln703_344_reg_11332;
wire   [15:0] sub_ln703_345_fu_3234_p2;
reg   [15:0] sub_ln703_345_reg_11337;
wire   [15:0] sub_ln703_350_fu_3244_p2;
reg   [15:0] sub_ln703_350_reg_11342;
wire   [15:0] add_ln703_426_fu_3258_p2;
reg   [15:0] add_ln703_426_reg_11347;
wire   [15:0] sub_ln703_353_fu_3269_p2;
reg   [15:0] sub_ln703_353_reg_11352;
wire   [15:0] add_ln703_431_fu_3274_p2;
reg   [15:0] add_ln703_431_reg_11357;
wire   [15:0] add_ln703_435_fu_3284_p2;
reg   [15:0] add_ln703_435_reg_11362;
wire   [15:0] sub_ln703_356_fu_3290_p2;
reg   [15:0] sub_ln703_356_reg_11367;
wire   [15:0] sub_ln703_358_fu_3300_p2;
reg   [15:0] sub_ln703_358_reg_11372;
wire   [15:0] sub_ln703_362_fu_3305_p2;
reg   [15:0] sub_ln703_362_reg_11377;
wire   [15:0] add_ln703_438_fu_3310_p2;
reg   [15:0] add_ln703_438_reg_11382;
wire   [15:0] add_ln703_445_fu_3315_p2;
reg   [15:0] add_ln703_445_reg_11387;
wire   [15:0] add_ln703_447_fu_3320_p2;
reg   [15:0] add_ln703_447_reg_11392;
wire   [15:0] sub_ln703_371_fu_3324_p2;
reg   [15:0] sub_ln703_371_reg_11397;
wire   [15:0] add_ln703_451_fu_3329_p2;
reg   [15:0] add_ln703_451_reg_11402;
wire   [15:0] add_ln703_466_fu_3333_p2;
reg   [15:0] add_ln703_466_reg_11410;
wire   [15:0] add_ln703_471_fu_3337_p2;
reg   [15:0] add_ln703_471_reg_11418;
wire   [15:0] add_ln703_484_fu_3342_p2;
reg   [15:0] add_ln703_484_reg_11423;
wire   [15:0] add_ln703_490_fu_3347_p2;
reg   [15:0] add_ln703_490_reg_11428;
wire   [15:0] add_ln703_498_fu_3351_p2;
reg   [15:0] add_ln703_498_reg_11436;
wire   [15:0] add_ln703_507_fu_3356_p2;
reg   [15:0] add_ln703_507_reg_11441;
reg   [15:0] add_ln703_507_reg_11441_pp0_iter9_reg;
wire   [15:0] add_ln703_528_fu_3360_p2;
reg   [15:0] add_ln703_528_reg_11452;
reg   [15:0] add_ln703_528_reg_11452_pp0_iter9_reg;
wire   [15:0] add_ln703_535_fu_3364_p2;
reg   [15:0] add_ln703_535_reg_11457;
wire   [15:0] add_ln703_568_fu_3368_p2;
reg   [15:0] add_ln703_568_reg_11464;
reg   [15:0] add_ln703_568_reg_11464_pp0_iter9_reg;
wire   [15:0] sub_ln703_384_fu_3645_p2;
reg   [15:0] sub_ln703_384_reg_11474;
wire   [15:0] add_ln703_469_fu_3655_p2;
reg   [15:0] add_ln703_469_reg_11479;
wire   [15:0] sub_ln703_386_fu_3660_p2;
reg   [15:0] sub_ln703_386_reg_11484;
wire   [15:0] sub_ln703_387_fu_3665_p2;
reg   [15:0] sub_ln703_387_reg_11489;
wire   [15:0] add_ln703_476_fu_3685_p2;
reg   [15:0] add_ln703_476_reg_11494;
wire   [15:0] sub_ln703_390_fu_3690_p2;
reg   [15:0] sub_ln703_390_reg_11499;
wire   [15:0] sub_ln703_393_fu_3705_p2;
reg   [15:0] sub_ln703_393_reg_11504;
wire   [15:0] sub_ln703_394_fu_3710_p2;
reg   [15:0] sub_ln703_394_reg_11509;
wire   [15:0] sub_ln703_395_fu_3720_p2;
reg   [15:0] sub_ln703_395_reg_11514;
wire   [15:0] add_ln703_478_fu_3730_p2;
reg   [15:0] add_ln703_478_reg_11519;
wire   [15:0] sub_ln703_399_fu_3761_p2;
reg   [15:0] sub_ln703_399_reg_11524;
wire   [15:0] sub_ln703_401_fu_3781_p2;
reg   [15:0] sub_ln703_401_reg_11529;
wire   [15:0] sub_ln703_402_fu_3786_p2;
reg   [15:0] sub_ln703_402_reg_11534;
wire   [15:0] sub_ln703_403_fu_3791_p2;
reg   [15:0] sub_ln703_403_reg_11539;
wire   [15:0] add_ln703_496_fu_3806_p2;
reg   [15:0] add_ln703_496_reg_11544;
wire   [15:0] add_ln703_497_fu_3811_p2;
reg   [15:0] add_ln703_497_reg_11549;
wire   [15:0] sub_ln703_405_fu_3816_p2;
reg   [15:0] sub_ln703_405_reg_11554;
wire   [15:0] add_ln703_506_fu_3839_p2;
reg   [15:0] add_ln703_506_reg_11559;
wire   [15:0] sub_ln703_408_fu_3845_p2;
reg   [15:0] sub_ln703_408_reg_11564;
wire   [15:0] sub_ln703_411_fu_3850_p2;
reg   [15:0] sub_ln703_411_reg_11569;
wire   [15:0] sub_ln703_412_fu_3855_p2;
reg   [15:0] sub_ln703_412_reg_11574;
wire   [15:0] sub_ln703_414_fu_3860_p2;
reg   [15:0] sub_ln703_414_reg_11579;
wire   [15:0] sub_ln703_416_fu_3865_p2;
reg   [15:0] sub_ln703_416_reg_11584;
wire   [15:0] add_ln703_512_fu_3878_p2;
reg   [15:0] add_ln703_512_reg_11589;
wire   [15:0] sub_ln703_419_fu_3884_p2;
reg   [15:0] sub_ln703_419_reg_11594;
wire   [15:0] add_ln703_515_fu_3889_p2;
reg   [15:0] add_ln703_515_reg_11599;
wire   [15:0] add_ln703_517_fu_3894_p2;
reg   [15:0] add_ln703_517_reg_11604;
wire   [15:0] add_ln703_537_fu_3912_p2;
reg   [15:0] add_ln703_537_reg_11609;
wire   [15:0] add_ln703_545_fu_3923_p2;
reg   [15:0] add_ln703_545_reg_11614;
wire   [15:0] add_ln703_556_fu_3933_p2;
reg   [15:0] add_ln703_556_reg_11619;
wire   [15:0] sub_ln703_440_fu_3938_p2;
reg   [15:0] sub_ln703_440_reg_11624;
wire   [15:0] add_ln703_560_fu_3943_p2;
reg   [15:0] add_ln703_560_reg_11629;
wire   [15:0] add_ln703_566_fu_3952_p2;
reg   [15:0] add_ln703_566_reg_11635;
wire   [15:0] add_ln703_569_fu_3957_p2;
reg   [15:0] add_ln703_569_reg_11640;
wire   [15:0] add_ln703_588_fu_3961_p2;
reg   [15:0] add_ln703_588_reg_11646;
wire   [15:0] add_ln703_600_fu_3965_p2;
reg   [15:0] add_ln703_600_reg_11652;
reg   [15:0] add_ln703_600_reg_11652_pp0_iter10_reg;
wire   [15:0] add_ln703_621_fu_3969_p2;
reg   [15:0] add_ln703_621_reg_11662;
reg   [15:0] add_ln703_621_reg_11662_pp0_iter10_reg;
wire   [15:0] sub_ln703_448_fu_4206_p2;
reg   [15:0] sub_ln703_448_reg_11673;
wire   [15:0] sub_ln703_452_fu_4231_p2;
reg   [15:0] sub_ln703_452_reg_11678;
wire   [15:0] sub_ln703_453_fu_4236_p2;
reg   [15:0] sub_ln703_453_reg_11683;
wire   [15:0] sub_ln703_458_fu_4270_p2;
reg   [15:0] sub_ln703_458_reg_11688;
wire   [15:0] sub_ln703_461_fu_4303_p2;
reg   [15:0] sub_ln703_461_reg_11693;
wire   [15:0] add_ln703_572_fu_4308_p2;
reg   [15:0] add_ln703_572_reg_11698;
wire   [15:0] sub_ln703_462_fu_4313_p2;
reg   [15:0] sub_ln703_462_reg_11703;
wire   [15:0] add_ln703_573_fu_4323_p2;
reg   [15:0] add_ln703_573_reg_11708;
wire   [15:0] sub_ln703_467_fu_4333_p2;
reg   [15:0] sub_ln703_467_reg_11713;
wire   [15:0] sub_ln703_468_fu_4353_p2;
reg   [15:0] sub_ln703_468_reg_11718;
wire   [15:0] add_ln703_581_fu_4358_p2;
reg   [15:0] add_ln703_581_reg_11723;
wire   [15:0] add_ln703_583_fu_4363_p2;
reg   [15:0] add_ln703_583_reg_11728;
wire   [15:0] sub_ln703_469_fu_4368_p2;
reg   [15:0] sub_ln703_469_reg_11733;
wire   [15:0] sub_ln703_470_fu_4373_p2;
reg   [15:0] sub_ln703_470_reg_11738;
wire   [15:0] add_ln703_586_fu_4398_p2;
reg   [15:0] add_ln703_586_reg_11743;
wire   [15:0] add_ln703_590_fu_4412_p2;
reg   [15:0] add_ln703_590_reg_11748;
wire   [15:0] sub_ln703_475_fu_4418_p2;
reg   [15:0] sub_ln703_475_reg_11753;
wire   [15:0] add_ln703_591_fu_4423_p2;
reg   [15:0] add_ln703_591_reg_11758;
wire   [15:0] add_ln703_592_fu_4428_p2;
reg   [15:0] add_ln703_592_reg_11763;
wire   [15:0] add_ln703_598_fu_4441_p2;
reg   [15:0] add_ln703_598_reg_11768;
wire   [15:0] sub_ln703_482_fu_4447_p2;
reg   [15:0] sub_ln703_482_reg_11773;
wire   [15:0] sub_ln703_483_fu_4452_p2;
reg   [15:0] sub_ln703_483_reg_11778;
wire   [15:0] sub_ln703_488_fu_4457_p2;
reg   [15:0] sub_ln703_488_reg_11783;
wire   [15:0] sub_ln703_490_fu_4462_p2;
reg   [15:0] sub_ln703_490_reg_11788;
wire   [15:0] sub_ln703_491_fu_4467_p2;
reg   [15:0] sub_ln703_491_reg_11793;
wire   [15:0] add_ln703_599_fu_4477_p2;
reg   [15:0] add_ln703_599_reg_11798;
wire   [15:0] add_ln703_609_fu_4501_p2;
reg   [15:0] add_ln703_609_reg_11803;
wire   [15:0] add_ln703_616_fu_4511_p2;
reg   [15:0] add_ln703_616_reg_11808;
wire   [15:0] sub_ln703_503_fu_4516_p2;
reg   [15:0] sub_ln703_503_reg_11813;
wire   [15:0] sub_ln703_505_fu_4521_p2;
reg   [15:0] sub_ln703_505_reg_11818;
wire   [15:0] add_ln703_633_fu_4531_p2;
reg   [15:0] add_ln703_633_reg_11823;
wire   [15:0] add_ln703_634_fu_4535_p2;
reg   [15:0] add_ln703_634_reg_11828;
wire   [15:0] add_ln703_639_fu_4541_p2;
reg   [15:0] add_ln703_639_reg_11833;
wire   [15:0] add_ln703_646_fu_4546_p2;
reg   [15:0] add_ln703_646_reg_11838;
wire   [15:0] add_ln703_650_fu_4550_p2;
reg   [15:0] add_ln703_650_reg_11844;
reg   [15:0] add_ln703_650_reg_11844_pp0_iter11_reg;
wire   [15:0] add_ln703_667_fu_4554_p2;
reg   [15:0] add_ln703_667_reg_11853;
wire   [15:0] sub_ln703_526_fu_4860_p2;
reg   [15:0] sub_ln703_526_reg_11864;
wire   [15:0] sub_ln703_527_fu_4865_p2;
reg   [15:0] sub_ln703_527_reg_11869;
wire   [15:0] add_ln703_647_fu_4870_p2;
reg   [15:0] add_ln703_647_reg_11874;
wire   [15:0] sub_ln703_529_fu_4880_p2;
reg   [15:0] sub_ln703_529_reg_11879;
wire   [15:0] sub_ln703_532_fu_4894_p2;
reg   [15:0] sub_ln703_532_reg_11884;
wire   [15:0] add_ln703_648_fu_4899_p2;
reg   [15:0] add_ln703_648_reg_11889;
wire   [15:0] sub_ln703_533_fu_4904_p2;
reg   [15:0] sub_ln703_533_reg_11894;
wire   [15:0] sub_ln703_535_fu_4919_p2;
reg   [15:0] sub_ln703_535_reg_11899;
wire   [15:0] sub_ln703_538_fu_4934_p2;
reg   [15:0] sub_ln703_538_reg_11904;
wire   [15:0] sub_ln703_539_fu_4939_p2;
reg   [15:0] sub_ln703_539_reg_11909;
wire   [15:0] sub_ln703_540_fu_4944_p2;
reg   [15:0] sub_ln703_540_reg_11914;
wire   [15:0] sub_ln703_541_fu_4949_p2;
reg   [15:0] sub_ln703_541_reg_11919;
wire   [15:0] sub_ln703_542_fu_4954_p2;
reg   [15:0] sub_ln703_542_reg_11924;
wire   [15:0] add_ln703_651_fu_4959_p2;
reg   [15:0] add_ln703_651_reg_11929;
wire   [15:0] sub_ln703_544_fu_4984_p2;
reg   [15:0] sub_ln703_544_reg_11934;
wire   [15:0] add_ln703_660_fu_4994_p2;
reg   [15:0] add_ln703_660_reg_11939;
wire   [15:0] add_ln703_661_fu_4999_p2;
reg   [15:0] add_ln703_661_reg_11944;
wire   [15:0] sub_ln703_551_fu_5004_p2;
reg   [15:0] sub_ln703_551_reg_11949;
wire   [15:0] add_ln703_666_fu_5013_p2;
reg   [15:0] add_ln703_666_reg_11954;
wire   [15:0] add_ln703_668_fu_5019_p2;
reg   [15:0] add_ln703_668_reg_11959;
wire   [15:0] sub_ln703_556_fu_5024_p2;
reg   [15:0] sub_ln703_556_reg_11964;
wire   [15:0] sub_ln703_557_fu_5029_p2;
reg   [15:0] sub_ln703_557_reg_11969;
wire   [15:0] sub_ln703_558_fu_5034_p2;
reg   [15:0] sub_ln703_558_reg_11974;
wire   [15:0] add_ln703_676_fu_5052_p2;
reg   [15:0] add_ln703_676_reg_11979;
wire   [15:0] add_ln703_682_fu_5066_p2;
reg   [15:0] add_ln703_682_reg_11984;
wire   [15:0] add_ln703_685_fu_5077_p2;
reg   [15:0] add_ln703_685_reg_11989;
wire   [15:0] add_ln703_691_fu_5092_p2;
reg   [15:0] add_ln703_691_reg_11994;
wire   [15:0] add_ln703_697_fu_5096_p2;
reg   [15:0] add_ln703_697_reg_12002;
wire   [15:0] sub_ln703_573_fu_5101_p2;
reg   [15:0] sub_ln703_573_reg_12007;
wire   [15:0] sub_ln703_582_fu_5106_p2;
reg   [15:0] sub_ln703_582_reg_12012;
wire   [15:0] sub_ln703_583_fu_5111_p2;
reg   [15:0] sub_ln703_583_reg_12017;
wire   [15:0] add_ln703_703_fu_5116_p2;
reg   [15:0] add_ln703_703_reg_12022;
wire   [15:0] add_ln703_706_fu_5120_p2;
reg   [15:0] add_ln703_706_reg_12031;
wire   [15:0] add_ln703_722_fu_5125_p2;
reg   [15:0] add_ln703_722_reg_12036;
wire   [15:0] add_ln703_726_fu_5130_p2;
reg   [15:0] add_ln703_726_reg_12041;
wire   [15:0] add_ln703_737_fu_5134_p2;
reg   [15:0] add_ln703_737_reg_12047;
wire   [15:0] add_ln703_704_fu_5336_p2;
reg   [15:0] add_ln703_704_reg_12056;
wire   [15:0] sub_ln703_586_fu_5351_p2;
reg   [15:0] sub_ln703_586_reg_12061;
wire   [15:0] sub_ln703_589_fu_5375_p2;
reg   [15:0] sub_ln703_589_reg_12066;
wire   [15:0] sub_ln703_593_fu_5410_p2;
reg   [15:0] sub_ln703_593_reg_12071;
wire   [15:0] sub_ln703_594_fu_5415_p2;
reg   [15:0] sub_ln703_594_reg_12076;
wire   [15:0] sub_ln703_595_fu_5420_p2;
reg   [15:0] sub_ln703_595_reg_12081;
wire   [15:0] add_ln703_719_fu_5439_p2;
reg   [15:0] add_ln703_719_reg_12086;
wire   [15:0] sub_ln703_598_fu_5454_p2;
reg   [15:0] sub_ln703_598_reg_12091;
wire   [15:0] add_ln703_728_fu_5485_p2;
reg   [15:0] add_ln703_728_reg_12096;
wire   [15:0] sub_ln703_603_fu_5491_p2;
reg   [15:0] sub_ln703_603_reg_12101;
wire   [15:0] sub_ln703_604_fu_5496_p2;
reg   [15:0] sub_ln703_604_reg_12106;
wire   [15:0] sub_ln703_605_fu_5501_p2;
reg   [15:0] sub_ln703_605_reg_12111;
wire   [15:0] sub_ln703_608_fu_5511_p2;
reg   [15:0] sub_ln703_608_reg_12116;
wire   [15:0] sub_ln703_609_fu_5516_p2;
reg   [15:0] sub_ln703_609_reg_12121;
wire   [15:0] sub_ln703_610_fu_5521_p2;
reg   [15:0] sub_ln703_610_reg_12126;
wire   [15:0] sub_ln703_612_fu_5526_p2;
reg   [15:0] sub_ln703_612_reg_12131;
wire   [15:0] sub_ln703_613_fu_5531_p2;
reg   [15:0] sub_ln703_613_reg_12136;
wire   [15:0] sub_ln703_614_fu_5536_p2;
reg   [15:0] sub_ln703_614_reg_12141;
wire   [15:0] add_ln703_733_fu_5551_p2;
reg   [15:0] add_ln703_733_reg_12146;
wire   [15:0] add_ln703_734_fu_5556_p2;
reg   [15:0] add_ln703_734_reg_12151;
wire   [15:0] sub_ln703_618_fu_5566_p2;
reg   [15:0] sub_ln703_618_reg_12156;
wire   [15:0] add_ln703_735_fu_5571_p2;
reg   [15:0] add_ln703_735_reg_12161;
wire   [15:0] sub_ln703_624_fu_5596_p2;
reg   [15:0] sub_ln703_624_reg_12166;
wire   [15:0] sub_ln703_630_fu_5627_p2;
reg   [15:0] sub_ln703_630_reg_12171;
wire   [15:0] sub_ln703_631_fu_5632_p2;
reg   [15:0] sub_ln703_631_reg_12176;
wire   [15:0] sub_ln703_634_fu_5637_p2;
reg   [15:0] sub_ln703_634_reg_12181;
wire   [15:0] sub_ln703_637_fu_5642_p2;
reg   [15:0] sub_ln703_637_reg_12186;
wire   [15:0] sub_ln703_638_fu_5647_p2;
reg   [15:0] sub_ln703_638_reg_12191;
wire   [15:0] add_ln703_755_fu_5652_p2;
reg   [15:0] add_ln703_755_reg_12196;
wire   [15:0] sub_ln703_644_fu_5656_p2;
reg   [15:0] sub_ln703_644_reg_12204;
wire   [15:0] sub_ln703_648_fu_5661_p2;
reg   [15:0] sub_ln703_648_reg_12209;
wire   [15:0] sub_ln703_650_fu_5666_p2;
reg   [15:0] sub_ln703_650_reg_12214;
wire   [15:0] add_ln703_765_fu_5671_p2;
reg   [15:0] add_ln703_765_reg_12219;
wire   [15:0] add_ln703_778_fu_5675_p2;
reg   [15:0] add_ln703_778_reg_12227;
wire   [15:0] add_ln703_783_fu_5679_p2;
reg   [15:0] add_ln703_783_reg_12236;
wire   [15:0] add_ln703_816_fu_5684_p2;
reg   [15:0] add_ln703_816_reg_12241;
reg   [15:0] add_ln703_816_reg_12241_pp0_iter13_reg;
wire   [15:0] sub_ln703_662_fu_5918_p2;
reg   [15:0] sub_ln703_662_reg_12248;
wire   [15:0] sub_ln703_665_fu_5932_p2;
reg   [15:0] sub_ln703_665_reg_12253;
wire   [15:0] add_ln703_770_fu_5950_p2;
reg   [15:0] add_ln703_770_reg_12258;
wire   [15:0] sub_ln703_667_fu_5956_p2;
reg   [15:0] sub_ln703_667_reg_12263;
wire   [15:0] sub_ln703_669_fu_5975_p2;
reg   [15:0] sub_ln703_669_reg_12268;
wire   [15:0] add_ln703_779_fu_6024_p2;
reg   [15:0] add_ln703_779_reg_12273;
wire   [15:0] sub_ln703_676_fu_6033_p2;
reg   [15:0] sub_ln703_676_reg_12278;
wire   [15:0] sub_ln703_678_fu_6052_p2;
reg   [15:0] sub_ln703_678_reg_12283;
wire   [15:0] sub_ln703_679_fu_6057_p2;
reg   [15:0] sub_ln703_679_reg_12288;
wire   [15:0] sub_ln703_680_fu_6062_p2;
reg   [15:0] sub_ln703_680_reg_12293;
wire   [15:0] sub_ln703_682_fu_6067_p2;
reg   [15:0] sub_ln703_682_reg_12298;
wire   [15:0] sub_ln703_684_fu_6072_p2;
reg   [15:0] sub_ln703_684_reg_12303;
wire   [15:0] sub_ln703_686_fu_6077_p2;
reg   [15:0] sub_ln703_686_reg_12308;
wire   [15:0] sub_ln703_687_fu_6086_p2;
reg   [15:0] sub_ln703_687_reg_12313;
wire   [15:0] sub_ln703_688_fu_6091_p2;
reg   [15:0] sub_ln703_688_reg_12318;
wire   [15:0] sub_ln703_690_fu_6101_p2;
reg   [15:0] sub_ln703_690_reg_12323;
wire   [15:0] sub_ln703_691_fu_6106_p2;
reg   [15:0] sub_ln703_691_reg_12328;
wire   [15:0] sub_ln703_692_fu_6111_p2;
reg   [15:0] sub_ln703_692_reg_12333;
wire   [15:0] sub_ln703_693_fu_6116_p2;
reg   [15:0] sub_ln703_693_reg_12338;
wire   [15:0] sub_ln703_694_fu_6126_p2;
reg   [15:0] sub_ln703_694_reg_12343;
wire   [15:0] add_ln703_791_fu_6131_p2;
reg   [15:0] add_ln703_791_reg_12348;
wire   [15:0] sub_ln703_696_fu_6136_p2;
reg   [15:0] sub_ln703_696_reg_12353;
wire   [15:0] sub_ln703_697_fu_6141_p2;
reg   [15:0] sub_ln703_697_reg_12358;
wire   [15:0] add_ln703_792_fu_6146_p2;
reg   [15:0] add_ln703_792_reg_12363;
wire   [15:0] add_ln703_796_fu_6160_p2;
reg   [15:0] add_ln703_796_reg_12368;
wire   [15:0] add_ln703_798_fu_6166_p2;
reg   [15:0] add_ln703_798_reg_12373;
wire   [15:0] sub_ln703_700_fu_6172_p2;
reg   [15:0] sub_ln703_700_reg_12378;
wire   [15:0] sub_ln703_704_fu_6177_p2;
reg   [15:0] sub_ln703_704_reg_12383;
wire   [15:0] sub_ln703_707_fu_6182_p2;
reg   [15:0] sub_ln703_707_reg_12388;
wire   [15:0] add_ln703_801_fu_6187_p2;
reg   [15:0] add_ln703_801_reg_12393;
wire   [15:0] add_ln703_802_fu_6192_p2;
reg   [15:0] add_ln703_802_reg_12398;
wire   [15:0] add_ln703_818_fu_6205_p2;
reg   [15:0] add_ln703_818_reg_12409;
reg   [15:0] add_ln703_818_reg_12409_pp0_iter14_reg;
wire   [15:0] add_ln703_821_fu_6216_p2;
reg   [15:0] add_ln703_821_reg_12414;
wire   [15:0] add_ln703_826_fu_6222_p2;
reg   [15:0] add_ln703_826_reg_12419;
wire   [15:0] add_ln703_836_fu_6226_p2;
reg   [15:0] add_ln703_836_reg_12428;
wire   [15:0] add_ln703_849_fu_6230_p2;
reg   [15:0] add_ln703_849_reg_12434;
reg   [15:0] add_ln703_849_reg_12434_pp0_iter14_reg;
wire   [15:0] add_ln703_867_fu_6234_p2;
reg   [15:0] add_ln703_867_reg_12444;
reg   [15:0] add_ln703_867_reg_12444_pp0_iter14_reg;
wire   [15:0] sub_ln703_724_fu_6432_p2;
reg   [15:0] sub_ln703_724_reg_12450;
wire   [15:0] add_ln703_819_fu_6447_p2;
reg   [15:0] add_ln703_819_reg_12455;
wire   [15:0] sub_ln703_727_fu_6452_p2;
reg   [15:0] sub_ln703_727_reg_12460;
wire   [15:0] sub_ln703_728_fu_6457_p2;
reg   [15:0] sub_ln703_728_reg_12465;
wire   [15:0] sub_ln703_733_fu_6487_p2;
reg   [15:0] sub_ln703_733_reg_12470;
wire   [15:0] sub_ln703_736_fu_6502_p2;
reg   [15:0] sub_ln703_736_reg_12475;
wire   [15:0] add_ln703_825_fu_6526_p2;
reg   [15:0] add_ln703_825_reg_12480;
wire   [15:0] add_ln703_827_fu_6531_p2;
reg   [15:0] add_ln703_827_reg_12485;
wire   [15:0] add_ln703_831_fu_6554_p2;
reg   [15:0] add_ln703_831_reg_12490;
wire   [15:0] add_ln703_833_fu_6573_p2;
reg   [15:0] add_ln703_833_reg_12495;
wire   [15:0] sub_ln703_746_fu_6579_p2;
reg   [15:0] sub_ln703_746_reg_12500;
wire   [15:0] add_ln703_834_fu_6594_p2;
reg   [15:0] add_ln703_834_reg_12505;
wire   [15:0] sub_ln703_749_fu_6599_p2;
reg   [15:0] sub_ln703_749_reg_12510;
wire   [15:0] sub_ln703_757_fu_6629_p2;
reg   [15:0] sub_ln703_757_reg_12515;
wire   [15:0] add_ln703_838_fu_6634_p2;
reg   [15:0] add_ln703_838_reg_12520;
wire   [15:0] sub_ln703_759_fu_6639_p2;
reg   [15:0] sub_ln703_759_reg_12525;
wire   [15:0] sub_ln703_761_fu_6644_p2;
reg   [15:0] sub_ln703_761_reg_12530;
wire   [15:0] add_ln703_840_fu_6649_p2;
reg   [15:0] add_ln703_840_reg_12535;
wire   [15:0] sub_ln703_763_fu_6654_p2;
reg   [15:0] sub_ln703_763_reg_12540;
wire   [15:0] sub_ln703_767_fu_6659_p2;
reg   [15:0] sub_ln703_767_reg_12545;
wire   [15:0] add_ln703_841_fu_6664_p2;
reg   [15:0] add_ln703_841_reg_12550;
wire   [15:0] sub_ln703_769_fu_6684_p2;
reg   [15:0] sub_ln703_769_reg_12555;
wire   [15:0] add_ln703_845_fu_6689_p2;
reg   [15:0] add_ln703_845_reg_12560;
wire   [15:0] add_ln703_851_fu_6702_p2;
reg   [15:0] add_ln703_851_reg_12565;
wire   [15:0] sub_ln703_770_fu_6708_p2;
reg   [15:0] sub_ln703_770_reg_12570;
wire   [15:0] add_ln703_858_fu_6733_p2;
reg   [15:0] add_ln703_858_reg_12575;
wire   [15:0] sub_ln703_781_fu_6739_p2;
reg   [15:0] sub_ln703_781_reg_12580;
wire   [15:0] add_ln703_868_fu_6755_p2;
reg   [15:0] add_ln703_868_reg_12585;
wire   [15:0] sub_ln703_787_fu_6759_p2;
reg   [15:0] sub_ln703_787_reg_12590;
wire   [15:0] sub_ln703_799_fu_6764_p2;
reg   [15:0] sub_ln703_799_reg_12595;
wire   [15:0] add_ln703_876_fu_6769_p2;
reg   [15:0] add_ln703_876_reg_12600;
wire   [15:0] add_ln703_877_fu_6774_p2;
reg   [15:0] add_ln703_877_reg_12605;
wire   [15:0] add_ln703_894_fu_6778_p2;
reg   [15:0] add_ln703_894_reg_12616;
reg   [15:0] add_ln703_894_reg_12616_pp0_iter15_reg;
wire   [15:0] add_ln703_905_fu_6782_p2;
reg   [15:0] add_ln703_905_reg_12625;
wire   [15:0] add_ln703_914_fu_6786_p2;
reg   [15:0] add_ln703_914_reg_12632;
wire   [15:0] add_ln703_920_fu_6791_p2;
reg   [15:0] add_ln703_920_reg_12637;
reg   [15:0] add_ln703_920_reg_12637_pp0_iter15_reg;
wire   [15:0] sub_ln703_797_fu_7030_p2;
reg   [15:0] sub_ln703_797_reg_12645;
wire   [15:0] add_ln703_872_fu_7050_p2;
reg   [15:0] add_ln703_872_reg_12650;
wire   [15:0] add_ln703_873_fu_7055_p2;
reg   [15:0] add_ln703_873_reg_12655;
wire   [15:0] sub_ln703_801_fu_7060_p2;
reg   [15:0] sub_ln703_801_reg_12660;
wire   [15:0] sub_ln703_802_fu_7065_p2;
reg   [15:0] sub_ln703_802_reg_12665;
wire   [15:0] sub_ln703_805_fu_7079_p2;
reg   [15:0] sub_ln703_805_reg_12670;
wire   [15:0] add_ln703_874_fu_7084_p2;
reg   [15:0] add_ln703_874_reg_12675;
wire   [15:0] add_ln703_875_fu_7094_p2;
reg   [15:0] add_ln703_875_reg_12680;
wire   [15:0] sub_ln703_807_fu_7099_p2;
reg   [15:0] sub_ln703_807_reg_12685;
wire   [15:0] add_ln703_882_fu_7121_p2;
reg   [15:0] add_ln703_882_reg_12690;
wire   [15:0] add_ln703_884_fu_7132_p2;
reg   [15:0] add_ln703_884_reg_12695;
wire   [15:0] sub_ln703_808_fu_7137_p2;
reg   [15:0] sub_ln703_808_reg_12700;
wire   [15:0] add_ln703_888_fu_7156_p2;
reg   [15:0] add_ln703_888_reg_12705;
wire   [15:0] add_ln703_892_fu_7175_p2;
reg   [15:0] add_ln703_892_reg_12710;
wire   [15:0] add_ln703_893_fu_7180_p2;
reg   [15:0] add_ln703_893_reg_12715;
wire   [15:0] add_ln703_895_fu_7185_p2;
reg   [15:0] add_ln703_895_reg_12720;
wire   [15:0] add_ln703_896_fu_7190_p2;
reg   [15:0] add_ln703_896_reg_12725;
wire   [15:0] add_ln703_898_fu_7195_p2;
reg   [15:0] add_ln703_898_reg_12730;
wire   [15:0] sub_ln703_814_fu_7200_p2;
reg   [15:0] sub_ln703_814_reg_12735;
wire   [15:0] sub_ln703_816_fu_7205_p2;
reg   [15:0] sub_ln703_816_reg_12740;
wire   [15:0] sub_ln703_818_fu_7210_p2;
reg   [15:0] sub_ln703_818_reg_12745;
wire   [15:0] sub_ln703_820_fu_7215_p2;
reg   [15:0] sub_ln703_820_reg_12750;
wire   [15:0] sub_ln703_821_fu_7220_p2;
reg   [15:0] sub_ln703_821_reg_12755;
wire   [15:0] sub_ln703_823_fu_7225_p2;
reg   [15:0] sub_ln703_823_reg_12760;
wire   [15:0] sub_ln703_824_fu_7230_p2;
reg   [15:0] sub_ln703_824_reg_12765;
wire   [15:0] sub_ln703_825_fu_7235_p2;
reg   [15:0] sub_ln703_825_reg_12770;
wire   [15:0] add_ln703_906_fu_7245_p2;
reg   [15:0] add_ln703_906_reg_12775;
wire   [15:0] add_ln703_917_fu_7273_p2;
reg   [15:0] add_ln703_917_reg_12780;
wire   [15:0] add_ln703_922_fu_7287_p2;
reg   [15:0] add_ln703_922_reg_12785;
wire   [15:0] sub_ln703_852_fu_7319_p2;
reg   [15:0] sub_ln703_852_reg_12790;
wire   [15:0] sub_ln703_862_fu_7324_p2;
reg   [15:0] sub_ln703_862_reg_12795;
wire   [15:0] sub_ln703_869_fu_7329_p2;
reg   [15:0] sub_ln703_869_reg_12800;
reg   [15:0] sub_ln703_869_reg_12800_pp0_iter16_reg;
wire   [15:0] add_ln703_946_fu_7334_p2;
reg   [15:0] add_ln703_946_reg_12805;
wire   [15:0] add_ln703_954_fu_7338_p2;
reg   [15:0] add_ln703_954_reg_12812;
wire   [15:0] add_ln703_985_fu_7342_p2;
reg   [15:0] add_ln703_985_reg_12819;
reg   [15:0] add_ln703_985_reg_12819_pp0_iter16_reg;
wire   [15:0] sub_ln703_857_fu_7600_p2;
reg   [15:0] sub_ln703_857_reg_12835;
wire   [15:0] sub_ln703_858_fu_7605_p2;
reg   [15:0] sub_ln703_858_reg_12840;
wire   [15:0] add_ln703_934_fu_7610_p2;
reg   [15:0] add_ln703_934_reg_12845;
wire   [15:0] sub_ln703_859_fu_7615_p2;
reg   [15:0] sub_ln703_859_reg_12850;
wire   [15:0] add_ln703_936_fu_7634_p2;
reg   [15:0] add_ln703_936_reg_12855;
wire   [15:0] sub_ln703_863_fu_7639_p2;
reg   [15:0] sub_ln703_863_reg_12860;
wire   [15:0] sub_ln703_865_fu_7649_p2;
reg   [15:0] sub_ln703_865_reg_12865;
wire   [15:0] sub_ln703_866_fu_7654_p2;
reg   [15:0] sub_ln703_866_reg_12870;
wire   [15:0] add_ln703_938_fu_7663_p2;
reg   [15:0] add_ln703_938_reg_12875;
wire   [15:0] sub_ln703_867_fu_7669_p2;
reg   [15:0] sub_ln703_867_reg_12880;
wire   [15:0] sub_ln703_868_fu_7674_p2;
reg   [15:0] sub_ln703_868_reg_12885;
wire   [15:0] add_ln703_939_fu_7679_p2;
reg   [15:0] add_ln703_939_reg_12890;
wire   [15:0] sub_ln703_870_fu_7685_p2;
reg   [15:0] sub_ln703_870_reg_12895;
wire   [15:0] sub_ln703_873_fu_7710_p2;
reg   [15:0] sub_ln703_873_reg_12900;
wire   [15:0] add_ln703_943_fu_7719_p2;
reg   [15:0] add_ln703_943_reg_12905;
wire   [15:0] sub_ln703_875_fu_7730_p2;
reg   [15:0] sub_ln703_875_reg_12910;
wire   [15:0] sub_ln703_879_fu_7735_p2;
reg   [15:0] sub_ln703_879_reg_12915;
wire   [15:0] sub_ln703_880_fu_7750_p2;
reg   [15:0] sub_ln703_880_reg_12920;
wire   [15:0] sub_ln703_881_fu_7755_p2;
reg   [15:0] sub_ln703_881_reg_12925;
wire   [15:0] add_ln703_948_fu_7760_p2;
reg   [15:0] add_ln703_948_reg_12930;
wire   [15:0] sub_ln703_892_fu_7780_p2;
reg   [15:0] sub_ln703_892_reg_12935;
wire   [15:0] sub_ln703_893_fu_7785_p2;
reg   [15:0] sub_ln703_893_reg_12940;
wire   [15:0] sub_ln703_894_fu_7790_p2;
reg   [15:0] sub_ln703_894_reg_12945;
wire   [15:0] sub_ln703_895_fu_7795_p2;
reg   [15:0] sub_ln703_895_reg_12950;
wire   [15:0] sub_ln703_898_fu_7805_p2;
reg   [15:0] sub_ln703_898_reg_12955;
wire   [15:0] sub_ln703_904_fu_7810_p2;
reg   [15:0] sub_ln703_904_reg_12960;
wire   [15:0] add_ln703_958_fu_7827_p2;
reg   [15:0] add_ln703_958_reg_12965;
wire   [15:0] sub_ln703_911_fu_7833_p2;
reg   [15:0] sub_ln703_911_reg_12970;
wire   [15:0] sub_ln703_917_fu_7838_p2;
reg   [15:0] sub_ln703_917_reg_12975;
wire   [15:0] sub_ln703_922_fu_7843_p2;
reg   [15:0] sub_ln703_922_reg_12980;
wire   [15:0] add_ln703_964_fu_7848_p2;
reg   [15:0] add_ln703_964_reg_12985;
wire   [15:0] acc_21_V_fu_7872_p2;
reg   [15:0] acc_21_V_reg_12991;
wire    ap_block_pp0_stage0;
wire   [15:0] sub_ln703_5_fu_564_p2;
wire   [15:0] add_ln703_143_fu_585_p2;
wire   [15:0] add_ln703_142_fu_581_p2;
wire   [15:0] add_ln703_133_fu_603_p2;
wire   [15:0] sub_ln703_7_fu_607_p2;
wire   [15:0] sub_ln703_9_fu_611_p2;
wire   [15:0] add_ln703_136_fu_623_p2;
wire   [15:0] add_ln703_139_fu_636_p2;
wire   [15:0] sub_ln703_12_fu_627_p2;
wire   [15:0] sub_ln703_13_fu_689_p2;
wire   [15:0] sub_ln703_14_fu_693_p2;
wire   [15:0] add_ln703_137_fu_697_p2;
wire   [15:0] add_ln703_138_fu_701_p2;
wire   [15:0] sub_ln703_19_fu_705_p2;
wire   [15:0] sub_ln703_22_fu_713_p2;
wire   [15:0] sub_ln703_24_fu_717_p2;
wire   [15:0] sub_ln703_25_fu_722_p2;
wire   [15:0] sub_ln703_27_fu_732_p2;
wire   [15:0] add_ln703_145_fu_736_p2;
wire   [15:0] add_ln703_146_fu_741_p2;
wire   [15:0] add_ln703_147_fu_745_p2;
wire   [15:0] sub_ln703_29_fu_749_p2;
wire   [15:0] sub_ln703_30_fu_753_p2;
wire   [15:0] add_ln703_148_fu_757_p2;
wire   [15:0] sub_ln703_31_fu_761_p2;
wire   [15:0] sub_ln703_32_fu_765_p2;
wire   [15:0] sub_ln703_33_fu_769_p2;
wire   [15:0] add_ln703_155_fu_868_p2;
wire   [15:0] add_ln703_149_fu_773_p2;
wire   [15:0] sub_ln703_34_fu_778_p2;
wire   [15:0] add_ln703_150_fu_782_p2;
wire   [15:0] sub_ln703_35_fu_787_p2;
wire   [15:0] add_ln703_151_fu_791_p2;
wire   [15:0] sub_ln703_37_fu_800_p2;
wire   [15:0] add_ln703_152_fu_804_p2;
wire   [15:0] sub_ln703_26_fu_727_p2;
wire   [15:0] sub_ln703_41_fu_829_p2;
wire   [15:0] add_ln703_154_fu_843_p2;
wire   [15:0] sub_ln703_44_fu_848_p2;
wire   [15:0] sub_ln703_45_fu_853_p2;
wire   [15:0] add_ln703_156_fu_872_p2;
wire   [15:0] sub_ln703_48_fu_877_p2;
wire   [15:0] sub_ln703_49_fu_882_p2;
wire   [15:0] sub_ln703_21_fu_709_p2;
wire   [15:0] add_ln703_166_fu_962_p2;
wire   [15:0] sub_ln703_51_fu_897_p2;
wire   [15:0] sub_ln703_36_fu_795_p2;
wire   [15:0] add_ln703_160_fu_902_p2;
wire   [15:0] sub_ln703_60_fu_927_p2;
wire   [15:0] sub_ln703_61_fu_932_p2;
wire   [15:0] add_ln703_164_fu_937_p2;
wire   [15:0] add_ln703_180_fu_1011_p2;
wire   [15:0] add_ln703_178_fu_1007_p2;
wire   [15:0] sub_ln703_47_fu_863_p2;
wire   [15:0] add_ln703_165_fu_952_p2;
wire   [15:0] add_ln703_168_fu_967_p2;
wire   [15:0] sub_ln703_50_fu_887_p2;
wire   [15:0] add_ln703_187_fu_1041_p2;
wire   [15:0] add_ln703_189_fu_1045_p2;
wire   [15:0] sub_ln703_52_fu_907_p2;
wire   [15:0] sub_ln703_46_fu_858_p2;
wire   [15:0] sub_ln703_42_fu_833_p2;
wire   [15:0] sub_ln703_54_fu_1086_p2;
wire   [15:0] sub_ln703_55_fu_1090_p2;
wire   [15:0] sub_ln703_56_fu_1094_p2;
wire   [15:0] add_ln703_163_fu_1098_p2;
wire   [15:0] sub_ln703_57_fu_1102_p2;
wire   [15:0] sub_ln703_65_fu_1110_p2;
wire   [15:0] add_ln703_174_fu_1114_p2;
wire   [15:0] sub_ln703_67_fu_1119_p2;
wire   [15:0] add_ln703_175_fu_1123_p2;
wire   [15:0] add_ln703_176_fu_1128_p2;
wire   [15:0] sub_ln703_69_fu_1138_p2;
wire   [15:0] sub_ln703_59_fu_1106_p2;
wire   [15:0] add_ln703_184_fu_1143_p2;
wire   [15:0] sub_ln703_72_fu_1147_p2;
wire   [15:0] sub_ln703_74_fu_1151_p2;
wire   [15:0] sub_ln703_77_fu_1159_p2;
wire   [15:0] sub_ln703_78_fu_1164_p2;
wire   [15:0] sub_ln703_79_fu_1168_p2;
wire   [15:0] add_ln703_190_fu_1172_p2;
wire   [15:0] add_ln703_191_fu_1176_p2;
wire   [15:0] add_ln703_193_fu_1180_p2;
wire   [15:0] sub_ln703_80_fu_1184_p2;
wire   [15:0] add_ln703_194_fu_1189_p2;
wire   [15:0] sub_ln703_82_fu_1199_p2;
wire   [15:0] sub_ln703_68_fu_1133_p2;
wire   [15:0] add_ln703_195_fu_1204_p2;
wire   [15:0] add_ln703_197_fu_1209_p2;
wire   [15:0] add_ln703_199_fu_1213_p2;
wire   [15:0] sub_ln703_83_fu_1218_p2;
wire   [15:0] sub_ln703_84_fu_1222_p2;
wire   [15:0] add_ln703_200_fu_1226_p2;
wire   [15:0] add_ln703_214_fu_1349_p2;
wire   [15:0] sub_ln703_85_fu_1230_p2;
wire   [15:0] sub_ln703_87_fu_1238_p2;
wire   [15:0] add_ln703_201_fu_1243_p2;
wire   [15:0] sub_ln703_88_fu_1248_p2;
wire   [15:0] sub_ln703_89_fu_1252_p2;
wire   [15:0] sub_ln703_90_fu_1257_p2;
wire   [15:0] sub_ln703_91_fu_1261_p2;
wire   [15:0] add_ln703_217_fu_1393_p2;
wire   [15:0] sub_ln703_76_fu_1155_p2;
wire   [15:0] add_ln703_202_fu_1265_p2;
wire   [15:0] add_ln703_203_fu_1270_p2;
wire   [15:0] sub_ln703_93_fu_1275_p2;
wire   [15:0] sub_ln703_94_fu_1280_p2;
wire   [15:0] add_ln703_206_fu_1290_p2;
wire   [15:0] sub_ln703_97_fu_1304_p2;
wire   [15:0] sub_ln703_81_fu_1194_p2;
wire   [15:0] sub_ln703_99_fu_1324_p2;
wire   [15:0] add_ln703_211_fu_1339_p2;
wire   [15:0] sub_ln703_102_fu_1344_p2;
wire   [15:0] add_ln703_215_fu_1353_p2;
wire   [15:0] sub_ln703_103_fu_1363_p2;
wire   [15:0] sub_ln703_104_fu_1368_p2;
wire   [15:0] sub_ln703_105_fu_1373_p2;
wire   [15:0] add_ln703_219_fu_1397_p2;
wire   [15:0] add_ln703_221_fu_1402_p2;
wire   [15:0] sub_ln703_111_fu_1417_p2;
wire   [15:0] sub_ln703_112_fu_1422_p2;
wire   [15:0] sub_ln703_113_fu_1427_p2;
wire   [15:0] sub_ln703_119_fu_1442_p2;
wire   [15:0] add_ln703_237_fu_1516_p2;
wire   [15:0] sub_ln703_100_fu_1329_p2;
wire   [15:0] sub_ln703_101_fu_1334_p2;
wire   [15:0] add_ln703_225_fu_1452_p2;
wire   [15:0] sub_ln703_86_fu_1234_p2;
wire   [15:0] add_ln703_242_fu_1537_p2;
wire   [15:0] add_ln703_228_fu_1477_p2;
wire   [15:0] sub_ln703_126_fu_1487_p2;
wire   [15:0] add_ln703_232_fu_1492_p2;
wire   [15:0] sub_ln703_110_fu_1412_p2;
wire   [15:0] sub_ln703_95_fu_1285_p2;
wire   [15:0] add_ln703_248_fu_1569_p2;
wire   [15:0] sub_ln703_129_fu_1506_p2;
wire   [15:0] add_ln703_259_fu_1589_p2;
wire   [15:0] add_ln703_256_fu_1585_p2;
wire   [15:0] add_ln703_240_fu_1526_p2;
wire   [15:0] sub_ln703_120_fu_1447_p2;
wire   [15:0] add_ln703_244_fu_1542_p2;
wire   [15:0] add_ln703_222_fu_1626_p2;
wire   [15:0] sub_ln703_114_fu_1630_p2;
wire   [15:0] sub_ln703_118_fu_1642_p2;
wire   [15:0] sub_ln703_121_fu_1646_p2;
wire   [15:0] sub_ln703_124_fu_1650_p2;
wire   [15:0] add_ln703_229_fu_1654_p2;
wire   [15:0] add_ln703_230_fu_1658_p2;
wire   [15:0] sub_ln703_127_fu_1662_p2;
wire   [15:0] sub_ln703_130_fu_1666_p2;
wire   [15:0] add_ln703_234_fu_1671_p2;
wire   [15:0] add_ln703_235_fu_1676_p2;
wire   [15:0] sub_ln703_131_fu_1680_p2;
wire   [15:0] sub_ln703_117_fu_1638_p2;
wire   [15:0] add_ln703_241_fu_1693_p2;
wire   [15:0] sub_ln703_135_fu_1698_p2;
wire   [15:0] sub_ln703_136_fu_1702_p2;
wire   [15:0] sub_ln703_139_fu_1711_p2;
wire   [15:0] sub_ln703_140_fu_1716_p2;
wire   [15:0] add_ln703_245_fu_1721_p2;
wire   [15:0] sub_ln703_145_fu_1734_p2;
wire   [15:0] sub_ln703_148_fu_1743_p2;
wire   [15:0] sub_ln703_149_fu_1748_p2;
wire   [15:0] add_ln703_251_fu_1753_p2;
wire   [15:0] add_ln703_253_fu_1758_p2;
wire   [15:0] sub_ln703_132_fu_1684_p2;
wire   [15:0] sub_ln703_150_fu_1763_p2;
wire   [15:0] sub_ln703_151_fu_1767_p2;
wire   [15:0] add_ln703_263_fu_1771_p2;
wire   [15:0] sub_ln703_134_fu_1689_p2;
wire   [15:0] add_ln703_269_fu_1891_p2;
wire   [15:0] sub_ln703_156_fu_1785_p2;
wire   [15:0] sub_ln703_157_fu_1790_p2;
wire   [15:0] sub_ln703_138_fu_1706_p2;
wire   [15:0] sub_ln703_160_fu_1804_p2;
wire   [15:0] sub_ln703_161_fu_1809_p2;
wire   [15:0] sub_ln703_162_fu_1813_p2;
wire   [15:0] sub_ln703_143_fu_1725_p2;
wire   [15:0] sub_ln703_163_fu_1817_p2;
wire   [15:0] add_ln703_264_fu_1821_p2;
wire   [15:0] sub_ln703_164_fu_1826_p2;
wire   [15:0] sub_ln703_165_fu_1830_p2;
wire   [15:0] sub_ln703_168_fu_1844_p2;
wire   [15:0] sub_ln703_116_fu_1634_p2;
wire   [15:0] add_ln703_281_fu_1969_p2;
wire   [15:0] add_ln703_279_fu_1964_p2;
wire   [15:0] sub_ln703_169_fu_1849_p2;
wire   [15:0] add_ln703_266_fu_1854_p2;
wire   [15:0] sub_ln703_172_fu_1868_p2;
wire   [15:0] sub_ln703_173_fu_1873_p2;
wire   [15:0] sub_ln703_174_fu_1877_p2;
wire   [15:0] add_ln703_268_fu_1886_p2;
wire   [15:0] sub_ln703_153_fu_1775_p2;
wire   [15:0] add_ln703_271_fu_1895_p2;
wire   [15:0] sub_ln703_155_fu_1780_p2;
wire   [15:0] sub_ln703_178_fu_1909_p2;
wire   [15:0] add_ln703_273_fu_1914_p2;
wire   [15:0] sub_ln703_158_fu_1794_p2;
wire   [15:0] sub_ln703_179_fu_1919_p2;
wire   [15:0] add_ln703_274_fu_1924_p2;
wire   [15:0] sub_ln703_180_fu_1929_p2;
wire   [15:0] add_ln703_276_fu_1934_p2;
wire   [15:0] add_ln703_277_fu_1939_p2;
wire   [15:0] sub_ln703_144_fu_1730_p2;
wire   [15:0] add_ln703_291_fu_2064_p2;
wire   [15:0] sub_ln703_181_fu_1944_p2;
wire   [15:0] add_ln703_278_fu_1954_p2;
wire   [15:0] sub_ln703_147_fu_1738_p2;
wire   [15:0] sub_ln703_167_fu_1839_p2;
wire   [15:0] add_ln703_282_fu_1973_p2;
wire   [15:0] sub_ln703_171_fu_1864_p2;
wire   [15:0] sub_ln703_185_fu_1989_p2;
wire   [15:0] sub_ln703_188_fu_2004_p2;
wire   [15:0] sub_ln703_189_fu_2014_p2;
wire   [15:0] sub_ln703_176_fu_1900_p2;
wire   [15:0] add_ln703_287_fu_2019_p2;
wire   [15:0] sub_ln703_177_fu_1904_p2;
wire   [15:0] sub_ln703_190_fu_2024_p2;
wire   [15:0] sub_ln703_159_fu_1799_p2;
wire   [15:0] sub_ln703_192_fu_2044_p2;
wire   [15:0] sub_ln703_195_fu_2059_p2;
wire   [15:0] add_ln703_293_fu_2069_p2;
wire   [15:0] sub_ln703_182_fu_1949_p2;
wire   [15:0] sub_ln703_197_fu_2079_p2;
wire   [15:0] add_ln703_316_fu_2178_p2;
wire   [15:0] sub_ln703_187_fu_1999_p2;
wire   [15:0] sub_ln703_193_fu_2049_p2;
wire   [15:0] add_ln703_314_fu_2167_p2;
wire   [15:0] sub_ln703_170_fu_1859_p2;
wire   [15:0] add_ln703_327_fu_2204_p2;
wire   [15:0] add_ln703_325_fu_2199_p2;
wire   [15:0] add_ln703_317_fu_2182_p2;
wire   [15:0] sub_ln703_175_fu_1881_p2;
wire   [15:0] add_ln703_330_fu_2219_p2;
wire   [15:0] add_ln703_296_fu_2238_p2;
wire   [15:0] add_ln703_298_fu_2242_p2;
wire   [15:0] sub_ln703_199_fu_2246_p2;
wire   [15:0] add_ln703_301_fu_2250_p2;
wire   [15:0] add_ln703_305_fu_2254_p2;
wire   [15:0] sub_ln703_201_fu_2258_p2;
wire   [15:0] sub_ln703_205_fu_2262_p2;
wire   [15:0] sub_ln703_206_fu_2266_p2;
wire   [15:0] add_ln703_312_fu_2270_p2;
wire   [15:0] sub_ln703_207_fu_2274_p2;
wire   [15:0] sub_ln703_211_fu_2278_p2;
wire   [15:0] sub_ln703_213_fu_2282_p2;
wire   [15:0] sub_ln703_215_fu_2292_p2;
wire   [15:0] sub_ln703_216_fu_2296_p2;
wire   [15:0] add_ln703_315_fu_2300_p2;
wire   [15:0] sub_ln703_217_fu_2305_p2;
wire   [15:0] sub_ln703_218_fu_2310_p2;
wire   [15:0] sub_ln703_220_fu_2318_p2;
wire   [15:0] add_ln703_318_fu_2323_p2;
wire   [15:0] add_ln703_319_fu_2328_p2;
wire   [15:0] sub_ln703_221_fu_2332_p2;
wire   [15:0] add_ln703_320_fu_2336_p2;
wire   [15:0] sub_ln703_222_fu_2340_p2;
wire   [15:0] sub_ln703_224_fu_2348_p2;
wire   [15:0] add_ln703_321_fu_2353_p2;
wire   [15:0] sub_ln703_225_fu_2358_p2;
wire   [15:0] sub_ln703_227_fu_2368_p2;
wire   [15:0] sub_ln703_228_fu_2372_p2;
wire   [15:0] sub_ln703_229_fu_2376_p2;
wire   [15:0] sub_ln703_231_fu_2381_p2;
wire   [15:0] sub_ln703_232_fu_2385_p2;
wire   [15:0] sub_ln703_235_fu_2400_p2;
wire   [15:0] add_ln703_324_fu_2405_p2;
wire   [15:0] add_ln703_329_fu_2410_p2;
wire   [15:0] sub_ln703_219_fu_2314_p2;
wire   [15:0] sub_ln703_236_fu_2415_p2;
wire   [15:0] add_ln703_335_fu_2420_p2;
wire   [15:0] sub_ln703_238_fu_2424_p2;
wire   [15:0] sub_ln703_239_fu_2429_p2;
wire   [15:0] sub_ln703_240_fu_2434_p2;
wire   [15:0] sub_ln703_241_fu_2439_p2;
wire   [15:0] sub_ln703_242_fu_2444_p2;
wire   [15:0] sub_ln703_223_fu_2344_p2;
wire   [15:0] add_ln703_336_fu_2449_p2;
wire   [15:0] sub_ln703_243_fu_2454_p2;
wire   [15:0] add_ln703_337_fu_2459_p2;
wire   [15:0] add_ln703_339_fu_2464_p2;
wire   [15:0] sub_ln703_244_fu_2468_p2;
wire   [15:0] add_ln703_349_fu_2598_p2;
wire   [15:0] add_ln703_347_fu_2594_p2;
wire   [15:0] sub_ln703_245_fu_2472_p2;
wire   [15:0] sub_ln703_247_fu_2482_p2;
wire   [15:0] sub_ln703_248_fu_2487_p2;
wire   [15:0] add_ln703_340_fu_2491_p2;
wire   [15:0] sub_ln703_252_fu_2511_p2;
wire   [15:0] sub_ln703_253_fu_2515_p2;
wire   [15:0] sub_ln703_255_fu_2530_p2;
wire   [15:0] sub_ln703_258_fu_2544_p2;
wire   [15:0] sub_ln703_259_fu_2549_p2;
wire   [15:0] add_ln703_343_fu_2554_p2;
wire   [15:0] add_ln703_345_fu_2564_p2;
wire   [15:0] sub_ln703_226_fu_2363_p2;
wire   [15:0] add_ln703_358_fu_2672_p2;
wire   [15:0] sub_ln703_264_fu_2584_p2;
wire   [15:0] add_ln703_351_fu_2608_p2;
wire   [15:0] sub_ln703_266_fu_2618_p2;
wire   [15:0] sub_ln703_267_fu_2623_p2;
wire   [15:0] add_ln703_355_fu_2642_p2;
wire   [15:0] sub_ln703_276_fu_2667_p2;
wire   [15:0] add_ln703_361_fu_2683_p2;
wire   [15:0] sub_ln703_283_fu_2693_p2;
wire   [15:0] sub_ln703_233_fu_2390_p2;
wire   [15:0] add_ln703_370_fu_2728_p2;
wire   [15:0] add_ln703_368_fu_2723_p2;
wire   [15:0] sub_ln703_260_fu_2559_p2;
wire   [15:0] sub_ln703_214_fu_2287_p2;
wire   [15:0] add_ln703_398_fu_2747_p2;
wire   [15:0] add_ln703_523_fu_2770_p2;
wire   [15:0] sub_ln703_268_fu_2783_p2;
wire   [15:0] sub_ln703_269_fu_2787_p2;
wire   [15:0] sub_ln703_271_fu_2791_p2;
wire   [15:0] add_ln703_353_fu_2795_p2;
wire   [15:0] add_ln703_357_fu_2811_p2;
wire   [15:0] sub_ln703_279_fu_2815_p2;
wire   [15:0] sub_ln703_280_fu_2819_p2;
wire   [15:0] add_ln703_363_fu_2823_p2;
wire   [15:0] add_ln703_364_fu_2831_p2;
wire   [15:0] sub_ln703_285_fu_2836_p2;
wire   [15:0] add_ln703_365_fu_2841_p2;
wire   [15:0] sub_ln703_286_fu_2845_p2;
wire   [15:0] sub_ln703_290_fu_2859_p2;
wire   [15:0] sub_ln703_273_fu_2799_p2;
wire   [15:0] sub_ln703_291_fu_2863_p2;
wire   [15:0] sub_ln703_292_fu_2867_p2;
wire   [15:0] add_ln703_366_fu_2871_p2;
wire   [15:0] sub_ln703_295_fu_2880_p2;
wire   [15:0] sub_ln703_297_fu_2884_p2;
wire   [15:0] sub_ln703_298_fu_2889_p2;
wire   [15:0] sub_ln703_299_fu_2894_p2;
wire   [15:0] sub_ln703_300_fu_2898_p2;
wire   [15:0] add_ln703_367_fu_2903_p2;
wire   [15:0] sub_ln703_302_fu_2907_p2;
wire   [15:0] add_ln703_385_fu_3011_p2;
wire   [15:0] add_ln703_383_fu_3007_p2;
wire   [15:0] sub_ln703_303_fu_2912_p2;
wire   [15:0] sub_ln703_304_fu_2917_p2;
wire   [15:0] add_ln703_372_fu_2927_p2;
wire   [15:0] sub_ln703_306_fu_2931_p2;
wire   [15:0] add_ln703_374_fu_2936_p2;
wire   [15:0] add_ln703_387_fu_3046_p2;
wire   [15:0] sub_ln703_307_fu_2941_p2;
wire   [15:0] sub_ln703_308_fu_2946_p2;
wire   [15:0] sub_ln703_309_fu_2951_p2;
wire   [15:0] add_ln703_377_fu_2956_p2;
wire   [15:0] add_ln703_378_fu_2960_p2;
wire   [15:0] sub_ln703_277_fu_2803_p2;
wire   [15:0] add_ln703_392_fu_3081_p2;
wire   [15:0] add_ln703_379_fu_2964_p2;
wire   [15:0] add_ln703_380_fu_2969_p2;
wire   [15:0] add_ln703_381_fu_2973_p2;
wire   [15:0] add_ln703_382_fu_2983_p2;
wire   [15:0] sub_ln703_311_fu_2988_p2;
wire   [15:0] sub_ln703_282_fu_2827_p2;
wire   [15:0] add_ln703_395_fu_3116_p2;
wire   [15:0] sub_ln703_312_fu_2993_p2;
wire   [15:0] add_ln703_403_fu_3131_p2;
wire   [15:0] sub_ln703_314_fu_3003_p2;
wire   [15:0] add_ln703_406_fu_3145_p2;
wire   [15:0] sub_ln703_316_fu_3026_p2;
wire   [15:0] sub_ln703_305_fu_2922_p2;
wire   [15:0] sub_ln703_288_fu_2854_p2;
wire   [15:0] add_ln703_414_fu_3165_p2;
wire   [15:0] sub_ln703_318_fu_3036_p2;
wire   [15:0] add_ln703_391_fu_3061_p2;
wire   [15:0] sub_ln703_321_fu_3066_p2;
wire   [15:0] sub_ln703_322_fu_3071_p2;
wire   [15:0] sub_ln703_323_fu_3076_p2;
wire   [15:0] add_ln703_394_fu_3086_p2;
wire   [15:0] sub_ln703_324_fu_3091_p2;
wire   [15:0] sub_ln703_325_fu_3096_p2;
wire   [15:0] sub_ln703_327_fu_3106_p2;
wire   [15:0] add_ln703_397_fu_3121_p2;
wire   [15:0] add_ln703_419_fu_3225_p2;
wire   [15:0] add_ln703_404_fu_3135_p2;
wire   [15:0] sub_ln703_331_fu_3140_p2;
wire   [15:0] add_ln703_413_fu_3160_p2;
wire   [15:0] sub_ln703_287_fu_2849_p2;
wire   [15:0] add_ln703_425_fu_3254_p2;
wire   [15:0] add_ln703_423_fu_3249_p2;
wire   [15:0] sub_ln703_317_fu_3031_p2;
wire   [15:0] sub_ln703_337_fu_3190_p2;
wire   [15:0] sub_ln703_338_fu_3195_p2;
wire   [15:0] sub_ln703_294_fu_2875_p2;
wire   [15:0] add_ln703_432_fu_3279_p2;
wire   [15:0] add_ln703_418_fu_3210_p2;
wire   [15:0] add_ln703_421_fu_3229_p2;
wire   [15:0] add_ln703_422_fu_3239_p2;
wire   [15:0] add_ln703_428_fu_3264_p2;
wire   [15:0] sub_ln703_320_fu_3056_p2;
wire   [15:0] sub_ln703_310_fu_2978_p2;
wire   [15:0] sub_ln703_357_fu_3295_p2;
wire   [15:0] sub_ln703_319_fu_3041_p2;
wire   [15:0] sub_ln703_329_fu_3126_p2;
wire   [15:0] sub_ln703_278_fu_2807_p2;
wire   [15:0] sub_ln703_332_fu_3376_p2;
wire   [15:0] add_ln703_411_fu_3380_p2;
wire   [15:0] sub_ln703_335_fu_3384_p2;
wire   [15:0] sub_ln703_346_fu_3396_p2;
wire   [15:0] sub_ln703_349_fu_3410_p2;
wire   [15:0] add_ln703_429_fu_3418_p2;
wire   [15:0] add_ln703_430_fu_3423_p2;
wire   [15:0] sub_ln703_352_fu_3427_p2;
wire   [15:0] sub_ln703_354_fu_3431_p2;
wire   [15:0] sub_ln703_355_fu_3435_p2;
wire   [15:0] sub_ln703_341_fu_3388_p2;
wire   [15:0] add_ln703_436_fu_3439_p2;
wire   [15:0] add_ln703_437_fu_3443_p2;
wire   [15:0] sub_ln703_348_fu_3405_p2;
wire   [15:0] sub_ln703_359_fu_3448_p2;
wire   [15:0] sub_ln703_360_fu_3453_p2;
wire   [15:0] sub_ln703_351_fu_3414_p2;
wire   [15:0] add_ln703_459_fu_3557_p2;
wire   [15:0] add_ln703_440_fu_3466_p2;
wire   [15:0] sub_ln703_364_fu_3470_p2;
wire   [15:0] add_ln703_441_fu_3480_p2;
wire   [15:0] sub_ln703_366_fu_3484_p2;
wire   [15:0] sub_ln703_367_fu_3488_p2;
wire   [15:0] sub_ln703_368_fu_3493_p2;
wire   [15:0] sub_ln703_369_fu_3497_p2;
wire   [15:0] add_ln703_442_fu_3502_p2;
wire   [15:0] add_ln703_444_fu_3506_p2;
wire   [15:0] add_ln703_448_fu_3511_p2;
wire   [15:0] sub_ln703_370_fu_3515_p2;
wire   [15:0] add_ln703_450_fu_3520_p2;
wire   [15:0] sub_ln703_330_fu_3372_p2;
wire   [15:0] add_ln703_467_fu_3635_p2;
wire   [15:0] add_ln703_465_fu_3630_p2;
wire   [15:0] add_ln703_452_fu_3524_p2;
wire   [15:0] add_ln703_453_fu_3528_p2;
wire   [15:0] sub_ln703_372_fu_3532_p2;
wire   [15:0] add_ln703_455_fu_3537_p2;
wire   [15:0] add_ln703_456_fu_3542_p2;
wire   [15:0] add_ln703_458_fu_3552_p2;
wire   [15:0] add_ln703_461_fu_3561_p2;
wire   [15:0] sub_ln703_363_fu_3461_p2;
wire   [15:0] add_ln703_462_fu_3571_p2;
wire   [15:0] sub_ln703_375_fu_3576_p2;
wire   [15:0] add_ln703_463_fu_3581_p2;
wire   [15:0] add_ln703_464_fu_3586_p2;
wire   [15:0] sub_ln703_377_fu_3596_p2;
wire   [15:0] sub_ln703_378_fu_3601_p2;
wire   [15:0] sub_ln703_379_fu_3606_p2;
wire   [15:0] sub_ln703_380_fu_3611_p2;
wire   [15:0] sub_ln703_381_fu_3616_p2;
wire   [15:0] sub_ln703_343_fu_3392_p2;
wire   [15:0] add_ln703_479_fu_3735_p2;
wire   [15:0] sub_ln703_382_fu_3621_p2;
wire   [15:0] sub_ln703_383_fu_3626_p2;
wire   [15:0] add_ln703_468_fu_3639_p2;
wire   [15:0] sub_ln703_385_fu_3650_p2;
wire   [15:0] sub_ln703_361_fu_3457_p2;
wire   [15:0] add_ln703_489_fu_3771_p2;
wire   [15:0] sub_ln703_388_fu_3670_p2;
wire   [15:0] sub_ln703_389_fu_3675_p2;
wire   [15:0] add_ln703_474_fu_3680_p2;
wire   [15:0] sub_ln703_374_fu_3566_p2;
wire   [15:0] sub_ln703_365_fu_3475_p2;
wire   [15:0] add_ln703_494_fu_3801_p2;
wire   [15:0] sub_ln703_391_fu_3695_p2;
wire   [15:0] sub_ln703_392_fu_3700_p2;
wire   [15:0] add_ln703_500_fu_3821_p2;
wire   [15:0] add_ln703_504_fu_3830_p2;
wire   [15:0] add_ln703_505_fu_3834_p2;
wire   [15:0] add_ln703_501_fu_3825_p2;
wire   [15:0] add_ln703_477_fu_3715_p2;
wire   [15:0] add_ln703_482_fu_3740_p2;
wire   [15:0] add_ln703_487_fu_3756_p2;
wire   [15:0] add_ln703_488_fu_3766_p2;
wire   [15:0] add_ln703_491_fu_3776_p2;
wire   [15:0] add_ln703_511_fu_3874_p2;
wire   [15:0] add_ln703_509_fu_3870_p2;
wire   [15:0] add_ln703_493_fu_3796_p2;
wire   [15:0] sub_ln703_396_fu_3725_p2;
wire   [15:0] sub_ln703_397_fu_3746_p2;
wire   [15:0] sub_ln703_398_fu_3751_p2;
wire   [15:0] add_ln703_536_fu_3908_p2;
wire   [15:0] add_ln703_532_fu_3904_p2;
wire   [15:0] sub_ln703_373_fu_3547_p2;
wire   [15:0] add_ln703_542_fu_3918_p2;
wire   [15:0] sub_ln703_376_fu_3591_p2;
wire   [15:0] add_ln703_553_fu_3928_p2;
wire   [15:0] add_ln703_519_fu_3899_p2;
wire   [15:0] sub_ln703_347_fu_3400_p2;
wire   [15:0] add_ln703_564_fu_3947_p2;
wire   [15:0] sub_ln703_400_fu_3973_p2;
wire   [15:0] sub_ln703_404_fu_3977_p2;
wire   [15:0] sub_ln703_407_fu_3985_p2;
wire   [15:0] sub_ln703_409_fu_3989_p2;
wire   [15:0] sub_ln703_410_fu_3993_p2;
wire   [15:0] sub_ln703_413_fu_3997_p2;
wire   [15:0] add_ln703_529_fu_4071_p2;
wire   [15:0] add_ln703_508_fu_4006_p2;
wire   [15:0] add_ln703_539_fu_4085_p2;
wire   [15:0] sub_ln703_417_fu_4010_p2;
wire   [15:0] sub_ln703_418_fu_4014_p2;
wire   [15:0] sub_ln703_420_fu_4019_p2;
wire   [15:0] sub_ln703_421_fu_4023_p2;
wire   [15:0] sub_ln703_422_fu_4027_p2;
wire   [15:0] sub_ln703_423_fu_4031_p2;
wire   [15:0] add_ln703_513_fu_4035_p2;
wire   [15:0] sub_ln703_424_fu_4040_p2;
wire   [15:0] sub_ln703_426_fu_4049_p2;
wire   [15:0] sub_ln703_427_fu_4054_p2;
wire   [15:0] add_ln703_520_fu_4058_p2;
wire   [15:0] add_ln703_521_fu_4062_p2;
wire   [15:0] add_ln703_522_fu_4067_p2;
wire   [15:0] add_ln703_538_fu_4075_p2;
wire   [15:0] sub_ln703_428_fu_4080_p2;
wire   [15:0] add_ln703_541_fu_4089_p2;
wire   [15:0] add_ln703_546_fu_4094_p2;
wire   [15:0] add_ln703_548_fu_4098_p2;
wire   [15:0] sub_ln703_429_fu_4102_p2;
wire   [15:0] sub_ln703_430_fu_4106_p2;
wire   [15:0] add_ln703_550_fu_4111_p2;
wire   [15:0] add_ln703_551_fu_4115_p2;
wire   [15:0] sub_ln703_431_fu_4120_p2;
wire   [15:0] sub_ln703_432_fu_4124_p2;
wire   [15:0] add_ln703_552_fu_4139_p2;
wire   [15:0] sub_ln703_436_fu_4149_p2;
wire   [15:0] sub_ln703_425_fu_4044_p2;
wire   [15:0] sub_ln703_437_fu_4154_p2;
wire   [15:0] add_ln703_557_fu_4158_p2;
wire   [15:0] sub_ln703_439_fu_4168_p2;
wire   [15:0] sub_ln703_441_fu_4172_p2;
wire   [15:0] sub_ln703_443_fu_4182_p2;
wire   [15:0] add_ln703_570_fu_4294_p2;
wire   [15:0] sub_ln703_445_fu_4192_p2;
wire   [15:0] sub_ln703_446_fu_4197_p2;
wire   [15:0] sub_ln703_447_fu_4202_p2;
wire   [15:0] add_ln703_558_fu_4216_p2;
wire   [15:0] sub_ln703_450_fu_4221_p2;
wire   [15:0] sub_ln703_451_fu_4226_p2;
wire   [15:0] add_ln703_559_fu_4241_p2;
wire   [15:0] sub_ln703_433_fu_4129_p2;
wire   [15:0] sub_ln703_406_fu_3981_p2;
wire   [15:0] add_ln703_577_fu_4343_p2;
wire   [15:0] sub_ln703_454_fu_4246_p2;
wire   [15:0] sub_ln703_455_fu_4251_p2;
wire   [15:0] sub_ln703_435_fu_4144_p2;
wire   [15:0] sub_ln703_456_fu_4255_p2;
wire   [15:0] add_ln703_561_fu_4260_p2;
wire   [15:0] sub_ln703_457_fu_4265_p2;
wire   [15:0] sub_ln703_438_fu_4163_p2;
wire   [15:0] add_ln703_562_fu_4275_p2;
wire   [15:0] add_ln703_563_fu_4280_p2;
wire   [15:0] sub_ln703_460_fu_4289_p2;
wire   [15:0] sub_ln703_415_fu_4001_p2;
wire   [15:0] add_ln703_589_fu_4408_p2;
wire   [15:0] add_ln703_587_fu_4403_p2;
wire   [15:0] add_ln703_571_fu_4298_p2;
wire   [15:0] sub_ln703_464_fu_4318_p2;
wire   [15:0] sub_ln703_465_fu_4328_p2;
wire   [15:0] add_ln703_597_fu_4437_p2;
wire   [15:0] add_ln703_594_fu_4433_p2;
wire   [15:0] add_ln703_576_fu_4338_p2;
wire   [15:0] add_ln703_580_fu_4348_p2;
wire   [15:0] sub_ln703_471_fu_4378_p2;
wire   [15:0] add_ln703_585_fu_4383_p2;
wire   [15:0] sub_ln703_473_fu_4388_p2;
wire   [15:0] sub_ln703_474_fu_4393_p2;
wire   [15:0] sub_ln703_442_fu_4177_p2;
wire   [15:0] add_ln703_602_fu_4482_p2;
wire   [15:0] add_ln703_607_fu_4491_p2;
wire   [15:0] add_ln703_604_fu_4486_p2;
wire   [15:0] sub_ln703_444_fu_4187_p2;
wire   [15:0] sub_ln703_449_fu_4211_p2;
wire   [15:0] add_ln703_614_fu_4506_p2;
wire   [15:0] sub_ln703_492_fu_4472_p2;
wire   [15:0] add_ln703_608_fu_4495_p2;
wire   [15:0] sub_ln703_434_fu_4134_p2;
wire   [15:0] add_ln703_631_fu_4526_p2;
wire   [15:0] sub_ln703_459_fu_4284_p2;
wire   [15:0] add_ln703_574_fu_4566_p2;
wire   [15:0] sub_ln703_472_fu_4570_p2;
wire   [15:0] sub_ln703_477_fu_4578_p2;
wire   [15:0] sub_ln703_478_fu_4582_p2;
wire   [15:0] sub_ln703_479_fu_4586_p2;
wire   [15:0] sub_ln703_480_fu_4590_p2;
wire   [15:0] sub_ln703_481_fu_4595_p2;
wire   [15:0] sub_ln703_484_fu_4599_p2;
wire   [15:0] sub_ln703_485_fu_4603_p2;
wire   [15:0] sub_ln703_486_fu_4607_p2;
wire   [15:0] add_ln703_601_fu_4620_p2;
wire   [15:0] sub_ln703_493_fu_4624_p2;
wire   [15:0] add_ln703_611_fu_4628_p2;
wire   [15:0] sub_ln703_494_fu_4632_p2;
wire   [15:0] sub_ln703_476_fu_4574_p2;
wire   [15:0] add_ln703_612_fu_4640_p2;
wire   [15:0] add_ln703_613_fu_4645_p2;
wire   [15:0] sub_ln703_496_fu_4650_p2;
wire   [15:0] sub_ln703_497_fu_4654_p2;
wire   [15:0] sub_ln703_498_fu_4659_p2;
wire   [15:0] sub_ln703_466_fu_4562_p2;
wire   [15:0] add_ln703_624_fu_4754_p2;
wire   [15:0] sub_ln703_500_fu_4668_p2;
wire   [15:0] sub_ln703_501_fu_4672_p2;
wire   [15:0] add_ln703_617_fu_4677_p2;
wire   [15:0] sub_ln703_502_fu_4682_p2;
wire   [15:0] add_ln703_618_fu_4687_p2;
wire   [15:0] sub_ln703_487_fu_4611_p2;
wire   [15:0] add_ln703_619_fu_4692_p2;
wire   [15:0] sub_ln703_489_fu_4615_p2;
wire   [15:0] add_ln703_620_fu_4696_p2;
wire   [15:0] sub_ln703_504_fu_4700_p2;
wire   [15:0] sub_ln703_506_fu_4705_p2;
wire   [15:0] sub_ln703_507_fu_4710_p2;
wire   [15:0] sub_ln703_508_fu_4715_p2;
wire   [15:0] add_ln703_622_fu_4720_p2;
wire   [15:0] sub_ln703_511_fu_4735_p2;
wire   [15:0] add_ln703_623_fu_4739_p2;
wire   [15:0] sub_ln703_512_fu_4744_p2;
wire   [15:0] add_ln703_626_fu_4759_p2;
wire   [15:0] sub_ln703_499_fu_4663_p2;
wire   [15:0] sub_ln703_514_fu_4764_p2;
wire   [15:0] add_ln703_627_fu_4769_p2;
wire   [15:0] add_ln703_629_fu_4774_p2;
wire   [15:0] sub_ln703_515_fu_4778_p2;
wire   [15:0] sub_ln703_516_fu_4783_p2;
wire   [15:0] sub_ln703_517_fu_4788_p2;
wire   [15:0] add_ln703_636_fu_4793_p2;
wire   [15:0] sub_ln703_518_fu_4798_p2;
wire   [15:0] add_ln703_638_fu_4803_p2;
wire   [15:0] sub_ln703_520_fu_4813_p2;
wire   [15:0] add_ln703_642_fu_4817_p2;
wire   [15:0] add_ln703_643_fu_4821_p2;
wire   [15:0] add_ln703_644_fu_4826_p2;
wire   [15:0] add_ln703_645_fu_4835_p2;
wire   [15:0] sub_ln703_522_fu_4840_p2;
wire   [15:0] sub_ln703_523_fu_4845_p2;
wire   [15:0] sub_ln703_510_fu_4730_p2;
wire   [15:0] sub_ln703_463_fu_4558_p2;
wire   [15:0] add_ln703_655_fu_4969_p2;
wire   [15:0] add_ln703_653_fu_4964_p2;
wire   [15:0] sub_ln703_524_fu_4850_p2;
wire   [15:0] sub_ln703_525_fu_4855_p2;
wire   [15:0] sub_ln703_513_fu_4749_p2;
wire   [15:0] sub_ln703_531_fu_4890_p2;
wire   [15:0] sub_ln703_534_fu_4909_p2;
wire   [15:0] add_ln703_649_fu_4914_p2;
wire   [15:0] add_ln703_663_fu_5009_p2;
wire   [15:0] sub_ln703_521_fu_4830_p2;
wire   [15:0] add_ln703_656_fu_4973_p2;
wire   [15:0] sub_ln703_543_fu_4979_p2;
wire   [15:0] add_ln703_658_fu_4989_p2;
wire   [15:0] sub_ln703_530_fu_4885_p2;
wire   [15:0] add_ln703_675_fu_5048_p2;
wire   [15:0] add_ln703_673_fu_5044_p2;
wire   [15:0] add_ln703_681_fu_5062_p2;
wire   [15:0] add_ln703_678_fu_5058_p2;
wire   [15:0] sub_ln703_519_fu_4808_p2;
wire   [15:0] add_ln703_683_fu_5072_p2;
wire   [15:0] sub_ln703_536_fu_4924_p2;
wire   [15:0] sub_ln703_537_fu_4929_p2;
wire   [15:0] sub_ln703_528_fu_4875_p2;
wire   [15:0] add_ln703_671_fu_5039_p2;
wire   [15:0] add_ln703_687_fu_5082_p2;
wire   [15:0] add_ln703_689_fu_5087_p2;
wire   [15:0] sub_ln703_509_fu_4725_p2;
wire   [15:0] sub_ln703_495_fu_4636_p2;
wire   [15:0] sub_ln703_546_fu_5142_p2;
wire   [15:0] sub_ln703_547_fu_5146_p2;
wire   [15:0] add_ln703_659_fu_5150_p2;
wire   [15:0] sub_ln703_548_fu_5154_p2;
wire   [15:0] sub_ln703_550_fu_5162_p2;
wire   [15:0] add_ln703_662_fu_5166_p2;
wire   [15:0] sub_ln703_553_fu_5174_p2;
wire   [15:0] sub_ln703_554_fu_5178_p2;
wire   [15:0] sub_ln703_555_fu_5182_p2;
wire   [15:0] add_ln703_669_fu_5186_p2;
wire   [15:0] sub_ln703_560_fu_5195_p2;
wire   [15:0] sub_ln703_561_fu_5200_p2;
wire   [15:0] sub_ln703_562_fu_5205_p2;
wire   [15:0] sub_ln703_564_fu_5214_p2;
wire   [15:0] sub_ln703_565_fu_5219_p2;
wire   [15:0] sub_ln703_566_fu_5223_p2;
wire   [15:0] sub_ln703_567_fu_5227_p2;
wire   [15:0] sub_ln703_568_fu_5232_p2;
wire   [15:0] add_ln703_702_fu_5332_p2;
wire   [15:0] sub_ln703_569_fu_5236_p2;
wire   [15:0] add_ln703_690_fu_5240_p2;
wire   [15:0] add_ln703_692_fu_5245_p2;
wire   [15:0] add_ln703_693_fu_5249_p2;
wire   [15:0] add_ln703_708_fu_5361_p2;
wire   [15:0] add_ln703_694_fu_5254_p2;
wire   [15:0] add_ln703_695_fu_5259_p2;
wire   [15:0] sub_ln703_570_fu_5263_p2;
wire   [15:0] sub_ln703_571_fu_5267_p2;
wire   [15:0] sub_ln703_545_fu_5138_p2;
wire   [15:0] add_ln703_710_fu_5390_p2;
wire   [15:0] add_ln703_696_fu_5272_p2;
wire   [15:0] sub_ln703_559_fu_5190_p2;
wire   [15:0] sub_ln703_572_fu_5276_p2;
wire   [15:0] add_ln703_699_fu_5281_p2;
wire   [15:0] add_ln703_700_fu_5285_p2;
wire   [15:0] sub_ln703_574_fu_5290_p2;
wire   [15:0] sub_ln703_563_fu_5209_p2;
wire   [15:0] sub_ln703_576_fu_5299_p2;
wire   [15:0] sub_ln703_577_fu_5304_p2;
wire   [15:0] add_ln703_701_fu_5313_p2;
wire   [15:0] sub_ln703_579_fu_5318_p2;
wire   [15:0] sub_ln703_580_fu_5323_p2;
wire   [15:0] sub_ln703_581_fu_5328_p2;
wire   [15:0] add_ln703_727_fu_5481_p2;
wire   [15:0] add_ln703_724_fu_5477_p2;
wire   [15:0] sub_ln703_587_fu_5356_p2;
wire   [15:0] add_ln703_709_fu_5365_p2;
wire   [15:0] sub_ln703_588_fu_5370_p2;
wire   [15:0] sub_ln703_590_fu_5380_p2;
wire   [15:0] sub_ln703_591_fu_5385_p2;
wire   [15:0] add_ln703_712_fu_5395_p2;
wire   [15:0] add_ln703_714_fu_5405_p2;
wire   [15:0] add_ln703_715_fu_5425_p2;
wire   [15:0] add_ln703_716_fu_5429_p2;
wire   [15:0] add_ln703_718_fu_5434_p2;
wire   [15:0] sub_ln703_596_fu_5444_p2;
wire   [15:0] sub_ln703_578_fu_5308_p2;
wire   [15:0] sub_ln703_597_fu_5449_p2;
wire   [15:0] sub_ln703_599_fu_5459_p2;
wire   [15:0] sub_ln703_600_fu_5464_p2;
wire   [15:0] add_ln703_720_fu_5469_p2;
wire   [15:0] sub_ln703_601_fu_5473_p2;
wire   [15:0] sub_ln703_552_fu_5170_p2;
wire   [15:0] add_ln703_738_fu_5581_p2;
wire   [15:0] add_ln703_736_fu_5576_p2;
wire   [15:0] sub_ln703_584_fu_5341_p2;
wire   [15:0] sub_ln703_607_fu_5506_p2;
wire   [15:0] sub_ln703_592_fu_5400_p2;
wire   [15:0] sub_ln703_575_fu_5295_p2;
wire   [15:0] add_ln703_745_fu_5606_p2;
wire   [15:0] sub_ln703_549_fu_5158_p2;
wire   [15:0] add_ln703_750_fu_5616_p2;
wire   [15:0] add_ln703_730_fu_5541_p2;
wire   [15:0] add_ln703_732_fu_5546_p2;
wire   [15:0] sub_ln703_617_fu_5561_p2;
wire   [15:0] add_ln703_739_fu_5585_p2;
wire   [15:0] add_ln703_741_fu_5591_p2;
wire   [15:0] add_ln703_744_fu_5601_p2;
wire   [15:0] add_ln703_747_fu_5611_p2;
wire   [15:0] add_ln703_753_fu_5621_p2;
wire   [15:0] sub_ln703_585_fu_5346_p2;
wire   [15:0] sub_ln703_602_fu_5688_p2;
wire   [15:0] add_ln703_721_fu_5692_p2;
wire   [15:0] add_ln703_729_fu_5700_p2;
wire   [15:0] sub_ln703_615_fu_5708_p2;
wire   [15:0] sub_ln703_619_fu_5716_p2;
wire   [15:0] sub_ln703_620_fu_5721_p2;
wire   [15:0] sub_ln703_622_fu_5730_p2;
wire   [15:0] sub_ln703_623_fu_5734_p2;
wire   [15:0] add_ln703_742_fu_5738_p2;
wire   [15:0] sub_ln703_606_fu_5696_p2;
wire   [15:0] sub_ln703_625_fu_5742_p2;
wire   [15:0] sub_ln703_626_fu_5746_p2;
wire   [15:0] sub_ln703_627_fu_5750_p2;
wire   [15:0] sub_ln703_611_fu_5704_p2;
wire   [15:0] sub_ln703_628_fu_5755_p2;
wire   [15:0] add_ln703_748_fu_5759_p2;
wire   [15:0] sub_ln703_629_fu_5763_p2;
wire   [15:0] sub_ln703_632_fu_5768_p2;
wire   [15:0] sub_ln703_633_fu_5772_p2;
wire   [15:0] add_ln703_754_fu_5776_p2;
wire   [15:0] sub_ln703_635_fu_5780_p2;
wire   [15:0] sub_ln703_621_fu_5726_p2;
wire   [15:0] sub_ln703_640_fu_5794_p2;
wire   [15:0] sub_ln703_642_fu_5804_p2;
wire   [15:0] add_ln703_756_fu_5809_p2;
wire   [15:0] add_ln703_757_fu_5814_p2;
wire   [15:0] add_ln703_759_fu_5818_p2;
wire   [15:0] sub_ln703_643_fu_5822_p2;
wire   [15:0] sub_ln703_646_fu_5832_p2;
wire   [15:0] add_ln703_761_fu_5837_p2;
wire   [15:0] add_ln703_769_fu_5946_p2;
wire   [15:0] add_ln703_767_fu_5942_p2;
wire   [15:0] add_ln703_763_fu_5842_p2;
wire   [15:0] sub_ln703_647_fu_5846_p2;
wire   [15:0] sub_ln703_649_fu_5851_p2;
wire   [15:0] sub_ln703_651_fu_5856_p2;
wire   [15:0] add_ln703_764_fu_5861_p2;
wire   [15:0] sub_ln703_652_fu_5865_p2;
wire   [15:0] sub_ln703_616_fu_5712_p2;
wire   [15:0] add_ln703_775_fu_5994_p2;
wire   [15:0] sub_ln703_653_fu_5870_p2;
wire   [15:0] sub_ln703_654_fu_5875_p2;
wire   [15:0] sub_ln703_655_fu_5879_p2;
wire   [15:0] sub_ln703_656_fu_5884_p2;
wire   [15:0] sub_ln703_636_fu_5784_p2;
wire   [15:0] sub_ln703_657_fu_5889_p2;
wire   [15:0] add_ln703_785_fu_6038_p2;
wire   [15:0] add_ln703_766_fu_5893_p2;
wire   [15:0] sub_ln703_658_fu_5898_p2;
wire   [15:0] sub_ln703_659_fu_5903_p2;
wire   [15:0] sub_ln703_660_fu_5908_p2;
wire   [15:0] sub_ln703_664_fu_5928_p2;
wire   [15:0] sub_ln703_666_fu_5937_p2;
wire   [15:0] add_ln703_771_fu_5961_p2;
wire   [15:0] add_ln703_772_fu_5966_p2;
wire   [15:0] sub_ln703_668_fu_5971_p2;
wire   [15:0] sub_ln703_670_fu_5980_p2;
wire   [15:0] add_ln703_774_fu_5985_p2;
wire   [15:0] sub_ln703_671_fu_5989_p2;
wire   [15:0] add_ln703_777_fu_5999_p2;
wire   [15:0] sub_ln703_672_fu_6004_p2;
wire   [15:0] sub_ln703_673_fu_6009_p2;
wire   [15:0] sub_ln703_674_fu_6014_p2;
wire   [15:0] sub_ln703_675_fu_6019_p2;
wire   [15:0] add_ln703_781_fu_6029_p2;
wire   [15:0] add_ln703_786_fu_6042_p2;
wire   [15:0] sub_ln703_677_fu_6047_p2;
wire   [15:0] sub_ln703_641_fu_5799_p2;
wire   [15:0] add_ln703_795_fu_6156_p2;
wire   [15:0] add_ln703_794_fu_6151_p2;
wire   [15:0] sub_ln703_663_fu_5923_p2;
wire   [15:0] add_ln703_788_fu_6082_p2;
wire   [15:0] sub_ln703_689_fu_6096_p2;
wire   [15:0] add_ln703_790_fu_6121_p2;
wire   [15:0] sub_ln703_639_fu_5789_p2;
wire   [15:0] sub_ln703_661_fu_5913_p2;
wire   [15:0] add_ln703_817_fu_6201_p2;
wire   [15:0] add_ln703_815_fu_6196_p2;
wire   [15:0] sub_ln703_645_fu_5827_p2;
wire   [15:0] add_ln703_820_fu_6211_p2;
wire   [15:0] sub_ln703_681_fu_6238_p2;
wire   [15:0] sub_ln703_683_fu_6242_p2;
wire   [15:0] sub_ln703_685_fu_6246_p2;
wire   [15:0] add_ln703_789_fu_6250_p2;
wire   [15:0] sub_ln703_695_fu_6254_p2;
wire   [15:0] add_ln703_803_fu_6319_p2;
wire   [15:0] add_ln703_793_fu_6258_p2;
wire   [15:0] add_ln703_797_fu_6262_p2;
wire   [15:0] sub_ln703_698_fu_6267_p2;
wire   [15:0] sub_ln703_699_fu_6271_p2;
wire   [15:0] add_ln703_799_fu_6276_p2;
wire   [15:0] add_ln703_807_fu_6369_p2;
wire   [15:0] sub_ln703_701_fu_6281_p2;
wire   [15:0] sub_ln703_702_fu_6285_p2;
wire   [15:0] sub_ln703_703_fu_6289_p2;
wire   [15:0] sub_ln703_708_fu_6302_p2;
wire   [15:0] sub_ln703_709_fu_6306_p2;
wire   [15:0] add_ln703_800_fu_6315_p2;
wire   [15:0] add_ln703_804_fu_6323_p2;
wire   [15:0] sub_ln703_713_fu_6337_p2;
wire   [15:0] add_ln703_805_fu_6341_p2;
wire   [15:0] sub_ln703_714_fu_6345_p2;
wire   [15:0] sub_ln703_715_fu_6350_p2;
wire   [15:0] add_ln703_806_fu_6359_p2;
wire   [15:0] add_ln703_808_fu_6373_p2;
wire   [15:0] add_ln703_809_fu_6378_p2;
wire   [15:0] sub_ln703_718_fu_6382_p2;
wire   [15:0] sub_ln703_719_fu_6386_p2;
wire   [15:0] sub_ln703_720_fu_6391_p2;
wire   [15:0] add_ln703_810_fu_6396_p2;
wire   [15:0] add_ln703_811_fu_6401_p2;
wire   [15:0] add_ln703_812_fu_6405_p2;
wire   [15:0] add_ln703_813_fu_6409_p2;
wire   [15:0] sub_ln703_721_fu_6413_p2;
wire   [15:0] add_ln703_823_fu_6512_p2;
wire   [15:0] add_ln703_814_fu_6417_p2;
wire   [15:0] sub_ln703_722_fu_6422_p2;
wire   [15:0] sub_ln703_710_fu_6311_p2;
wire   [15:0] sub_ln703_712_fu_6332_p2;
wire   [15:0] sub_ln703_725_fu_6437_p2;
wire   [15:0] add_ln703_830_fu_6550_p2;
wire   [15:0] add_ln703_829_fu_6546_p2;
wire   [15:0] sub_ln703_726_fu_6442_p2;
wire   [15:0] add_ln703_832_fu_6569_p2;
wire   [15:0] sub_ln703_729_fu_6462_p2;
wire   [15:0] sub_ln703_730_fu_6467_p2;
wire   [15:0] sub_ln703_731_fu_6472_p2;
wire   [15:0] sub_ln703_732_fu_6477_p2;
wire   [15:0] add_ln703_822_fu_6482_p2;
wire   [15:0] sub_ln703_734_fu_6492_p2;
wire   [15:0] sub_ln703_735_fu_6497_p2;
wire   [15:0] sub_ln703_737_fu_6507_p2;
wire   [15:0] add_ln703_824_fu_6516_p2;
wire   [15:0] sub_ln703_723_fu_6427_p2;
wire   [15:0] add_ln703_828_fu_6536_p2;
wire   [15:0] sub_ln703_739_fu_6541_p2;
wire   [15:0] sub_ln703_740_fu_6560_p2;
wire   [15:0] sub_ln703_744_fu_6565_p2;
wire   [15:0] sub_ln703_747_fu_6584_p2;
wire   [15:0] sub_ln703_748_fu_6589_p2;
wire   [15:0] sub_ln703_751_fu_6604_p2;
wire   [15:0] sub_ln703_752_fu_6609_p2;
wire   [15:0] sub_ln703_705_fu_6294_p2;
wire   [15:0] add_ln703_843_fu_6674_p2;
wire   [15:0] add_ln703_842_fu_6669_p2;
wire   [15:0] sub_ln703_753_fu_6614_p2;
wire   [15:0] sub_ln703_754_fu_6619_p2;
wire   [15:0] add_ln703_850_fu_6698_p2;
wire   [15:0] add_ln703_848_fu_6694_p2;
wire   [15:0] add_ln703_837_fu_6624_p2;
wire   [15:0] sub_ln703_711_fu_6328_p2;
wire   [15:0] add_ln703_853_fu_6718_p2;
wire   [15:0] add_ln703_852_fu_6713_p2;
wire   [15:0] sub_ln703_716_fu_6354_p2;
wire   [15:0] add_ln703_857_fu_6728_p2;
wire   [15:0] add_ln703_844_fu_6678_p2;
wire   [15:0] sub_ln703_706_fu_6298_p2;
wire   [15:0] add_ln703_863_fu_6744_p2;
wire   [15:0] add_ln703_854_fu_6722_p2;
wire   [15:0] add_ln703_864_fu_6749_p2;
wire   [15:0] sub_ln703_717_fu_6364_p2;
wire   [15:0] sub_ln703_738_fu_6521_p2;
wire   [15:0] sub_ln703_741_fu_6795_p2;
wire   [15:0] sub_ln703_743_fu_6803_p2;
wire   [15:0] sub_ln703_750_fu_6811_p2;
wire   [15:0] add_ln703_835_fu_6815_p2;
wire   [15:0] sub_ln703_755_fu_6819_p2;
wire   [15:0] sub_ln703_756_fu_6823_p2;
wire   [15:0] sub_ln703_758_fu_6827_p2;
wire   [15:0] sub_ln703_760_fu_6831_p2;
wire   [15:0] sub_ln703_742_fu_6799_p2;
wire   [15:0] add_ln703_839_fu_6836_p2;
wire   [15:0] sub_ln703_745_fu_6807_p2;
wire   [15:0] sub_ln703_762_fu_6841_p2;
wire   [15:0] sub_ln703_764_fu_6845_p2;
wire   [15:0] sub_ln703_765_fu_6849_p2;
wire   [15:0] sub_ln703_766_fu_6853_p2;
wire   [15:0] add_ln703_846_fu_6863_p2;
wire   [15:0] add_ln703_847_fu_6868_p2;
wire   [15:0] add_ln703_866_fu_6972_p2;
wire   [15:0] sub_ln703_772_fu_6877_p2;
wire   [15:0] add_ln703_855_fu_6882_p2;
wire   [15:0] add_ln703_856_fu_6891_p2;
wire   [15:0] add_ln703_859_fu_6901_p2;
wire   [15:0] add_ln703_860_fu_6905_p2;
wire   [15:0] sub_ln703_775_fu_6910_p2;
wire   [15:0] add_ln703_861_fu_6919_p2;
wire   [15:0] add_ln703_862_fu_6923_p2;
wire   [15:0] sub_ln703_777_fu_6928_p2;
wire   [15:0] sub_ln703_778_fu_6933_p2;
wire   [15:0] sub_ln703_779_fu_6938_p2;
wire   [15:0] sub_ln703_782_fu_6946_p2;
wire   [15:0] sub_ln703_783_fu_6950_p2;
wire   [15:0] sub_ln703_784_fu_6954_p2;
wire   [15:0] sub_ln703_785_fu_6959_p2;
wire   [15:0] sub_ln703_786_fu_6964_p2;
wire   [15:0] add_ln703_865_fu_6968_p2;
wire   [15:0] add_ln703_869_fu_6976_p2;
wire   [15:0] sub_ln703_790_fu_6991_p2;
wire   [15:0] sub_ln703_791_fu_6996_p2;
wire   [15:0] sub_ln703_792_fu_7000_p2;
wire   [15:0] sub_ln703_793_fu_7005_p2;
wire   [15:0] sub_ln703_794_fu_7010_p2;
wire   [15:0] add_ln703_878_fu_7104_p2;
wire   [15:0] add_ln703_881_fu_7117_p2;
wire   [15:0] add_ln703_880_fu_7113_p2;
wire   [15:0] sub_ln703_795_fu_7015_p2;
wire   [15:0] sub_ln703_796_fu_7020_p2;
wire   [15:0] add_ln703_870_fu_7025_p2;
wire   [15:0] sub_ln703_798_fu_7035_p2;
wire   [15:0] sub_ln703_768_fu_6858_p2;
wire   [15:0] add_ln703_887_fu_7151_p2;
wire   [15:0] add_ln703_871_fu_7040_p2;
wire   [15:0] sub_ln703_800_fu_7045_p2;
wire   [15:0] sub_ln703_803_fu_7070_p2;
wire   [15:0] sub_ln703_804_fu_7075_p2;
wire   [15:0] sub_ln703_788_fu_6981_p2;
wire   [15:0] sub_ln703_773_fu_6886_p2;
wire   [15:0] sub_ln703_774_fu_6896_p2;
wire   [15:0] sub_ln703_806_fu_7089_p2;
wire   [15:0] add_ln703_879_fu_7108_p2;
wire   [15:0] add_ln703_883_fu_7127_p2;
wire   [15:0] add_ln703_885_fu_7142_p2;
wire   [15:0] add_ln703_886_fu_7147_p2;
wire   [15:0] add_ln703_889_fu_7161_p2;
wire   [15:0] sub_ln703_809_fu_7165_p2;
wire   [15:0] sub_ln703_810_fu_7170_p2;
wire   [15:0] sub_ln703_789_fu_6986_p2;
wire   [15:0] add_ln703_904_fu_7240_p2;
wire   [15:0] sub_ln703_780_fu_6942_p2;
wire   [15:0] add_ln703_909_fu_7255_p2;
wire   [15:0] add_ln703_908_fu_7250_p2;
wire   [15:0] add_ln703_916_fu_7269_p2;
wire   [15:0] add_ln703_915_fu_7265_p2;
wire   [15:0] add_ln703_921_fu_7283_p2;
wire   [15:0] add_ln703_919_fu_7279_p2;
wire   [15:0] sub_ln703_771_fu_6873_p2;
wire   [15:0] add_ln703_924_fu_7298_p2;
wire   [15:0] add_ln703_923_fu_7293_p2;
wire   [15:0] sub_ln703_776_fu_6915_p2;
wire   [15:0] add_ln703_931_fu_7308_p2;
wire   [15:0] add_ln703_910_fu_7259_p2;
wire   [15:0] add_ln703_925_fu_7302_p2;
wire   [15:0] add_ln703_932_fu_7313_p2;
wire   [15:0] sub_ln703_811_fu_7346_p2;
wire   [15:0] sub_ln703_812_fu_7350_p2;
wire   [15:0] add_ln703_890_fu_7354_p2;
wire   [15:0] add_ln703_891_fu_7358_p2;
wire   [15:0] add_ln703_897_fu_7362_p2;
wire   [15:0] add_ln703_899_fu_7366_p2;
wire   [15:0] sub_ln703_813_fu_7370_p2;
wire   [15:0] sub_ln703_815_fu_7374_p2;
wire   [15:0] add_ln703_900_fu_7378_p2;
wire   [15:0] add_ln703_901_fu_7390_p2;
wire   [15:0] add_ln703_902_fu_7394_p2;
wire   [15:0] sub_ln703_822_fu_7398_p2;
wire   [15:0] add_ln703_903_fu_7402_p2;
wire   [15:0] sub_ln703_826_fu_7407_p2;
wire   [15:0] sub_ln703_827_fu_7412_p2;
wire   [15:0] sub_ln703_828_fu_7417_p2;
wire   [15:0] sub_ln703_829_fu_7422_p2;
wire   [15:0] sub_ln703_831_fu_7430_p2;
wire   [15:0] sub_ln703_832_fu_7434_p2;
wire   [15:0] add_ln703_927_fu_7537_p2;
wire   [15:0] sub_ln703_833_fu_7439_p2;
wire   [15:0] sub_ln703_834_fu_7444_p2;
wire   [15:0] sub_ln703_836_fu_7453_p2;
wire   [15:0] sub_ln703_837_fu_7458_p2;
wire   [15:0] sub_ln703_839_fu_7467_p2;
wire   [15:0] add_ln703_907_fu_7477_p2;
wire   [15:0] add_ln703_911_fu_7481_p2;
wire   [15:0] sub_ln703_841_fu_7485_p2;
wire   [15:0] add_ln703_912_fu_7490_p2;
wire   [15:0] add_ln703_913_fu_7494_p2;
wire   [15:0] sub_ln703_842_fu_7498_p2;
wire   [15:0] sub_ln703_843_fu_7503_p2;
wire   [15:0] sub_ln703_844_fu_7508_p2;
wire   [15:0] add_ln703_918_fu_7513_p2;
wire   [15:0] sub_ln703_845_fu_7518_p2;
wire   [15:0] sub_ln703_846_fu_7523_p2;
wire   [15:0] sub_ln703_847_fu_7528_p2;
wire   [15:0] add_ln703_926_fu_7532_p2;
wire   [15:0] add_ln703_928_fu_7541_p2;
wire   [15:0] add_ln703_929_fu_7546_p2;
wire   [15:0] sub_ln703_848_fu_7551_p2;
wire   [15:0] add_ln703_937_fu_7659_p2;
wire   [15:0] sub_ln703_835_fu_7449_p2;
wire   [15:0] sub_ln703_849_fu_7556_p2;
wire   [15:0] add_ln703_930_fu_7561_p2;
wire   [15:0] sub_ln703_838_fu_7463_p2;
wire   [15:0] sub_ln703_850_fu_7566_p2;
wire   [15:0] sub_ln703_840_fu_7472_p2;
wire   [15:0] sub_ln703_851_fu_7571_p2;
wire   [15:0] sub_ln703_853_fu_7576_p2;
wire   [15:0] add_ln703_933_fu_7581_p2;
wire   [15:0] add_ln703_942_fu_7715_p2;
wire   [15:0] sub_ln703_855_fu_7591_p2;
wire   [15:0] sub_ln703_856_fu_7596_p2;
wire   [15:0] sub_ln703_860_fu_7620_p2;
wire   [15:0] sub_ln703_830_fu_7426_p2;
wire   [15:0] add_ln703_945_fu_7740_p2;
wire   [15:0] sub_ln703_861_fu_7625_p2;
wire   [15:0] add_ln703_935_fu_7629_p2;
wire   [15:0] sub_ln703_864_fu_7644_p2;
wire   [15:0] sub_ln703_817_fu_7382_p2;
wire   [15:0] add_ln703_950_fu_7770_p2;
wire   [15:0] add_ln703_949_fu_7765_p2;
wire   [15:0] add_ln703_940_fu_7690_p2;
wire   [15:0] sub_ln703_871_fu_7696_p2;
wire   [15:0] add_ln703_941_fu_7701_p2;
wire   [15:0] sub_ln703_872_fu_7705_p2;
wire   [15:0] sub_ln703_854_fu_7586_p2;
wire   [15:0] sub_ln703_874_fu_7725_p2;
wire   [15:0] add_ln703_947_fu_7745_p2;
wire   [15:0] add_ln703_957_fu_7823_p2;
wire   [15:0] add_ln703_956_fu_7819_p2;
wire   [15:0] add_ln703_951_fu_7774_p2;
wire   [15:0] add_ln703_952_fu_7800_p2;
wire   [15:0] add_ln703_955_fu_7815_p2;
wire   [15:0] sub_ln703_819_fu_7386_p2;
wire   [15:0] add_ln703_1000_fu_7852_p2;
wire   [15:0] add_ln703_1002_fu_7863_p2;
wire   [15:0] add_ln703_1003_fu_7867_p2;
wire   [15:0] add_ln703_1001_fu_7857_p2;
wire   [15:0] sub_ln703_876_fu_7878_p2;
wire   [15:0] add_ln703_944_fu_7882_p2;
wire   [15:0] sub_ln703_877_fu_7886_p2;
wire   [15:0] sub_ln703_878_fu_7890_p2;
wire   [15:0] sub_ln703_883_fu_7898_p2;
wire   [15:0] sub_ln703_885_fu_7906_p2;
wire   [15:0] sub_ln703_888_fu_7918_p2;
wire   [15:0] sub_ln703_889_fu_7922_p2;
wire   [15:0] sub_ln703_890_fu_7926_p2;
wire   [15:0] sub_ln703_891_fu_7930_p2;
wire   [15:0] sub_ln703_896_fu_7934_p2;
wire   [15:0] add_ln703_953_fu_7956_p2;
wire   [15:0] sub_ln703_902_fu_7961_p2;
wire   [15:0] sub_ln703_903_fu_7966_p2;
wire   [15:0] sub_ln703_905_fu_7970_p2;
wire   [15:0] sub_ln703_906_fu_7974_p2;
wire   [15:0] sub_ln703_908_fu_7983_p2;
wire   [15:0] sub_ln703_886_fu_7910_p2;
wire   [15:0] add_ln703_959_fu_7997_p2;
wire   [15:0] sub_ln703_913_fu_8007_p2;
wire   [15:0] add_ln703_960_fu_8012_p2;
wire   [15:0] add_ln703_961_fu_8016_p2;
wire   [15:0] sub_ln703_914_fu_8020_p2;
wire   [15:0] sub_ln703_915_fu_8024_p2;
wire   [15:0] sub_ln703_897_fu_7938_p2;
wire   [15:0] sub_ln703_918_fu_8033_p2;
wire   [15:0] sub_ln703_921_fu_8047_p2;
wire   [15:0] add_ln703_970_fu_8125_p2;
wire   [15:0] add_ln703_962_fu_8052_p2;
wire   [15:0] sub_ln703_923_fu_8057_p2;
wire   [15:0] sub_ln703_882_fu_7894_p2;
wire   [15:0] add_ln703_972_fu_8148_p2;
wire   [15:0] sub_ln703_907_fu_7978_p2;
wire   [15:0] add_ln703_963_fu_8062_p2;
wire   [15:0] sub_ln703_884_fu_7902_p2;
wire   [15:0] add_ln703_975_fu_8170_p2;
wire   [15:0] add_ln703_965_fu_8067_p2;
wire   [15:0] sub_ln703_887_fu_7914_p2;
wire   [15:0] add_ln703_977_fu_8186_p2;
wire   [15:0] sub_ln703_910_fu_7992_p2;
wire   [15:0] sub_ln703_912_fu_8002_p2;
wire   [15:0] sub_ln703_928_fu_8090_p2;
wire   [15:0] sub_ln703_929_fu_8095_p2;
wire   [15:0] add_ln703_966_fu_8100_p2;
wire   [15:0] add_ln703_967_fu_8105_p2;
wire   [15:0] add_ln703_968_fu_8110_p2;
wire   [15:0] add_ln703_969_fu_8115_p2;
wire   [15:0] sub_ln703_899_fu_7942_p2;
wire   [15:0] add_ln703_982_fu_8239_p2;
wire   [15:0] sub_ln703_900_fu_7946_p2;
wire   [15:0] add_ln703_984_fu_8250_p2;
wire   [15:0] sub_ln703_901_fu_7951_p2;
wire   [15:0] add_ln703_987_fu_8260_p2;
wire   [15:0] sub_ln703_919_fu_8037_p2;
wire   [15:0] sub_ln703_920_fu_8042_p2;
wire   [15:0] sub_ln703_930_fu_8120_p2;
wire   [15:0] add_ln703_971_fu_8129_p2;
wire   [15:0] sub_ln703_931_fu_8134_p2;
wire   [15:0] sub_ln703_932_fu_8139_p2;
wire   [15:0] sub_ln703_933_fu_8143_p2;
wire   [15:0] add_ln703_973_fu_8153_p2;
wire   [15:0] add_ln703_974_fu_8159_p2;
wire   [15:0] sub_ln703_934_fu_8165_p2;
wire   [15:0] add_ln703_976_fu_8175_p2;
wire   [15:0] sub_ln703_909_fu_7987_p2;
wire   [15:0] add_ln703_994_fu_8325_p2;
wire   [15:0] sub_ln703_935_fu_8181_p2;
wire   [15:0] add_ln703_978_fu_8191_p2;
wire   [15:0] add_ln703_979_fu_8197_p2;
wire   [15:0] sub_ln703_924_fu_8072_p2;
wire   [15:0] sub_ln703_925_fu_8076_p2;
wire   [15:0] sub_ln703_926_fu_8080_p2;
wire   [15:0] add_ln703_980_fu_8203_p2;
wire   [15:0] sub_ln703_927_fu_8085_p2;
wire   [15:0] sub_ln703_936_fu_8209_p2;
wire   [15:0] add_ln703_981_fu_8214_p2;
wire   [15:0] sub_ln703_937_fu_8219_p2;
wire   [15:0] sub_ln703_938_fu_8224_p2;
wire   [15:0] sub_ln703_916_fu_8028_p2;
wire   [15:0] add_ln703_1007_fu_8395_p2;
wire   [15:0] sub_ln703_939_fu_8229_p2;
wire   [15:0] add_ln703_1009_fu_8410_p2;
wire   [15:0] sub_ln703_940_fu_8234_p2;
wire   [15:0] add_ln703_983_fu_8244_p2;
wire   [15:0] add_ln703_986_fu_8255_p2;
wire   [15:0] acc_1_V_fu_8265_p2;
wire   [15:0] acc_2_V_fu_8270_p2;
wire   [15:0] acc_3_V_fu_8275_p2;
wire   [15:0] acc_4_V_fu_8280_p2;
wire   [15:0] acc_5_V_fu_8285_p2;
wire   [15:0] acc_6_V_fu_8290_p2;
wire   [15:0] acc_7_V_fu_8295_p2;
wire   [15:0] acc_8_V_fu_8300_p2;
wire   [15:0] acc_9_V_fu_8305_p2;
wire   [15:0] acc_10_V_fu_8310_p2;
wire   [15:0] acc_11_V_fu_8315_p2;
wire   [15:0] acc_12_V_fu_8320_p2;
wire   [15:0] acc_13_V_fu_8330_p2;
wire   [15:0] acc_14_V_fu_8335_p2;
wire   [15:0] acc_15_V_fu_8340_p2;
wire   [15:0] acc_16_V_fu_8345_p2;
wire   [15:0] acc_17_V_fu_8350_p2;
wire   [15:0] acc_18_V_fu_8355_p2;
wire   [15:0] acc_19_V_fu_8360_p2;
wire   [15:0] acc_20_V_fu_8365_p2;
wire   [15:0] acc_22_V_fu_8370_p2;
wire   [15:0] acc_23_V_fu_8375_p2;
wire   [15:0] acc_24_V_fu_8380_p2;
wire   [15:0] acc_25_V_fu_8385_p2;
wire   [15:0] acc_26_V_fu_8390_p2;
wire   [15:0] acc_27_V_fu_8400_p2;
wire   [15:0] acc_28_V_fu_8405_p2;
wire   [15:0] acc_29_V_fu_8414_p2;
wire   [15:0] acc_30_V_fu_8419_p2;
wire   [15:0] acc_31_V_fu_8424_p2;
reg    ap_ce_reg;
reg   [15:0] data_0_V_read_int_reg;
reg   [15:0] data_1_V_read_int_reg;
reg   [15:0] data_2_V_read_int_reg;
reg   [15:0] data_3_V_read_int_reg;
reg   [15:0] data_4_V_read_int_reg;
reg   [15:0] data_5_V_read_int_reg;
reg   [15:0] data_6_V_read_int_reg;
reg   [15:0] data_7_V_read_int_reg;
reg   [15:0] data_8_V_read_int_reg;
reg   [15:0] data_9_V_read_int_reg;
reg   [15:0] data_10_V_read_int_reg;
reg   [15:0] data_11_V_read_int_reg;
reg   [15:0] data_12_V_read_int_reg;
reg   [15:0] data_13_V_read_int_reg;
reg   [15:0] data_14_V_read_int_reg;
reg   [15:0] data_15_V_read_int_reg;
reg   [15:0] data_16_V_read_int_reg;
reg   [15:0] data_17_V_read_int_reg;
reg   [15:0] data_18_V_read_int_reg;
reg   [15:0] data_19_V_read_int_reg;
reg   [15:0] data_20_V_read_int_reg;
reg   [15:0] data_21_V_read_int_reg;
reg   [15:0] data_22_V_read_int_reg;
reg   [15:0] data_23_V_read_int_reg;
reg   [15:0] data_24_V_read_int_reg;
reg   [15:0] data_25_V_read_int_reg;
reg   [15:0] data_26_V_read_int_reg;
reg   [15:0] data_27_V_read_int_reg;
reg   [15:0] data_28_V_read_int_reg;
reg   [15:0] data_29_V_read_int_reg;
reg   [15:0] data_30_V_read_int_reg;
reg   [15:0] data_31_V_read_int_reg;
reg   [15:0] data_32_V_read_int_reg;
reg   [15:0] data_33_V_read_int_reg;
reg   [15:0] data_34_V_read_int_reg;
reg   [15:0] data_35_V_read_int_reg;
reg   [15:0] data_36_V_read_int_reg;
reg   [15:0] data_37_V_read_int_reg;
reg   [15:0] data_38_V_read_int_reg;
reg   [15:0] data_39_V_read_int_reg;
reg   [15:0] data_40_V_read_int_reg;
reg   [15:0] data_41_V_read_int_reg;
reg   [15:0] data_42_V_read_int_reg;
reg   [15:0] data_43_V_read_int_reg;
reg   [15:0] data_44_V_read_int_reg;
reg   [15:0] data_45_V_read_int_reg;
reg   [15:0] data_46_V_read_int_reg;
reg   [15:0] data_47_V_read_int_reg;
reg   [15:0] data_48_V_read_int_reg;
reg   [15:0] data_49_V_read_int_reg;
reg   [15:0] data_50_V_read_int_reg;
reg   [15:0] data_51_V_read_int_reg;
reg   [15:0] data_52_V_read_int_reg;
reg   [15:0] data_53_V_read_int_reg;
reg   [15:0] data_54_V_read_int_reg;
reg   [15:0] data_55_V_read_int_reg;
reg   [15:0] data_56_V_read_int_reg;
reg   [15:0] data_57_V_read_int_reg;
reg   [15:0] data_58_V_read_int_reg;
reg   [15:0] data_59_V_read_int_reg;
reg   [15:0] data_60_V_read_int_reg;
reg   [15:0] data_61_V_read_int_reg;
reg   [15:0] data_62_V_read_int_reg;
reg   [15:0] data_63_V_read_int_reg;
reg   [15:0] ap_return_0_int_reg;
reg   [15:0] ap_return_1_int_reg;
reg   [15:0] ap_return_2_int_reg;
reg   [15:0] ap_return_3_int_reg;
reg   [15:0] ap_return_4_int_reg;
reg   [15:0] ap_return_5_int_reg;
reg   [15:0] ap_return_6_int_reg;
reg   [15:0] ap_return_7_int_reg;
reg   [15:0] ap_return_8_int_reg;
reg   [15:0] ap_return_9_int_reg;
reg   [15:0] ap_return_10_int_reg;
reg   [15:0] ap_return_11_int_reg;
reg   [15:0] ap_return_12_int_reg;
reg   [15:0] ap_return_13_int_reg;
reg   [15:0] ap_return_14_int_reg;
reg   [15:0] ap_return_15_int_reg;
reg   [15:0] ap_return_16_int_reg;
reg   [15:0] ap_return_17_int_reg;
reg   [15:0] ap_return_18_int_reg;
reg   [15:0] ap_return_19_int_reg;
reg   [15:0] ap_return_20_int_reg;
reg   [15:0] ap_return_21_int_reg;
reg   [15:0] ap_return_22_int_reg;
reg   [15:0] ap_return_23_int_reg;
reg   [15:0] ap_return_24_int_reg;
reg   [15:0] ap_return_25_int_reg;
reg   [15:0] ap_return_26_int_reg;
reg   [15:0] ap_return_27_int_reg;
reg   [15:0] ap_return_28_int_reg;
reg   [15:0] ap_return_29_int_reg;
reg   [15:0] ap_return_30_int_reg;
reg   [15:0] ap_return_31_int_reg;

always @ (posedge ap_clk) begin
    ap_ce_reg <= ap_ce;
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        acc_21_V_reg_12991 <= acc_21_V_fu_7872_p2;
        add_ln703_130_reg_10373 <= add_ln703_130_fu_556_p2;
        add_ln703_131_reg_10354 <= add_ln703_131_fu_544_p2;
        add_ln703_131_reg_10354_pp0_iter2_reg <= add_ln703_131_reg_10354;
        add_ln703_132_reg_10414 <= add_ln703_132_fu_599_p2;
        add_ln703_134_reg_10385 <= add_ln703_134_fu_568_p2;
        add_ln703_135_reg_10425 <= add_ln703_135_fu_619_p2;
        add_ln703_140_reg_10442 <= add_ln703_140_fu_644_p2;
        add_ln703_141_reg_10447 <= add_ln703_141_fu_649_p2;
        add_ln703_144_reg_10403 <= add_ln703_144_fu_589_p2;
        add_ln703_144_reg_10403_pp0_iter3_reg <= add_ln703_144_reg_10403;
        add_ln703_153_reg_10503 <= add_ln703_153_fu_809_p2;
        add_ln703_157_reg_10529 <= add_ln703_157_fu_892_p2;
        add_ln703_158_reg_10482 <= add_ln703_158_fu_676_p2;
        add_ln703_161_reg_10487 <= add_ln703_161_fu_681_p2;
        add_ln703_162_reg_10539 <= add_ln703_162_fu_917_p2;
        add_ln703_170_reg_10566 <= add_ln703_170_fu_972_p2;
        add_ln703_171_reg_10571 <= add_ln703_171_fu_977_p2;
        add_ln703_173_reg_10576 <= add_ln703_173_fu_982_p2;
        add_ln703_177_reg_10591 <= add_ln703_177_fu_997_p2;
        add_ln703_179_reg_10495 <= add_ln703_179_fu_685_p2;
        add_ln703_181_reg_10601 <= add_ln703_181_fu_1015_p2;
        add_ln703_183_reg_10606 <= add_ln703_183_fu_1021_p2;
        add_ln703_186_reg_10621 <= add_ln703_186_fu_1036_p2;
        add_ln703_192_reg_10626 <= add_ln703_192_fu_1050_p2;
        add_ln703_204_reg_10641 <= add_ln703_204_fu_1059_p2;
        add_ln703_207_reg_10682 <= add_ln703_207_fu_1299_p2;
        add_ln703_208_reg_10687 <= add_ln703_208_fu_1309_p2;
        add_ln703_209_reg_10646 <= add_ln703_209_fu_1064_p2;
        add_ln703_210_reg_10692 <= add_ln703_210_fu_1314_p2;
        add_ln703_213_reg_10653 <= add_ln703_213_fu_1068_p2;
        add_ln703_216_reg_10702 <= add_ln703_216_fu_1358_p2;
        add_ln703_223_reg_10658 <= add_ln703_223_fu_1073_p2;
        add_ln703_224_reg_10732 <= add_ln703_224_fu_1437_p2;
        add_ln703_226_reg_10737 <= add_ln703_226_fu_1457_p2;
        add_ln703_227_reg_10752 <= add_ln703_227_fu_1472_p2;
        add_ln703_233_reg_10767 <= add_ln703_233_fu_1501_p2;
        add_ln703_236_reg_10772 <= add_ln703_236_fu_1511_p2;
        add_ln703_238_reg_10777 <= add_ln703_238_fu_1520_p2;
        add_ln703_247_reg_10802 <= add_ln703_247_fu_1563_p2;
        add_ln703_250_reg_10807 <= add_ln703_250_fu_1574_p2;
        add_ln703_252_reg_10665 <= add_ln703_252_fu_1077_p2;
        add_ln703_252_reg_10665_pp0_iter5_reg <= add_ln703_252_reg_10665;
        add_ln703_254_reg_10672 <= add_ln703_254_fu_1081_p2;
        add_ln703_260_reg_10817 <= add_ln703_260_fu_1593_p2;
        add_ln703_262_reg_10827 <= add_ln703_262_fu_1604_p2;
        add_ln703_265_reg_10837 <= add_ln703_265_fu_1614_p2;
        add_ln703_280_reg_10846 <= add_ln703_280_fu_1618_p2;
        add_ln703_283_reg_10873 <= add_ln703_283_fu_1979_p2;
        add_ln703_285_reg_10888 <= add_ln703_285_fu_2009_p2;
        add_ln703_289_reg_10898 <= add_ln703_289_fu_2034_p2;
        add_ln703_290_reg_10903 <= add_ln703_290_fu_2039_p2;
        add_ln703_294_reg_10918 <= add_ln703_294_fu_2084_p2;
        add_ln703_295_reg_10923 <= add_ln703_295_fu_2089_p2;
        add_ln703_300_reg_10930 <= add_ln703_300_fu_2093_p2;
        add_ln703_303_reg_10940 <= add_ln703_303_fu_2104_p2;
        add_ln703_304_reg_10945 <= add_ln703_304_fu_2110_p2;
        add_ln703_307_reg_10960 <= add_ln703_307_fu_2125_p2;
        add_ln703_309_reg_10970 <= add_ln703_309_fu_2136_p2;
        add_ln703_310_reg_10980 <= add_ln703_310_fu_2147_p2;
        add_ln703_323_reg_11005 <= add_ln703_323_fu_2188_p2;
        add_ln703_326_reg_10855 <= add_ln703_326_fu_1622_p2;
        add_ln703_326_reg_10855_pp0_iter6_reg <= add_ln703_326_reg_10855;
        add_ln703_328_reg_11015 <= add_ln703_328_fu_2208_p2;
        add_ln703_333_reg_11025 <= add_ln703_333_fu_2224_p2;
        add_ln703_341_reg_11030 <= add_ln703_341_fu_2230_p2;
        add_ln703_342_reg_11071 <= add_ln703_342_fu_2520_p2;
        add_ln703_346_reg_11106 <= add_ln703_346_fu_2589_p2;
        add_ln703_350_reg_11111 <= add_ln703_350_fu_2602_p2;
        add_ln703_352_reg_11126 <= add_ln703_352_fu_2633_p2;
        add_ln703_354_reg_11131 <= add_ln703_354_fu_2638_p2;
        add_ln703_356_reg_11148 <= add_ln703_356_fu_2657_p2;
        add_ln703_360_reg_11158 <= add_ln703_360_fu_2677_p2;
        add_ln703_369_reg_11037 <= add_ln703_369_fu_2234_p2;
        add_ln703_369_reg_11037_pp0_iter7_reg <= add_ln703_369_reg_11037;
        add_ln703_371_reg_11193 <= add_ln703_371_fu_2732_p2;
        add_ln703_375_reg_11198 <= add_ln703_375_fu_2738_p2;
        add_ln703_384_reg_11203 <= add_ln703_384_fu_2743_p2;
        add_ln703_386_reg_11262 <= add_ln703_386_fu_3015_p2;
        add_ln703_390_reg_11272 <= add_ln703_390_fu_3050_p2;
        add_ln703_400_reg_11210 <= add_ln703_400_fu_2752_p2;
        add_ln703_402_reg_11215 <= add_ln703_402_fu_2758_p2;
        add_ln703_402_reg_11215_pp0_iter8_reg <= add_ln703_402_reg_11215;
        add_ln703_410_reg_11287 <= add_ln703_410_fu_3149_p2;
        add_ln703_416_reg_11297 <= add_ln703_416_fu_3170_p2;
        add_ln703_417_reg_11312 <= add_ln703_417_fu_3185_p2;
        add_ln703_424_reg_11225 <= add_ln703_424_fu_2762_p2;
        add_ln703_426_reg_11347 <= add_ln703_426_fu_3258_p2;
        add_ln703_431_reg_11357 <= add_ln703_431_fu_3274_p2;
        add_ln703_435_reg_11362 <= add_ln703_435_fu_3284_p2;
        add_ln703_438_reg_11382 <= add_ln703_438_fu_3310_p2;
        add_ln703_439_reg_11233 <= add_ln703_439_fu_2766_p2;
        add_ln703_439_reg_11233_pp0_iter8_reg <= add_ln703_439_reg_11233;
        add_ln703_445_reg_11387 <= add_ln703_445_fu_3315_p2;
        add_ln703_447_reg_11392 <= add_ln703_447_fu_3320_p2;
        add_ln703_451_reg_11402 <= add_ln703_451_fu_3329_p2;
        add_ln703_466_reg_11410 <= add_ln703_466_fu_3333_p2;
        add_ln703_469_reg_11479 <= add_ln703_469_fu_3655_p2;
        add_ln703_471_reg_11418 <= add_ln703_471_fu_3337_p2;
        add_ln703_476_reg_11494 <= add_ln703_476_fu_3685_p2;
        add_ln703_478_reg_11519 <= add_ln703_478_fu_3730_p2;
        add_ln703_484_reg_11423 <= add_ln703_484_fu_3342_p2;
        add_ln703_490_reg_11428 <= add_ln703_490_fu_3347_p2;
        add_ln703_496_reg_11544 <= add_ln703_496_fu_3806_p2;
        add_ln703_497_reg_11549 <= add_ln703_497_fu_3811_p2;
        add_ln703_498_reg_11436 <= add_ln703_498_fu_3351_p2;
        add_ln703_506_reg_11559 <= add_ln703_506_fu_3839_p2;
        add_ln703_507_reg_11441 <= add_ln703_507_fu_3356_p2;
        add_ln703_507_reg_11441_pp0_iter9_reg <= add_ln703_507_reg_11441;
        add_ln703_512_reg_11589 <= add_ln703_512_fu_3878_p2;
        add_ln703_515_reg_11599 <= add_ln703_515_fu_3889_p2;
        add_ln703_517_reg_11604 <= add_ln703_517_fu_3894_p2;
        add_ln703_525_reg_11243 <= add_ln703_525_fu_2774_p2;
        add_ln703_525_reg_11243_pp0_iter8_reg <= add_ln703_525_reg_11243;
        add_ln703_525_reg_11243_pp0_iter9_reg <= add_ln703_525_reg_11243_pp0_iter8_reg;
        add_ln703_528_reg_11452 <= add_ln703_528_fu_3360_p2;
        add_ln703_528_reg_11452_pp0_iter9_reg <= add_ln703_528_reg_11452;
        add_ln703_534_reg_11248 <= add_ln703_534_fu_2779_p2;
        add_ln703_534_reg_11248_pp0_iter8_reg <= add_ln703_534_reg_11248;
        add_ln703_534_reg_11248_pp0_iter9_reg <= add_ln703_534_reg_11248_pp0_iter8_reg;
        add_ln703_535_reg_11457 <= add_ln703_535_fu_3364_p2;
        add_ln703_537_reg_11609 <= add_ln703_537_fu_3912_p2;
        add_ln703_545_reg_11614 <= add_ln703_545_fu_3923_p2;
        add_ln703_556_reg_11619 <= add_ln703_556_fu_3933_p2;
        add_ln703_560_reg_11629 <= add_ln703_560_fu_3943_p2;
        add_ln703_566_reg_11635 <= add_ln703_566_fu_3952_p2;
        add_ln703_568_reg_11464 <= add_ln703_568_fu_3368_p2;
        add_ln703_568_reg_11464_pp0_iter9_reg <= add_ln703_568_reg_11464;
        add_ln703_569_reg_11640 <= add_ln703_569_fu_3957_p2;
        add_ln703_572_reg_11698 <= add_ln703_572_fu_4308_p2;
        add_ln703_573_reg_11708 <= add_ln703_573_fu_4323_p2;
        add_ln703_581_reg_11723 <= add_ln703_581_fu_4358_p2;
        add_ln703_583_reg_11728 <= add_ln703_583_fu_4363_p2;
        add_ln703_586_reg_11743 <= add_ln703_586_fu_4398_p2;
        add_ln703_588_reg_11646 <= add_ln703_588_fu_3961_p2;
        add_ln703_590_reg_11748 <= add_ln703_590_fu_4412_p2;
        add_ln703_591_reg_11758 <= add_ln703_591_fu_4423_p2;
        add_ln703_592_reg_11763 <= add_ln703_592_fu_4428_p2;
        add_ln703_598_reg_11768 <= add_ln703_598_fu_4441_p2;
        add_ln703_599_reg_11798 <= add_ln703_599_fu_4477_p2;
        add_ln703_600_reg_11652 <= add_ln703_600_fu_3965_p2;
        add_ln703_600_reg_11652_pp0_iter10_reg <= add_ln703_600_reg_11652;
        add_ln703_609_reg_11803 <= add_ln703_609_fu_4501_p2;
        add_ln703_616_reg_11808 <= add_ln703_616_fu_4511_p2;
        add_ln703_621_reg_11662 <= add_ln703_621_fu_3969_p2;
        add_ln703_621_reg_11662_pp0_iter10_reg <= add_ln703_621_reg_11662;
        add_ln703_633_reg_11823 <= add_ln703_633_fu_4531_p2;
        add_ln703_634_reg_11828 <= add_ln703_634_fu_4535_p2;
        add_ln703_639_reg_11833 <= add_ln703_639_fu_4541_p2;
        add_ln703_646_reg_11838 <= add_ln703_646_fu_4546_p2;
        add_ln703_647_reg_11874 <= add_ln703_647_fu_4870_p2;
        add_ln703_648_reg_11889 <= add_ln703_648_fu_4899_p2;
        add_ln703_650_reg_11844 <= add_ln703_650_fu_4550_p2;
        add_ln703_650_reg_11844_pp0_iter11_reg <= add_ln703_650_reg_11844;
        add_ln703_651_reg_11929 <= add_ln703_651_fu_4959_p2;
        add_ln703_660_reg_11939 <= add_ln703_660_fu_4994_p2;
        add_ln703_661_reg_11944 <= add_ln703_661_fu_4999_p2;
        add_ln703_666_reg_11954 <= add_ln703_666_fu_5013_p2;
        add_ln703_667_reg_11853 <= add_ln703_667_fu_4554_p2;
        add_ln703_668_reg_11959 <= add_ln703_668_fu_5019_p2;
        add_ln703_676_reg_11979 <= add_ln703_676_fu_5052_p2;
        add_ln703_682_reg_11984 <= add_ln703_682_fu_5066_p2;
        add_ln703_685_reg_11989 <= add_ln703_685_fu_5077_p2;
        add_ln703_691_reg_11994 <= add_ln703_691_fu_5092_p2;
        add_ln703_697_reg_12002 <= add_ln703_697_fu_5096_p2;
        add_ln703_703_reg_12022 <= add_ln703_703_fu_5116_p2;
        add_ln703_704_reg_12056 <= add_ln703_704_fu_5336_p2;
        add_ln703_706_reg_12031 <= add_ln703_706_fu_5120_p2;
        add_ln703_719_reg_12086 <= add_ln703_719_fu_5439_p2;
        add_ln703_722_reg_12036 <= add_ln703_722_fu_5125_p2;
        add_ln703_726_reg_12041 <= add_ln703_726_fu_5130_p2;
        add_ln703_728_reg_12096 <= add_ln703_728_fu_5485_p2;
        add_ln703_733_reg_12146 <= add_ln703_733_fu_5551_p2;
        add_ln703_734_reg_12151 <= add_ln703_734_fu_5556_p2;
        add_ln703_735_reg_12161 <= add_ln703_735_fu_5571_p2;
        add_ln703_737_reg_12047 <= add_ln703_737_fu_5134_p2;
        add_ln703_755_reg_12196 <= add_ln703_755_fu_5652_p2;
        add_ln703_765_reg_12219 <= add_ln703_765_fu_5671_p2;
        add_ln703_770_reg_12258 <= add_ln703_770_fu_5950_p2;
        add_ln703_778_reg_12227 <= add_ln703_778_fu_5675_p2;
        add_ln703_779_reg_12273 <= add_ln703_779_fu_6024_p2;
        add_ln703_783_reg_12236 <= add_ln703_783_fu_5679_p2;
        add_ln703_791_reg_12348 <= add_ln703_791_fu_6131_p2;
        add_ln703_792_reg_12363 <= add_ln703_792_fu_6146_p2;
        add_ln703_796_reg_12368 <= add_ln703_796_fu_6160_p2;
        add_ln703_798_reg_12373 <= add_ln703_798_fu_6166_p2;
        add_ln703_801_reg_12393 <= add_ln703_801_fu_6187_p2;
        add_ln703_802_reg_12398 <= add_ln703_802_fu_6192_p2;
        add_ln703_816_reg_12241 <= add_ln703_816_fu_5684_p2;
        add_ln703_816_reg_12241_pp0_iter13_reg <= add_ln703_816_reg_12241;
        add_ln703_818_reg_12409 <= add_ln703_818_fu_6205_p2;
        add_ln703_818_reg_12409_pp0_iter14_reg <= add_ln703_818_reg_12409;
        add_ln703_819_reg_12455 <= add_ln703_819_fu_6447_p2;
        add_ln703_821_reg_12414 <= add_ln703_821_fu_6216_p2;
        add_ln703_825_reg_12480 <= add_ln703_825_fu_6526_p2;
        add_ln703_826_reg_12419 <= add_ln703_826_fu_6222_p2;
        add_ln703_827_reg_12485 <= add_ln703_827_fu_6531_p2;
        add_ln703_831_reg_12490 <= add_ln703_831_fu_6554_p2;
        add_ln703_833_reg_12495 <= add_ln703_833_fu_6573_p2;
        add_ln703_834_reg_12505 <= add_ln703_834_fu_6594_p2;
        add_ln703_836_reg_12428 <= add_ln703_836_fu_6226_p2;
        add_ln703_838_reg_12520 <= add_ln703_838_fu_6634_p2;
        add_ln703_840_reg_12535 <= add_ln703_840_fu_6649_p2;
        add_ln703_841_reg_12550 <= add_ln703_841_fu_6664_p2;
        add_ln703_845_reg_12560 <= add_ln703_845_fu_6689_p2;
        add_ln703_849_reg_12434 <= add_ln703_849_fu_6230_p2;
        add_ln703_849_reg_12434_pp0_iter14_reg <= add_ln703_849_reg_12434;
        add_ln703_851_reg_12565 <= add_ln703_851_fu_6702_p2;
        add_ln703_858_reg_12575 <= add_ln703_858_fu_6733_p2;
        add_ln703_867_reg_12444 <= add_ln703_867_fu_6234_p2;
        add_ln703_867_reg_12444_pp0_iter14_reg <= add_ln703_867_reg_12444;
        add_ln703_868_reg_12585 <= add_ln703_868_fu_6755_p2;
        add_ln703_872_reg_12650 <= add_ln703_872_fu_7050_p2;
        add_ln703_873_reg_12655 <= add_ln703_873_fu_7055_p2;
        add_ln703_874_reg_12675 <= add_ln703_874_fu_7084_p2;
        add_ln703_875_reg_12680 <= add_ln703_875_fu_7094_p2;
        add_ln703_876_reg_12600 <= add_ln703_876_fu_6769_p2;
        add_ln703_877_reg_12605 <= add_ln703_877_fu_6774_p2;
        add_ln703_882_reg_12690 <= add_ln703_882_fu_7121_p2;
        add_ln703_884_reg_12695 <= add_ln703_884_fu_7132_p2;
        add_ln703_888_reg_12705 <= add_ln703_888_fu_7156_p2;
        add_ln703_892_reg_12710 <= add_ln703_892_fu_7175_p2;
        add_ln703_893_reg_12715 <= add_ln703_893_fu_7180_p2;
        add_ln703_894_reg_12616 <= add_ln703_894_fu_6778_p2;
        add_ln703_894_reg_12616_pp0_iter15_reg <= add_ln703_894_reg_12616;
        add_ln703_895_reg_12720 <= add_ln703_895_fu_7185_p2;
        add_ln703_896_reg_12725 <= add_ln703_896_fu_7190_p2;
        add_ln703_898_reg_12730 <= add_ln703_898_fu_7195_p2;
        add_ln703_905_reg_12625 <= add_ln703_905_fu_6782_p2;
        add_ln703_906_reg_12775 <= add_ln703_906_fu_7245_p2;
        add_ln703_914_reg_12632 <= add_ln703_914_fu_6786_p2;
        add_ln703_917_reg_12780 <= add_ln703_917_fu_7273_p2;
        add_ln703_920_reg_12637 <= add_ln703_920_fu_6791_p2;
        add_ln703_920_reg_12637_pp0_iter15_reg <= add_ln703_920_reg_12637;
        add_ln703_922_reg_12785 <= add_ln703_922_fu_7287_p2;
        add_ln703_934_reg_12845 <= add_ln703_934_fu_7610_p2;
        add_ln703_936_reg_12855 <= add_ln703_936_fu_7634_p2;
        add_ln703_938_reg_12875 <= add_ln703_938_fu_7663_p2;
        add_ln703_939_reg_12890 <= add_ln703_939_fu_7679_p2;
        add_ln703_943_reg_12905 <= add_ln703_943_fu_7719_p2;
        add_ln703_946_reg_12805 <= add_ln703_946_fu_7334_p2;
        add_ln703_948_reg_12930 <= add_ln703_948_fu_7760_p2;
        add_ln703_954_reg_12812 <= add_ln703_954_fu_7338_p2;
        add_ln703_958_reg_12965 <= add_ln703_958_fu_7827_p2;
        add_ln703_964_reg_12985 <= add_ln703_964_fu_7848_p2;
        add_ln703_985_reg_12819 <= add_ln703_985_fu_7342_p2;
        add_ln703_985_reg_12819_pp0_iter16_reg <= add_ln703_985_reg_12819;
        add_ln703_reg_10335 <= add_ln703_fu_530_p2;
        add_ln703_reg_10335_pp0_iter1_reg <= add_ln703_reg_10335;
        data_0_V_read_10_reg_10329 <= data_0_V_read_int_reg;
        data_10_V_read11_reg_10105 <= data_10_V_read_int_reg;
        data_10_V_read11_reg_10105_pp0_iter1_reg <= data_10_V_read11_reg_10105;
        data_10_V_read11_reg_10105_pp0_iter2_reg <= data_10_V_read11_reg_10105_pp0_iter1_reg;
        data_10_V_read11_reg_10105_pp0_iter3_reg <= data_10_V_read11_reg_10105_pp0_iter2_reg;
        data_10_V_read11_reg_10105_pp0_iter4_reg <= data_10_V_read11_reg_10105_pp0_iter3_reg;
        data_11_V_read12_reg_10075 <= data_11_V_read_int_reg;
        data_11_V_read12_reg_10075_pp0_iter1_reg <= data_11_V_read12_reg_10075;
        data_11_V_read12_reg_10075_pp0_iter2_reg <= data_11_V_read12_reg_10075_pp0_iter1_reg;
        data_11_V_read12_reg_10075_pp0_iter3_reg <= data_11_V_read12_reg_10075_pp0_iter2_reg;
        data_11_V_read12_reg_10075_pp0_iter4_reg <= data_11_V_read12_reg_10075_pp0_iter3_reg;
        data_11_V_read12_reg_10075_pp0_iter5_reg <= data_11_V_read12_reg_10075_pp0_iter4_reg;
        data_12_V_read13_reg_10045 <= data_12_V_read_int_reg;
        data_12_V_read13_reg_10045_pp0_iter1_reg <= data_12_V_read13_reg_10045;
        data_12_V_read13_reg_10045_pp0_iter2_reg <= data_12_V_read13_reg_10045_pp0_iter1_reg;
        data_12_V_read13_reg_10045_pp0_iter3_reg <= data_12_V_read13_reg_10045_pp0_iter2_reg;
        data_12_V_read13_reg_10045_pp0_iter4_reg <= data_12_V_read13_reg_10045_pp0_iter3_reg;
        data_12_V_read13_reg_10045_pp0_iter5_reg <= data_12_V_read13_reg_10045_pp0_iter4_reg;
        data_13_V_read14_reg_10015 <= data_13_V_read_int_reg;
        data_13_V_read14_reg_10015_pp0_iter1_reg <= data_13_V_read14_reg_10015;
        data_13_V_read14_reg_10015_pp0_iter2_reg <= data_13_V_read14_reg_10015_pp0_iter1_reg;
        data_13_V_read14_reg_10015_pp0_iter3_reg <= data_13_V_read14_reg_10015_pp0_iter2_reg;
        data_13_V_read14_reg_10015_pp0_iter4_reg <= data_13_V_read14_reg_10015_pp0_iter3_reg;
        data_13_V_read14_reg_10015_pp0_iter5_reg <= data_13_V_read14_reg_10015_pp0_iter4_reg;
        data_14_V_read15_reg_9987 <= data_14_V_read_int_reg;
        data_14_V_read15_reg_9987_pp0_iter1_reg <= data_14_V_read15_reg_9987;
        data_14_V_read15_reg_9987_pp0_iter2_reg <= data_14_V_read15_reg_9987_pp0_iter1_reg;
        data_14_V_read15_reg_9987_pp0_iter3_reg <= data_14_V_read15_reg_9987_pp0_iter2_reg;
        data_14_V_read15_reg_9987_pp0_iter4_reg <= data_14_V_read15_reg_9987_pp0_iter3_reg;
        data_14_V_read15_reg_9987_pp0_iter5_reg <= data_14_V_read15_reg_9987_pp0_iter4_reg;
        data_15_V_read16_reg_9962 <= data_15_V_read_int_reg;
        data_15_V_read16_reg_9962_pp0_iter1_reg <= data_15_V_read16_reg_9962;
        data_15_V_read16_reg_9962_pp0_iter2_reg <= data_15_V_read16_reg_9962_pp0_iter1_reg;
        data_15_V_read16_reg_9962_pp0_iter3_reg <= data_15_V_read16_reg_9962_pp0_iter2_reg;
        data_15_V_read16_reg_9962_pp0_iter4_reg <= data_15_V_read16_reg_9962_pp0_iter3_reg;
        data_15_V_read16_reg_9962_pp0_iter5_reg <= data_15_V_read16_reg_9962_pp0_iter4_reg;
        data_16_V_read17_reg_9935 <= data_16_V_read_int_reg;
        data_16_V_read17_reg_9935_pp0_iter1_reg <= data_16_V_read17_reg_9935;
        data_16_V_read17_reg_9935_pp0_iter2_reg <= data_16_V_read17_reg_9935_pp0_iter1_reg;
        data_16_V_read17_reg_9935_pp0_iter3_reg <= data_16_V_read17_reg_9935_pp0_iter2_reg;
        data_16_V_read17_reg_9935_pp0_iter4_reg <= data_16_V_read17_reg_9935_pp0_iter3_reg;
        data_16_V_read17_reg_9935_pp0_iter5_reg <= data_16_V_read17_reg_9935_pp0_iter4_reg;
        data_16_V_read17_reg_9935_pp0_iter6_reg <= data_16_V_read17_reg_9935_pp0_iter5_reg;
        data_17_V_read18_reg_9904 <= data_17_V_read_int_reg;
        data_17_V_read18_reg_9904_pp0_iter1_reg <= data_17_V_read18_reg_9904;
        data_17_V_read18_reg_9904_pp0_iter2_reg <= data_17_V_read18_reg_9904_pp0_iter1_reg;
        data_17_V_read18_reg_9904_pp0_iter3_reg <= data_17_V_read18_reg_9904_pp0_iter2_reg;
        data_17_V_read18_reg_9904_pp0_iter4_reg <= data_17_V_read18_reg_9904_pp0_iter3_reg;
        data_17_V_read18_reg_9904_pp0_iter5_reg <= data_17_V_read18_reg_9904_pp0_iter4_reg;
        data_17_V_read18_reg_9904_pp0_iter6_reg <= data_17_V_read18_reg_9904_pp0_iter5_reg;
        data_18_V_read_8_reg_9874 <= data_18_V_read_int_reg;
        data_18_V_read_8_reg_9874_pp0_iter1_reg <= data_18_V_read_8_reg_9874;
        data_18_V_read_8_reg_9874_pp0_iter2_reg <= data_18_V_read_8_reg_9874_pp0_iter1_reg;
        data_18_V_read_8_reg_9874_pp0_iter3_reg <= data_18_V_read_8_reg_9874_pp0_iter2_reg;
        data_18_V_read_8_reg_9874_pp0_iter4_reg <= data_18_V_read_8_reg_9874_pp0_iter3_reg;
        data_18_V_read_8_reg_9874_pp0_iter5_reg <= data_18_V_read_8_reg_9874_pp0_iter4_reg;
        data_18_V_read_8_reg_9874_pp0_iter6_reg <= data_18_V_read_8_reg_9874_pp0_iter5_reg;
        data_19_V_read_8_reg_9845 <= data_19_V_read_int_reg;
        data_19_V_read_8_reg_9845_pp0_iter1_reg <= data_19_V_read_8_reg_9845;
        data_19_V_read_8_reg_9845_pp0_iter2_reg <= data_19_V_read_8_reg_9845_pp0_iter1_reg;
        data_19_V_read_8_reg_9845_pp0_iter3_reg <= data_19_V_read_8_reg_9845_pp0_iter2_reg;
        data_19_V_read_8_reg_9845_pp0_iter4_reg <= data_19_V_read_8_reg_9845_pp0_iter3_reg;
        data_19_V_read_8_reg_9845_pp0_iter5_reg <= data_19_V_read_8_reg_9845_pp0_iter4_reg;
        data_19_V_read_8_reg_9845_pp0_iter6_reg <= data_19_V_read_8_reg_9845_pp0_iter5_reg;
        data_1_V_read_10_reg_10323 <= data_1_V_read_int_reg;
        data_20_V_read21_reg_9814 <= data_20_V_read_int_reg;
        data_20_V_read21_reg_9814_pp0_iter1_reg <= data_20_V_read21_reg_9814;
        data_20_V_read21_reg_9814_pp0_iter2_reg <= data_20_V_read21_reg_9814_pp0_iter1_reg;
        data_20_V_read21_reg_9814_pp0_iter3_reg <= data_20_V_read21_reg_9814_pp0_iter2_reg;
        data_20_V_read21_reg_9814_pp0_iter4_reg <= data_20_V_read21_reg_9814_pp0_iter3_reg;
        data_20_V_read21_reg_9814_pp0_iter5_reg <= data_20_V_read21_reg_9814_pp0_iter4_reg;
        data_20_V_read21_reg_9814_pp0_iter6_reg <= data_20_V_read21_reg_9814_pp0_iter5_reg;
        data_20_V_read21_reg_9814_pp0_iter7_reg <= data_20_V_read21_reg_9814_pp0_iter6_reg;
        data_21_V_read22_reg_9784 <= data_21_V_read_int_reg;
        data_21_V_read22_reg_9784_pp0_iter1_reg <= data_21_V_read22_reg_9784;
        data_21_V_read22_reg_9784_pp0_iter2_reg <= data_21_V_read22_reg_9784_pp0_iter1_reg;
        data_21_V_read22_reg_9784_pp0_iter3_reg <= data_21_V_read22_reg_9784_pp0_iter2_reg;
        data_21_V_read22_reg_9784_pp0_iter4_reg <= data_21_V_read22_reg_9784_pp0_iter3_reg;
        data_21_V_read22_reg_9784_pp0_iter5_reg <= data_21_V_read22_reg_9784_pp0_iter4_reg;
        data_21_V_read22_reg_9784_pp0_iter6_reg <= data_21_V_read22_reg_9784_pp0_iter5_reg;
        data_21_V_read22_reg_9784_pp0_iter7_reg <= data_21_V_read22_reg_9784_pp0_iter6_reg;
        data_22_V_read23_reg_9756 <= data_22_V_read_int_reg;
        data_22_V_read23_reg_9756_pp0_iter1_reg <= data_22_V_read23_reg_9756;
        data_22_V_read23_reg_9756_pp0_iter2_reg <= data_22_V_read23_reg_9756_pp0_iter1_reg;
        data_22_V_read23_reg_9756_pp0_iter3_reg <= data_22_V_read23_reg_9756_pp0_iter2_reg;
        data_22_V_read23_reg_9756_pp0_iter4_reg <= data_22_V_read23_reg_9756_pp0_iter3_reg;
        data_22_V_read23_reg_9756_pp0_iter5_reg <= data_22_V_read23_reg_9756_pp0_iter4_reg;
        data_22_V_read23_reg_9756_pp0_iter6_reg <= data_22_V_read23_reg_9756_pp0_iter5_reg;
        data_22_V_read23_reg_9756_pp0_iter7_reg <= data_22_V_read23_reg_9756_pp0_iter6_reg;
        data_22_V_read23_reg_9756_pp0_iter8_reg <= data_22_V_read23_reg_9756_pp0_iter7_reg;
        data_23_V_read24_reg_9730 <= data_23_V_read_int_reg;
        data_23_V_read24_reg_9730_pp0_iter1_reg <= data_23_V_read24_reg_9730;
        data_23_V_read24_reg_9730_pp0_iter2_reg <= data_23_V_read24_reg_9730_pp0_iter1_reg;
        data_23_V_read24_reg_9730_pp0_iter3_reg <= data_23_V_read24_reg_9730_pp0_iter2_reg;
        data_23_V_read24_reg_9730_pp0_iter4_reg <= data_23_V_read24_reg_9730_pp0_iter3_reg;
        data_23_V_read24_reg_9730_pp0_iter5_reg <= data_23_V_read24_reg_9730_pp0_iter4_reg;
        data_23_V_read24_reg_9730_pp0_iter6_reg <= data_23_V_read24_reg_9730_pp0_iter5_reg;
        data_23_V_read24_reg_9730_pp0_iter7_reg <= data_23_V_read24_reg_9730_pp0_iter6_reg;
        data_24_V_read25_reg_9704 <= data_24_V_read_int_reg;
        data_24_V_read25_reg_9704_pp0_iter1_reg <= data_24_V_read25_reg_9704;
        data_24_V_read25_reg_9704_pp0_iter2_reg <= data_24_V_read25_reg_9704_pp0_iter1_reg;
        data_24_V_read25_reg_9704_pp0_iter3_reg <= data_24_V_read25_reg_9704_pp0_iter2_reg;
        data_24_V_read25_reg_9704_pp0_iter4_reg <= data_24_V_read25_reg_9704_pp0_iter3_reg;
        data_24_V_read25_reg_9704_pp0_iter5_reg <= data_24_V_read25_reg_9704_pp0_iter4_reg;
        data_24_V_read25_reg_9704_pp0_iter6_reg <= data_24_V_read25_reg_9704_pp0_iter5_reg;
        data_24_V_read25_reg_9704_pp0_iter7_reg <= data_24_V_read25_reg_9704_pp0_iter6_reg;
        data_24_V_read25_reg_9704_pp0_iter8_reg <= data_24_V_read25_reg_9704_pp0_iter7_reg;
        data_25_V_read26_reg_9677 <= data_25_V_read_int_reg;
        data_25_V_read26_reg_9677_pp0_iter1_reg <= data_25_V_read26_reg_9677;
        data_25_V_read26_reg_9677_pp0_iter2_reg <= data_25_V_read26_reg_9677_pp0_iter1_reg;
        data_25_V_read26_reg_9677_pp0_iter3_reg <= data_25_V_read26_reg_9677_pp0_iter2_reg;
        data_25_V_read26_reg_9677_pp0_iter4_reg <= data_25_V_read26_reg_9677_pp0_iter3_reg;
        data_25_V_read26_reg_9677_pp0_iter5_reg <= data_25_V_read26_reg_9677_pp0_iter4_reg;
        data_25_V_read26_reg_9677_pp0_iter6_reg <= data_25_V_read26_reg_9677_pp0_iter5_reg;
        data_25_V_read26_reg_9677_pp0_iter7_reg <= data_25_V_read26_reg_9677_pp0_iter6_reg;
        data_25_V_read26_reg_9677_pp0_iter8_reg <= data_25_V_read26_reg_9677_pp0_iter7_reg;
        data_26_V_read27_reg_9652 <= data_26_V_read_int_reg;
        data_26_V_read27_reg_9652_pp0_iter1_reg <= data_26_V_read27_reg_9652;
        data_26_V_read27_reg_9652_pp0_iter2_reg <= data_26_V_read27_reg_9652_pp0_iter1_reg;
        data_26_V_read27_reg_9652_pp0_iter3_reg <= data_26_V_read27_reg_9652_pp0_iter2_reg;
        data_26_V_read27_reg_9652_pp0_iter4_reg <= data_26_V_read27_reg_9652_pp0_iter3_reg;
        data_26_V_read27_reg_9652_pp0_iter5_reg <= data_26_V_read27_reg_9652_pp0_iter4_reg;
        data_26_V_read27_reg_9652_pp0_iter6_reg <= data_26_V_read27_reg_9652_pp0_iter5_reg;
        data_26_V_read27_reg_9652_pp0_iter7_reg <= data_26_V_read27_reg_9652_pp0_iter6_reg;
        data_26_V_read27_reg_9652_pp0_iter8_reg <= data_26_V_read27_reg_9652_pp0_iter7_reg;
        data_27_V_read28_reg_9625 <= data_27_V_read_int_reg;
        data_27_V_read28_reg_9625_pp0_iter1_reg <= data_27_V_read28_reg_9625;
        data_27_V_read28_reg_9625_pp0_iter2_reg <= data_27_V_read28_reg_9625_pp0_iter1_reg;
        data_27_V_read28_reg_9625_pp0_iter3_reg <= data_27_V_read28_reg_9625_pp0_iter2_reg;
        data_27_V_read28_reg_9625_pp0_iter4_reg <= data_27_V_read28_reg_9625_pp0_iter3_reg;
        data_27_V_read28_reg_9625_pp0_iter5_reg <= data_27_V_read28_reg_9625_pp0_iter4_reg;
        data_27_V_read28_reg_9625_pp0_iter6_reg <= data_27_V_read28_reg_9625_pp0_iter5_reg;
        data_27_V_read28_reg_9625_pp0_iter7_reg <= data_27_V_read28_reg_9625_pp0_iter6_reg;
        data_27_V_read28_reg_9625_pp0_iter8_reg <= data_27_V_read28_reg_9625_pp0_iter7_reg;
        data_28_V_read_8_reg_9598 <= data_28_V_read_int_reg;
        data_28_V_read_8_reg_9598_pp0_iter1_reg <= data_28_V_read_8_reg_9598;
        data_28_V_read_8_reg_9598_pp0_iter2_reg <= data_28_V_read_8_reg_9598_pp0_iter1_reg;
        data_28_V_read_8_reg_9598_pp0_iter3_reg <= data_28_V_read_8_reg_9598_pp0_iter2_reg;
        data_28_V_read_8_reg_9598_pp0_iter4_reg <= data_28_V_read_8_reg_9598_pp0_iter3_reg;
        data_28_V_read_8_reg_9598_pp0_iter5_reg <= data_28_V_read_8_reg_9598_pp0_iter4_reg;
        data_28_V_read_8_reg_9598_pp0_iter6_reg <= data_28_V_read_8_reg_9598_pp0_iter5_reg;
        data_28_V_read_8_reg_9598_pp0_iter7_reg <= data_28_V_read_8_reg_9598_pp0_iter6_reg;
        data_28_V_read_8_reg_9598_pp0_iter8_reg <= data_28_V_read_8_reg_9598_pp0_iter7_reg;
        data_29_V_read_8_reg_9573 <= data_29_V_read_int_reg;
        data_29_V_read_8_reg_9573_pp0_iter1_reg <= data_29_V_read_8_reg_9573;
        data_29_V_read_8_reg_9573_pp0_iter2_reg <= data_29_V_read_8_reg_9573_pp0_iter1_reg;
        data_29_V_read_8_reg_9573_pp0_iter3_reg <= data_29_V_read_8_reg_9573_pp0_iter2_reg;
        data_29_V_read_8_reg_9573_pp0_iter4_reg <= data_29_V_read_8_reg_9573_pp0_iter3_reg;
        data_29_V_read_8_reg_9573_pp0_iter5_reg <= data_29_V_read_8_reg_9573_pp0_iter4_reg;
        data_29_V_read_8_reg_9573_pp0_iter6_reg <= data_29_V_read_8_reg_9573_pp0_iter5_reg;
        data_29_V_read_8_reg_9573_pp0_iter7_reg <= data_29_V_read_8_reg_9573_pp0_iter6_reg;
        data_29_V_read_8_reg_9573_pp0_iter8_reg <= data_29_V_read_8_reg_9573_pp0_iter7_reg;
        data_29_V_read_8_reg_9573_pp0_iter9_reg <= data_29_V_read_8_reg_9573_pp0_iter8_reg;
        data_2_V_read_10_reg_10312 <= data_2_V_read_int_reg;
        data_2_V_read_10_reg_10312_pp0_iter1_reg <= data_2_V_read_10_reg_10312;
        data_30_V_read31_reg_9549 <= data_30_V_read_int_reg;
        data_30_V_read31_reg_9549_pp0_iter1_reg <= data_30_V_read31_reg_9549;
        data_30_V_read31_reg_9549_pp0_iter2_reg <= data_30_V_read31_reg_9549_pp0_iter1_reg;
        data_30_V_read31_reg_9549_pp0_iter3_reg <= data_30_V_read31_reg_9549_pp0_iter2_reg;
        data_30_V_read31_reg_9549_pp0_iter4_reg <= data_30_V_read31_reg_9549_pp0_iter3_reg;
        data_30_V_read31_reg_9549_pp0_iter5_reg <= data_30_V_read31_reg_9549_pp0_iter4_reg;
        data_30_V_read31_reg_9549_pp0_iter6_reg <= data_30_V_read31_reg_9549_pp0_iter5_reg;
        data_30_V_read31_reg_9549_pp0_iter7_reg <= data_30_V_read31_reg_9549_pp0_iter6_reg;
        data_30_V_read31_reg_9549_pp0_iter8_reg <= data_30_V_read31_reg_9549_pp0_iter7_reg;
        data_30_V_read31_reg_9549_pp0_iter9_reg <= data_30_V_read31_reg_9549_pp0_iter8_reg;
        data_31_V_read32_reg_9521 <= data_31_V_read_int_reg;
        data_31_V_read32_reg_9521_pp0_iter1_reg <= data_31_V_read32_reg_9521;
        data_31_V_read32_reg_9521_pp0_iter2_reg <= data_31_V_read32_reg_9521_pp0_iter1_reg;
        data_31_V_read32_reg_9521_pp0_iter3_reg <= data_31_V_read32_reg_9521_pp0_iter2_reg;
        data_31_V_read32_reg_9521_pp0_iter4_reg <= data_31_V_read32_reg_9521_pp0_iter3_reg;
        data_31_V_read32_reg_9521_pp0_iter5_reg <= data_31_V_read32_reg_9521_pp0_iter4_reg;
        data_31_V_read32_reg_9521_pp0_iter6_reg <= data_31_V_read32_reg_9521_pp0_iter5_reg;
        data_31_V_read32_reg_9521_pp0_iter7_reg <= data_31_V_read32_reg_9521_pp0_iter6_reg;
        data_31_V_read32_reg_9521_pp0_iter8_reg <= data_31_V_read32_reg_9521_pp0_iter7_reg;
        data_31_V_read32_reg_9521_pp0_iter9_reg <= data_31_V_read32_reg_9521_pp0_iter8_reg;
        data_32_V_read_3_reg_9492 <= data_32_V_read_int_reg;
        data_32_V_read_3_reg_9492_pp0_iter1_reg <= data_32_V_read_3_reg_9492;
        data_32_V_read_3_reg_9492_pp0_iter2_reg <= data_32_V_read_3_reg_9492_pp0_iter1_reg;
        data_32_V_read_3_reg_9492_pp0_iter3_reg <= data_32_V_read_3_reg_9492_pp0_iter2_reg;
        data_32_V_read_3_reg_9492_pp0_iter4_reg <= data_32_V_read_3_reg_9492_pp0_iter3_reg;
        data_32_V_read_3_reg_9492_pp0_iter5_reg <= data_32_V_read_3_reg_9492_pp0_iter4_reg;
        data_32_V_read_3_reg_9492_pp0_iter6_reg <= data_32_V_read_3_reg_9492_pp0_iter5_reg;
        data_32_V_read_3_reg_9492_pp0_iter7_reg <= data_32_V_read_3_reg_9492_pp0_iter6_reg;
        data_32_V_read_3_reg_9492_pp0_iter8_reg <= data_32_V_read_3_reg_9492_pp0_iter7_reg;
        data_32_V_read_3_reg_9492_pp0_iter9_reg <= data_32_V_read_3_reg_9492_pp0_iter8_reg;
        data_33_V_read_3_reg_9463 <= data_33_V_read_int_reg;
        data_33_V_read_3_reg_9463_pp0_iter10_reg <= data_33_V_read_3_reg_9463_pp0_iter9_reg;
        data_33_V_read_3_reg_9463_pp0_iter1_reg <= data_33_V_read_3_reg_9463;
        data_33_V_read_3_reg_9463_pp0_iter2_reg <= data_33_V_read_3_reg_9463_pp0_iter1_reg;
        data_33_V_read_3_reg_9463_pp0_iter3_reg <= data_33_V_read_3_reg_9463_pp0_iter2_reg;
        data_33_V_read_3_reg_9463_pp0_iter4_reg <= data_33_V_read_3_reg_9463_pp0_iter3_reg;
        data_33_V_read_3_reg_9463_pp0_iter5_reg <= data_33_V_read_3_reg_9463_pp0_iter4_reg;
        data_33_V_read_3_reg_9463_pp0_iter6_reg <= data_33_V_read_3_reg_9463_pp0_iter5_reg;
        data_33_V_read_3_reg_9463_pp0_iter7_reg <= data_33_V_read_3_reg_9463_pp0_iter6_reg;
        data_33_V_read_3_reg_9463_pp0_iter8_reg <= data_33_V_read_3_reg_9463_pp0_iter7_reg;
        data_33_V_read_3_reg_9463_pp0_iter9_reg <= data_33_V_read_3_reg_9463_pp0_iter8_reg;
        data_34_V_read_3_reg_9434 <= data_34_V_read_int_reg;
        data_34_V_read_3_reg_9434_pp0_iter10_reg <= data_34_V_read_3_reg_9434_pp0_iter9_reg;
        data_34_V_read_3_reg_9434_pp0_iter1_reg <= data_34_V_read_3_reg_9434;
        data_34_V_read_3_reg_9434_pp0_iter2_reg <= data_34_V_read_3_reg_9434_pp0_iter1_reg;
        data_34_V_read_3_reg_9434_pp0_iter3_reg <= data_34_V_read_3_reg_9434_pp0_iter2_reg;
        data_34_V_read_3_reg_9434_pp0_iter4_reg <= data_34_V_read_3_reg_9434_pp0_iter3_reg;
        data_34_V_read_3_reg_9434_pp0_iter5_reg <= data_34_V_read_3_reg_9434_pp0_iter4_reg;
        data_34_V_read_3_reg_9434_pp0_iter6_reg <= data_34_V_read_3_reg_9434_pp0_iter5_reg;
        data_34_V_read_3_reg_9434_pp0_iter7_reg <= data_34_V_read_3_reg_9434_pp0_iter6_reg;
        data_34_V_read_3_reg_9434_pp0_iter8_reg <= data_34_V_read_3_reg_9434_pp0_iter7_reg;
        data_34_V_read_3_reg_9434_pp0_iter9_reg <= data_34_V_read_3_reg_9434_pp0_iter8_reg;
        data_35_V_read_3_reg_9410 <= data_35_V_read_int_reg;
        data_35_V_read_3_reg_9410_pp0_iter10_reg <= data_35_V_read_3_reg_9410_pp0_iter9_reg;
        data_35_V_read_3_reg_9410_pp0_iter1_reg <= data_35_V_read_3_reg_9410;
        data_35_V_read_3_reg_9410_pp0_iter2_reg <= data_35_V_read_3_reg_9410_pp0_iter1_reg;
        data_35_V_read_3_reg_9410_pp0_iter3_reg <= data_35_V_read_3_reg_9410_pp0_iter2_reg;
        data_35_V_read_3_reg_9410_pp0_iter4_reg <= data_35_V_read_3_reg_9410_pp0_iter3_reg;
        data_35_V_read_3_reg_9410_pp0_iter5_reg <= data_35_V_read_3_reg_9410_pp0_iter4_reg;
        data_35_V_read_3_reg_9410_pp0_iter6_reg <= data_35_V_read_3_reg_9410_pp0_iter5_reg;
        data_35_V_read_3_reg_9410_pp0_iter7_reg <= data_35_V_read_3_reg_9410_pp0_iter6_reg;
        data_35_V_read_3_reg_9410_pp0_iter8_reg <= data_35_V_read_3_reg_9410_pp0_iter7_reg;
        data_35_V_read_3_reg_9410_pp0_iter9_reg <= data_35_V_read_3_reg_9410_pp0_iter8_reg;
        data_36_V_read_3_reg_9383 <= data_36_V_read_int_reg;
        data_36_V_read_3_reg_9383_pp0_iter10_reg <= data_36_V_read_3_reg_9383_pp0_iter9_reg;
        data_36_V_read_3_reg_9383_pp0_iter1_reg <= data_36_V_read_3_reg_9383;
        data_36_V_read_3_reg_9383_pp0_iter2_reg <= data_36_V_read_3_reg_9383_pp0_iter1_reg;
        data_36_V_read_3_reg_9383_pp0_iter3_reg <= data_36_V_read_3_reg_9383_pp0_iter2_reg;
        data_36_V_read_3_reg_9383_pp0_iter4_reg <= data_36_V_read_3_reg_9383_pp0_iter3_reg;
        data_36_V_read_3_reg_9383_pp0_iter5_reg <= data_36_V_read_3_reg_9383_pp0_iter4_reg;
        data_36_V_read_3_reg_9383_pp0_iter6_reg <= data_36_V_read_3_reg_9383_pp0_iter5_reg;
        data_36_V_read_3_reg_9383_pp0_iter7_reg <= data_36_V_read_3_reg_9383_pp0_iter6_reg;
        data_36_V_read_3_reg_9383_pp0_iter8_reg <= data_36_V_read_3_reg_9383_pp0_iter7_reg;
        data_36_V_read_3_reg_9383_pp0_iter9_reg <= data_36_V_read_3_reg_9383_pp0_iter8_reg;
        data_37_V_read_3_reg_9353 <= data_37_V_read_int_reg;
        data_37_V_read_3_reg_9353_pp0_iter10_reg <= data_37_V_read_3_reg_9353_pp0_iter9_reg;
        data_37_V_read_3_reg_9353_pp0_iter1_reg <= data_37_V_read_3_reg_9353;
        data_37_V_read_3_reg_9353_pp0_iter2_reg <= data_37_V_read_3_reg_9353_pp0_iter1_reg;
        data_37_V_read_3_reg_9353_pp0_iter3_reg <= data_37_V_read_3_reg_9353_pp0_iter2_reg;
        data_37_V_read_3_reg_9353_pp0_iter4_reg <= data_37_V_read_3_reg_9353_pp0_iter3_reg;
        data_37_V_read_3_reg_9353_pp0_iter5_reg <= data_37_V_read_3_reg_9353_pp0_iter4_reg;
        data_37_V_read_3_reg_9353_pp0_iter6_reg <= data_37_V_read_3_reg_9353_pp0_iter5_reg;
        data_37_V_read_3_reg_9353_pp0_iter7_reg <= data_37_V_read_3_reg_9353_pp0_iter6_reg;
        data_37_V_read_3_reg_9353_pp0_iter8_reg <= data_37_V_read_3_reg_9353_pp0_iter7_reg;
        data_37_V_read_3_reg_9353_pp0_iter9_reg <= data_37_V_read_3_reg_9353_pp0_iter8_reg;
        data_38_V_read_3_reg_9328 <= data_38_V_read_int_reg;
        data_38_V_read_3_reg_9328_pp0_iter10_reg <= data_38_V_read_3_reg_9328_pp0_iter9_reg;
        data_38_V_read_3_reg_9328_pp0_iter11_reg <= data_38_V_read_3_reg_9328_pp0_iter10_reg;
        data_38_V_read_3_reg_9328_pp0_iter1_reg <= data_38_V_read_3_reg_9328;
        data_38_V_read_3_reg_9328_pp0_iter2_reg <= data_38_V_read_3_reg_9328_pp0_iter1_reg;
        data_38_V_read_3_reg_9328_pp0_iter3_reg <= data_38_V_read_3_reg_9328_pp0_iter2_reg;
        data_38_V_read_3_reg_9328_pp0_iter4_reg <= data_38_V_read_3_reg_9328_pp0_iter3_reg;
        data_38_V_read_3_reg_9328_pp0_iter5_reg <= data_38_V_read_3_reg_9328_pp0_iter4_reg;
        data_38_V_read_3_reg_9328_pp0_iter6_reg <= data_38_V_read_3_reg_9328_pp0_iter5_reg;
        data_38_V_read_3_reg_9328_pp0_iter7_reg <= data_38_V_read_3_reg_9328_pp0_iter6_reg;
        data_38_V_read_3_reg_9328_pp0_iter8_reg <= data_38_V_read_3_reg_9328_pp0_iter7_reg;
        data_38_V_read_3_reg_9328_pp0_iter9_reg <= data_38_V_read_3_reg_9328_pp0_iter8_reg;
        data_39_V_read_3_reg_9301 <= data_39_V_read_int_reg;
        data_39_V_read_3_reg_9301_pp0_iter10_reg <= data_39_V_read_3_reg_9301_pp0_iter9_reg;
        data_39_V_read_3_reg_9301_pp0_iter11_reg <= data_39_V_read_3_reg_9301_pp0_iter10_reg;
        data_39_V_read_3_reg_9301_pp0_iter1_reg <= data_39_V_read_3_reg_9301;
        data_39_V_read_3_reg_9301_pp0_iter2_reg <= data_39_V_read_3_reg_9301_pp0_iter1_reg;
        data_39_V_read_3_reg_9301_pp0_iter3_reg <= data_39_V_read_3_reg_9301_pp0_iter2_reg;
        data_39_V_read_3_reg_9301_pp0_iter4_reg <= data_39_V_read_3_reg_9301_pp0_iter3_reg;
        data_39_V_read_3_reg_9301_pp0_iter5_reg <= data_39_V_read_3_reg_9301_pp0_iter4_reg;
        data_39_V_read_3_reg_9301_pp0_iter6_reg <= data_39_V_read_3_reg_9301_pp0_iter5_reg;
        data_39_V_read_3_reg_9301_pp0_iter7_reg <= data_39_V_read_3_reg_9301_pp0_iter6_reg;
        data_39_V_read_3_reg_9301_pp0_iter8_reg <= data_39_V_read_3_reg_9301_pp0_iter7_reg;
        data_39_V_read_3_reg_9301_pp0_iter9_reg <= data_39_V_read_3_reg_9301_pp0_iter8_reg;
        data_3_V_read_10_reg_10295 <= data_3_V_read_int_reg;
        data_3_V_read_10_reg_10295_pp0_iter1_reg <= data_3_V_read_10_reg_10295;
        data_3_V_read_10_reg_10295_pp0_iter2_reg <= data_3_V_read_10_reg_10295_pp0_iter1_reg;
        data_40_V_read41_reg_9272 <= data_40_V_read_int_reg;
        data_40_V_read41_reg_9272_pp0_iter10_reg <= data_40_V_read41_reg_9272_pp0_iter9_reg;
        data_40_V_read41_reg_9272_pp0_iter11_reg <= data_40_V_read41_reg_9272_pp0_iter10_reg;
        data_40_V_read41_reg_9272_pp0_iter1_reg <= data_40_V_read41_reg_9272;
        data_40_V_read41_reg_9272_pp0_iter2_reg <= data_40_V_read41_reg_9272_pp0_iter1_reg;
        data_40_V_read41_reg_9272_pp0_iter3_reg <= data_40_V_read41_reg_9272_pp0_iter2_reg;
        data_40_V_read41_reg_9272_pp0_iter4_reg <= data_40_V_read41_reg_9272_pp0_iter3_reg;
        data_40_V_read41_reg_9272_pp0_iter5_reg <= data_40_V_read41_reg_9272_pp0_iter4_reg;
        data_40_V_read41_reg_9272_pp0_iter6_reg <= data_40_V_read41_reg_9272_pp0_iter5_reg;
        data_40_V_read41_reg_9272_pp0_iter7_reg <= data_40_V_read41_reg_9272_pp0_iter6_reg;
        data_40_V_read41_reg_9272_pp0_iter8_reg <= data_40_V_read41_reg_9272_pp0_iter7_reg;
        data_40_V_read41_reg_9272_pp0_iter9_reg <= data_40_V_read41_reg_9272_pp0_iter8_reg;
        data_41_V_read42_reg_9242 <= data_41_V_read_int_reg;
        data_41_V_read42_reg_9242_pp0_iter10_reg <= data_41_V_read42_reg_9242_pp0_iter9_reg;
        data_41_V_read42_reg_9242_pp0_iter11_reg <= data_41_V_read42_reg_9242_pp0_iter10_reg;
        data_41_V_read42_reg_9242_pp0_iter1_reg <= data_41_V_read42_reg_9242;
        data_41_V_read42_reg_9242_pp0_iter2_reg <= data_41_V_read42_reg_9242_pp0_iter1_reg;
        data_41_V_read42_reg_9242_pp0_iter3_reg <= data_41_V_read42_reg_9242_pp0_iter2_reg;
        data_41_V_read42_reg_9242_pp0_iter4_reg <= data_41_V_read42_reg_9242_pp0_iter3_reg;
        data_41_V_read42_reg_9242_pp0_iter5_reg <= data_41_V_read42_reg_9242_pp0_iter4_reg;
        data_41_V_read42_reg_9242_pp0_iter6_reg <= data_41_V_read42_reg_9242_pp0_iter5_reg;
        data_41_V_read42_reg_9242_pp0_iter7_reg <= data_41_V_read42_reg_9242_pp0_iter6_reg;
        data_41_V_read42_reg_9242_pp0_iter8_reg <= data_41_V_read42_reg_9242_pp0_iter7_reg;
        data_41_V_read42_reg_9242_pp0_iter9_reg <= data_41_V_read42_reg_9242_pp0_iter8_reg;
        data_42_V_read_3_reg_9212 <= data_42_V_read_int_reg;
        data_42_V_read_3_reg_9212_pp0_iter10_reg <= data_42_V_read_3_reg_9212_pp0_iter9_reg;
        data_42_V_read_3_reg_9212_pp0_iter11_reg <= data_42_V_read_3_reg_9212_pp0_iter10_reg;
        data_42_V_read_3_reg_9212_pp0_iter12_reg <= data_42_V_read_3_reg_9212_pp0_iter11_reg;
        data_42_V_read_3_reg_9212_pp0_iter1_reg <= data_42_V_read_3_reg_9212;
        data_42_V_read_3_reg_9212_pp0_iter2_reg <= data_42_V_read_3_reg_9212_pp0_iter1_reg;
        data_42_V_read_3_reg_9212_pp0_iter3_reg <= data_42_V_read_3_reg_9212_pp0_iter2_reg;
        data_42_V_read_3_reg_9212_pp0_iter4_reg <= data_42_V_read_3_reg_9212_pp0_iter3_reg;
        data_42_V_read_3_reg_9212_pp0_iter5_reg <= data_42_V_read_3_reg_9212_pp0_iter4_reg;
        data_42_V_read_3_reg_9212_pp0_iter6_reg <= data_42_V_read_3_reg_9212_pp0_iter5_reg;
        data_42_V_read_3_reg_9212_pp0_iter7_reg <= data_42_V_read_3_reg_9212_pp0_iter6_reg;
        data_42_V_read_3_reg_9212_pp0_iter8_reg <= data_42_V_read_3_reg_9212_pp0_iter7_reg;
        data_42_V_read_3_reg_9212_pp0_iter9_reg <= data_42_V_read_3_reg_9212_pp0_iter8_reg;
        data_43_V_read_3_reg_9184 <= data_43_V_read_int_reg;
        data_43_V_read_3_reg_9184_pp0_iter10_reg <= data_43_V_read_3_reg_9184_pp0_iter9_reg;
        data_43_V_read_3_reg_9184_pp0_iter11_reg <= data_43_V_read_3_reg_9184_pp0_iter10_reg;
        data_43_V_read_3_reg_9184_pp0_iter12_reg <= data_43_V_read_3_reg_9184_pp0_iter11_reg;
        data_43_V_read_3_reg_9184_pp0_iter1_reg <= data_43_V_read_3_reg_9184;
        data_43_V_read_3_reg_9184_pp0_iter2_reg <= data_43_V_read_3_reg_9184_pp0_iter1_reg;
        data_43_V_read_3_reg_9184_pp0_iter3_reg <= data_43_V_read_3_reg_9184_pp0_iter2_reg;
        data_43_V_read_3_reg_9184_pp0_iter4_reg <= data_43_V_read_3_reg_9184_pp0_iter3_reg;
        data_43_V_read_3_reg_9184_pp0_iter5_reg <= data_43_V_read_3_reg_9184_pp0_iter4_reg;
        data_43_V_read_3_reg_9184_pp0_iter6_reg <= data_43_V_read_3_reg_9184_pp0_iter5_reg;
        data_43_V_read_3_reg_9184_pp0_iter7_reg <= data_43_V_read_3_reg_9184_pp0_iter6_reg;
        data_43_V_read_3_reg_9184_pp0_iter8_reg <= data_43_V_read_3_reg_9184_pp0_iter7_reg;
        data_43_V_read_3_reg_9184_pp0_iter9_reg <= data_43_V_read_3_reg_9184_pp0_iter8_reg;
        data_44_V_read_3_reg_9154 <= data_44_V_read_int_reg;
        data_44_V_read_3_reg_9154_pp0_iter10_reg <= data_44_V_read_3_reg_9154_pp0_iter9_reg;
        data_44_V_read_3_reg_9154_pp0_iter11_reg <= data_44_V_read_3_reg_9154_pp0_iter10_reg;
        data_44_V_read_3_reg_9154_pp0_iter12_reg <= data_44_V_read_3_reg_9154_pp0_iter11_reg;
        data_44_V_read_3_reg_9154_pp0_iter1_reg <= data_44_V_read_3_reg_9154;
        data_44_V_read_3_reg_9154_pp0_iter2_reg <= data_44_V_read_3_reg_9154_pp0_iter1_reg;
        data_44_V_read_3_reg_9154_pp0_iter3_reg <= data_44_V_read_3_reg_9154_pp0_iter2_reg;
        data_44_V_read_3_reg_9154_pp0_iter4_reg <= data_44_V_read_3_reg_9154_pp0_iter3_reg;
        data_44_V_read_3_reg_9154_pp0_iter5_reg <= data_44_V_read_3_reg_9154_pp0_iter4_reg;
        data_44_V_read_3_reg_9154_pp0_iter6_reg <= data_44_V_read_3_reg_9154_pp0_iter5_reg;
        data_44_V_read_3_reg_9154_pp0_iter7_reg <= data_44_V_read_3_reg_9154_pp0_iter6_reg;
        data_44_V_read_3_reg_9154_pp0_iter8_reg <= data_44_V_read_3_reg_9154_pp0_iter7_reg;
        data_44_V_read_3_reg_9154_pp0_iter9_reg <= data_44_V_read_3_reg_9154_pp0_iter8_reg;
        data_45_V_read_3_reg_9125 <= data_45_V_read_int_reg;
        data_45_V_read_3_reg_9125_pp0_iter10_reg <= data_45_V_read_3_reg_9125_pp0_iter9_reg;
        data_45_V_read_3_reg_9125_pp0_iter11_reg <= data_45_V_read_3_reg_9125_pp0_iter10_reg;
        data_45_V_read_3_reg_9125_pp0_iter12_reg <= data_45_V_read_3_reg_9125_pp0_iter11_reg;
        data_45_V_read_3_reg_9125_pp0_iter1_reg <= data_45_V_read_3_reg_9125;
        data_45_V_read_3_reg_9125_pp0_iter2_reg <= data_45_V_read_3_reg_9125_pp0_iter1_reg;
        data_45_V_read_3_reg_9125_pp0_iter3_reg <= data_45_V_read_3_reg_9125_pp0_iter2_reg;
        data_45_V_read_3_reg_9125_pp0_iter4_reg <= data_45_V_read_3_reg_9125_pp0_iter3_reg;
        data_45_V_read_3_reg_9125_pp0_iter5_reg <= data_45_V_read_3_reg_9125_pp0_iter4_reg;
        data_45_V_read_3_reg_9125_pp0_iter6_reg <= data_45_V_read_3_reg_9125_pp0_iter5_reg;
        data_45_V_read_3_reg_9125_pp0_iter7_reg <= data_45_V_read_3_reg_9125_pp0_iter6_reg;
        data_45_V_read_3_reg_9125_pp0_iter8_reg <= data_45_V_read_3_reg_9125_pp0_iter7_reg;
        data_45_V_read_3_reg_9125_pp0_iter9_reg <= data_45_V_read_3_reg_9125_pp0_iter8_reg;
        data_46_V_read_3_reg_9094 <= data_46_V_read_int_reg;
        data_46_V_read_3_reg_9094_pp0_iter10_reg <= data_46_V_read_3_reg_9094_pp0_iter9_reg;
        data_46_V_read_3_reg_9094_pp0_iter11_reg <= data_46_V_read_3_reg_9094_pp0_iter10_reg;
        data_46_V_read_3_reg_9094_pp0_iter12_reg <= data_46_V_read_3_reg_9094_pp0_iter11_reg;
        data_46_V_read_3_reg_9094_pp0_iter13_reg <= data_46_V_read_3_reg_9094_pp0_iter12_reg;
        data_46_V_read_3_reg_9094_pp0_iter1_reg <= data_46_V_read_3_reg_9094;
        data_46_V_read_3_reg_9094_pp0_iter2_reg <= data_46_V_read_3_reg_9094_pp0_iter1_reg;
        data_46_V_read_3_reg_9094_pp0_iter3_reg <= data_46_V_read_3_reg_9094_pp0_iter2_reg;
        data_46_V_read_3_reg_9094_pp0_iter4_reg <= data_46_V_read_3_reg_9094_pp0_iter3_reg;
        data_46_V_read_3_reg_9094_pp0_iter5_reg <= data_46_V_read_3_reg_9094_pp0_iter4_reg;
        data_46_V_read_3_reg_9094_pp0_iter6_reg <= data_46_V_read_3_reg_9094_pp0_iter5_reg;
        data_46_V_read_3_reg_9094_pp0_iter7_reg <= data_46_V_read_3_reg_9094_pp0_iter6_reg;
        data_46_V_read_3_reg_9094_pp0_iter8_reg <= data_46_V_read_3_reg_9094_pp0_iter7_reg;
        data_46_V_read_3_reg_9094_pp0_iter9_reg <= data_46_V_read_3_reg_9094_pp0_iter8_reg;
        data_47_V_read_3_reg_9066 <= data_47_V_read_int_reg;
        data_47_V_read_3_reg_9066_pp0_iter10_reg <= data_47_V_read_3_reg_9066_pp0_iter9_reg;
        data_47_V_read_3_reg_9066_pp0_iter11_reg <= data_47_V_read_3_reg_9066_pp0_iter10_reg;
        data_47_V_read_3_reg_9066_pp0_iter12_reg <= data_47_V_read_3_reg_9066_pp0_iter11_reg;
        data_47_V_read_3_reg_9066_pp0_iter13_reg <= data_47_V_read_3_reg_9066_pp0_iter12_reg;
        data_47_V_read_3_reg_9066_pp0_iter1_reg <= data_47_V_read_3_reg_9066;
        data_47_V_read_3_reg_9066_pp0_iter2_reg <= data_47_V_read_3_reg_9066_pp0_iter1_reg;
        data_47_V_read_3_reg_9066_pp0_iter3_reg <= data_47_V_read_3_reg_9066_pp0_iter2_reg;
        data_47_V_read_3_reg_9066_pp0_iter4_reg <= data_47_V_read_3_reg_9066_pp0_iter3_reg;
        data_47_V_read_3_reg_9066_pp0_iter5_reg <= data_47_V_read_3_reg_9066_pp0_iter4_reg;
        data_47_V_read_3_reg_9066_pp0_iter6_reg <= data_47_V_read_3_reg_9066_pp0_iter5_reg;
        data_47_V_read_3_reg_9066_pp0_iter7_reg <= data_47_V_read_3_reg_9066_pp0_iter6_reg;
        data_47_V_read_3_reg_9066_pp0_iter8_reg <= data_47_V_read_3_reg_9066_pp0_iter7_reg;
        data_47_V_read_3_reg_9066_pp0_iter9_reg <= data_47_V_read_3_reg_9066_pp0_iter8_reg;
        data_48_V_read_3_reg_9040 <= data_48_V_read_int_reg;
        data_48_V_read_3_reg_9040_pp0_iter10_reg <= data_48_V_read_3_reg_9040_pp0_iter9_reg;
        data_48_V_read_3_reg_9040_pp0_iter11_reg <= data_48_V_read_3_reg_9040_pp0_iter10_reg;
        data_48_V_read_3_reg_9040_pp0_iter12_reg <= data_48_V_read_3_reg_9040_pp0_iter11_reg;
        data_48_V_read_3_reg_9040_pp0_iter13_reg <= data_48_V_read_3_reg_9040_pp0_iter12_reg;
        data_48_V_read_3_reg_9040_pp0_iter1_reg <= data_48_V_read_3_reg_9040;
        data_48_V_read_3_reg_9040_pp0_iter2_reg <= data_48_V_read_3_reg_9040_pp0_iter1_reg;
        data_48_V_read_3_reg_9040_pp0_iter3_reg <= data_48_V_read_3_reg_9040_pp0_iter2_reg;
        data_48_V_read_3_reg_9040_pp0_iter4_reg <= data_48_V_read_3_reg_9040_pp0_iter3_reg;
        data_48_V_read_3_reg_9040_pp0_iter5_reg <= data_48_V_read_3_reg_9040_pp0_iter4_reg;
        data_48_V_read_3_reg_9040_pp0_iter6_reg <= data_48_V_read_3_reg_9040_pp0_iter5_reg;
        data_48_V_read_3_reg_9040_pp0_iter7_reg <= data_48_V_read_3_reg_9040_pp0_iter6_reg;
        data_48_V_read_3_reg_9040_pp0_iter8_reg <= data_48_V_read_3_reg_9040_pp0_iter7_reg;
        data_48_V_read_3_reg_9040_pp0_iter9_reg <= data_48_V_read_3_reg_9040_pp0_iter8_reg;
        data_49_V_read_3_reg_9012 <= data_49_V_read_int_reg;
        data_49_V_read_3_reg_9012_pp0_iter10_reg <= data_49_V_read_3_reg_9012_pp0_iter9_reg;
        data_49_V_read_3_reg_9012_pp0_iter11_reg <= data_49_V_read_3_reg_9012_pp0_iter10_reg;
        data_49_V_read_3_reg_9012_pp0_iter12_reg <= data_49_V_read_3_reg_9012_pp0_iter11_reg;
        data_49_V_read_3_reg_9012_pp0_iter13_reg <= data_49_V_read_3_reg_9012_pp0_iter12_reg;
        data_49_V_read_3_reg_9012_pp0_iter1_reg <= data_49_V_read_3_reg_9012;
        data_49_V_read_3_reg_9012_pp0_iter2_reg <= data_49_V_read_3_reg_9012_pp0_iter1_reg;
        data_49_V_read_3_reg_9012_pp0_iter3_reg <= data_49_V_read_3_reg_9012_pp0_iter2_reg;
        data_49_V_read_3_reg_9012_pp0_iter4_reg <= data_49_V_read_3_reg_9012_pp0_iter3_reg;
        data_49_V_read_3_reg_9012_pp0_iter5_reg <= data_49_V_read_3_reg_9012_pp0_iter4_reg;
        data_49_V_read_3_reg_9012_pp0_iter6_reg <= data_49_V_read_3_reg_9012_pp0_iter5_reg;
        data_49_V_read_3_reg_9012_pp0_iter7_reg <= data_49_V_read_3_reg_9012_pp0_iter6_reg;
        data_49_V_read_3_reg_9012_pp0_iter8_reg <= data_49_V_read_3_reg_9012_pp0_iter7_reg;
        data_49_V_read_3_reg_9012_pp0_iter9_reg <= data_49_V_read_3_reg_9012_pp0_iter8_reg;
        data_4_V_read_10_reg_10273 <= data_4_V_read_int_reg;
        data_4_V_read_10_reg_10273_pp0_iter1_reg <= data_4_V_read_10_reg_10273;
        data_4_V_read_10_reg_10273_pp0_iter2_reg <= data_4_V_read_10_reg_10273_pp0_iter1_reg;
        data_4_V_read_10_reg_10273_pp0_iter3_reg <= data_4_V_read_10_reg_10273_pp0_iter2_reg;
        data_50_V_read51_reg_8984 <= data_50_V_read_int_reg;
        data_50_V_read51_reg_8984_pp0_iter10_reg <= data_50_V_read51_reg_8984_pp0_iter9_reg;
        data_50_V_read51_reg_8984_pp0_iter11_reg <= data_50_V_read51_reg_8984_pp0_iter10_reg;
        data_50_V_read51_reg_8984_pp0_iter12_reg <= data_50_V_read51_reg_8984_pp0_iter11_reg;
        data_50_V_read51_reg_8984_pp0_iter13_reg <= data_50_V_read51_reg_8984_pp0_iter12_reg;
        data_50_V_read51_reg_8984_pp0_iter14_reg <= data_50_V_read51_reg_8984_pp0_iter13_reg;
        data_50_V_read51_reg_8984_pp0_iter1_reg <= data_50_V_read51_reg_8984;
        data_50_V_read51_reg_8984_pp0_iter2_reg <= data_50_V_read51_reg_8984_pp0_iter1_reg;
        data_50_V_read51_reg_8984_pp0_iter3_reg <= data_50_V_read51_reg_8984_pp0_iter2_reg;
        data_50_V_read51_reg_8984_pp0_iter4_reg <= data_50_V_read51_reg_8984_pp0_iter3_reg;
        data_50_V_read51_reg_8984_pp0_iter5_reg <= data_50_V_read51_reg_8984_pp0_iter4_reg;
        data_50_V_read51_reg_8984_pp0_iter6_reg <= data_50_V_read51_reg_8984_pp0_iter5_reg;
        data_50_V_read51_reg_8984_pp0_iter7_reg <= data_50_V_read51_reg_8984_pp0_iter6_reg;
        data_50_V_read51_reg_8984_pp0_iter8_reg <= data_50_V_read51_reg_8984_pp0_iter7_reg;
        data_50_V_read51_reg_8984_pp0_iter9_reg <= data_50_V_read51_reg_8984_pp0_iter8_reg;
        data_51_V_read52_reg_8956 <= data_51_V_read_int_reg;
        data_51_V_read52_reg_8956_pp0_iter10_reg <= data_51_V_read52_reg_8956_pp0_iter9_reg;
        data_51_V_read52_reg_8956_pp0_iter11_reg <= data_51_V_read52_reg_8956_pp0_iter10_reg;
        data_51_V_read52_reg_8956_pp0_iter12_reg <= data_51_V_read52_reg_8956_pp0_iter11_reg;
        data_51_V_read52_reg_8956_pp0_iter13_reg <= data_51_V_read52_reg_8956_pp0_iter12_reg;
        data_51_V_read52_reg_8956_pp0_iter14_reg <= data_51_V_read52_reg_8956_pp0_iter13_reg;
        data_51_V_read52_reg_8956_pp0_iter1_reg <= data_51_V_read52_reg_8956;
        data_51_V_read52_reg_8956_pp0_iter2_reg <= data_51_V_read52_reg_8956_pp0_iter1_reg;
        data_51_V_read52_reg_8956_pp0_iter3_reg <= data_51_V_read52_reg_8956_pp0_iter2_reg;
        data_51_V_read52_reg_8956_pp0_iter4_reg <= data_51_V_read52_reg_8956_pp0_iter3_reg;
        data_51_V_read52_reg_8956_pp0_iter5_reg <= data_51_V_read52_reg_8956_pp0_iter4_reg;
        data_51_V_read52_reg_8956_pp0_iter6_reg <= data_51_V_read52_reg_8956_pp0_iter5_reg;
        data_51_V_read52_reg_8956_pp0_iter7_reg <= data_51_V_read52_reg_8956_pp0_iter6_reg;
        data_51_V_read52_reg_8956_pp0_iter8_reg <= data_51_V_read52_reg_8956_pp0_iter7_reg;
        data_51_V_read52_reg_8956_pp0_iter9_reg <= data_51_V_read52_reg_8956_pp0_iter8_reg;
        data_52_V_read_3_reg_8928 <= data_52_V_read_int_reg;
        data_52_V_read_3_reg_8928_pp0_iter10_reg <= data_52_V_read_3_reg_8928_pp0_iter9_reg;
        data_52_V_read_3_reg_8928_pp0_iter11_reg <= data_52_V_read_3_reg_8928_pp0_iter10_reg;
        data_52_V_read_3_reg_8928_pp0_iter12_reg <= data_52_V_read_3_reg_8928_pp0_iter11_reg;
        data_52_V_read_3_reg_8928_pp0_iter13_reg <= data_52_V_read_3_reg_8928_pp0_iter12_reg;
        data_52_V_read_3_reg_8928_pp0_iter14_reg <= data_52_V_read_3_reg_8928_pp0_iter13_reg;
        data_52_V_read_3_reg_8928_pp0_iter1_reg <= data_52_V_read_3_reg_8928;
        data_52_V_read_3_reg_8928_pp0_iter2_reg <= data_52_V_read_3_reg_8928_pp0_iter1_reg;
        data_52_V_read_3_reg_8928_pp0_iter3_reg <= data_52_V_read_3_reg_8928_pp0_iter2_reg;
        data_52_V_read_3_reg_8928_pp0_iter4_reg <= data_52_V_read_3_reg_8928_pp0_iter3_reg;
        data_52_V_read_3_reg_8928_pp0_iter5_reg <= data_52_V_read_3_reg_8928_pp0_iter4_reg;
        data_52_V_read_3_reg_8928_pp0_iter6_reg <= data_52_V_read_3_reg_8928_pp0_iter5_reg;
        data_52_V_read_3_reg_8928_pp0_iter7_reg <= data_52_V_read_3_reg_8928_pp0_iter6_reg;
        data_52_V_read_3_reg_8928_pp0_iter8_reg <= data_52_V_read_3_reg_8928_pp0_iter7_reg;
        data_52_V_read_3_reg_8928_pp0_iter9_reg <= data_52_V_read_3_reg_8928_pp0_iter8_reg;
        data_53_V_read_3_reg_8899 <= data_53_V_read_int_reg;
        data_53_V_read_3_reg_8899_pp0_iter10_reg <= data_53_V_read_3_reg_8899_pp0_iter9_reg;
        data_53_V_read_3_reg_8899_pp0_iter11_reg <= data_53_V_read_3_reg_8899_pp0_iter10_reg;
        data_53_V_read_3_reg_8899_pp0_iter12_reg <= data_53_V_read_3_reg_8899_pp0_iter11_reg;
        data_53_V_read_3_reg_8899_pp0_iter13_reg <= data_53_V_read_3_reg_8899_pp0_iter12_reg;
        data_53_V_read_3_reg_8899_pp0_iter14_reg <= data_53_V_read_3_reg_8899_pp0_iter13_reg;
        data_53_V_read_3_reg_8899_pp0_iter1_reg <= data_53_V_read_3_reg_8899;
        data_53_V_read_3_reg_8899_pp0_iter2_reg <= data_53_V_read_3_reg_8899_pp0_iter1_reg;
        data_53_V_read_3_reg_8899_pp0_iter3_reg <= data_53_V_read_3_reg_8899_pp0_iter2_reg;
        data_53_V_read_3_reg_8899_pp0_iter4_reg <= data_53_V_read_3_reg_8899_pp0_iter3_reg;
        data_53_V_read_3_reg_8899_pp0_iter5_reg <= data_53_V_read_3_reg_8899_pp0_iter4_reg;
        data_53_V_read_3_reg_8899_pp0_iter6_reg <= data_53_V_read_3_reg_8899_pp0_iter5_reg;
        data_53_V_read_3_reg_8899_pp0_iter7_reg <= data_53_V_read_3_reg_8899_pp0_iter6_reg;
        data_53_V_read_3_reg_8899_pp0_iter8_reg <= data_53_V_read_3_reg_8899_pp0_iter7_reg;
        data_53_V_read_3_reg_8899_pp0_iter9_reg <= data_53_V_read_3_reg_8899_pp0_iter8_reg;
        data_54_V_read_3_reg_8873 <= data_54_V_read_int_reg;
        data_54_V_read_3_reg_8873_pp0_iter10_reg <= data_54_V_read_3_reg_8873_pp0_iter9_reg;
        data_54_V_read_3_reg_8873_pp0_iter11_reg <= data_54_V_read_3_reg_8873_pp0_iter10_reg;
        data_54_V_read_3_reg_8873_pp0_iter12_reg <= data_54_V_read_3_reg_8873_pp0_iter11_reg;
        data_54_V_read_3_reg_8873_pp0_iter13_reg <= data_54_V_read_3_reg_8873_pp0_iter12_reg;
        data_54_V_read_3_reg_8873_pp0_iter14_reg <= data_54_V_read_3_reg_8873_pp0_iter13_reg;
        data_54_V_read_3_reg_8873_pp0_iter1_reg <= data_54_V_read_3_reg_8873;
        data_54_V_read_3_reg_8873_pp0_iter2_reg <= data_54_V_read_3_reg_8873_pp0_iter1_reg;
        data_54_V_read_3_reg_8873_pp0_iter3_reg <= data_54_V_read_3_reg_8873_pp0_iter2_reg;
        data_54_V_read_3_reg_8873_pp0_iter4_reg <= data_54_V_read_3_reg_8873_pp0_iter3_reg;
        data_54_V_read_3_reg_8873_pp0_iter5_reg <= data_54_V_read_3_reg_8873_pp0_iter4_reg;
        data_54_V_read_3_reg_8873_pp0_iter6_reg <= data_54_V_read_3_reg_8873_pp0_iter5_reg;
        data_54_V_read_3_reg_8873_pp0_iter7_reg <= data_54_V_read_3_reg_8873_pp0_iter6_reg;
        data_54_V_read_3_reg_8873_pp0_iter8_reg <= data_54_V_read_3_reg_8873_pp0_iter7_reg;
        data_54_V_read_3_reg_8873_pp0_iter9_reg <= data_54_V_read_3_reg_8873_pp0_iter8_reg;
        data_55_V_read_3_reg_8844 <= data_55_V_read_int_reg;
        data_55_V_read_3_reg_8844_pp0_iter10_reg <= data_55_V_read_3_reg_8844_pp0_iter9_reg;
        data_55_V_read_3_reg_8844_pp0_iter11_reg <= data_55_V_read_3_reg_8844_pp0_iter10_reg;
        data_55_V_read_3_reg_8844_pp0_iter12_reg <= data_55_V_read_3_reg_8844_pp0_iter11_reg;
        data_55_V_read_3_reg_8844_pp0_iter13_reg <= data_55_V_read_3_reg_8844_pp0_iter12_reg;
        data_55_V_read_3_reg_8844_pp0_iter14_reg <= data_55_V_read_3_reg_8844_pp0_iter13_reg;
        data_55_V_read_3_reg_8844_pp0_iter15_reg <= data_55_V_read_3_reg_8844_pp0_iter14_reg;
        data_55_V_read_3_reg_8844_pp0_iter1_reg <= data_55_V_read_3_reg_8844;
        data_55_V_read_3_reg_8844_pp0_iter2_reg <= data_55_V_read_3_reg_8844_pp0_iter1_reg;
        data_55_V_read_3_reg_8844_pp0_iter3_reg <= data_55_V_read_3_reg_8844_pp0_iter2_reg;
        data_55_V_read_3_reg_8844_pp0_iter4_reg <= data_55_V_read_3_reg_8844_pp0_iter3_reg;
        data_55_V_read_3_reg_8844_pp0_iter5_reg <= data_55_V_read_3_reg_8844_pp0_iter4_reg;
        data_55_V_read_3_reg_8844_pp0_iter6_reg <= data_55_V_read_3_reg_8844_pp0_iter5_reg;
        data_55_V_read_3_reg_8844_pp0_iter7_reg <= data_55_V_read_3_reg_8844_pp0_iter6_reg;
        data_55_V_read_3_reg_8844_pp0_iter8_reg <= data_55_V_read_3_reg_8844_pp0_iter7_reg;
        data_55_V_read_3_reg_8844_pp0_iter9_reg <= data_55_V_read_3_reg_8844_pp0_iter8_reg;
        data_56_V_read_3_reg_8814 <= data_56_V_read_int_reg;
        data_56_V_read_3_reg_8814_pp0_iter10_reg <= data_56_V_read_3_reg_8814_pp0_iter9_reg;
        data_56_V_read_3_reg_8814_pp0_iter11_reg <= data_56_V_read_3_reg_8814_pp0_iter10_reg;
        data_56_V_read_3_reg_8814_pp0_iter12_reg <= data_56_V_read_3_reg_8814_pp0_iter11_reg;
        data_56_V_read_3_reg_8814_pp0_iter13_reg <= data_56_V_read_3_reg_8814_pp0_iter12_reg;
        data_56_V_read_3_reg_8814_pp0_iter14_reg <= data_56_V_read_3_reg_8814_pp0_iter13_reg;
        data_56_V_read_3_reg_8814_pp0_iter15_reg <= data_56_V_read_3_reg_8814_pp0_iter14_reg;
        data_56_V_read_3_reg_8814_pp0_iter1_reg <= data_56_V_read_3_reg_8814;
        data_56_V_read_3_reg_8814_pp0_iter2_reg <= data_56_V_read_3_reg_8814_pp0_iter1_reg;
        data_56_V_read_3_reg_8814_pp0_iter3_reg <= data_56_V_read_3_reg_8814_pp0_iter2_reg;
        data_56_V_read_3_reg_8814_pp0_iter4_reg <= data_56_V_read_3_reg_8814_pp0_iter3_reg;
        data_56_V_read_3_reg_8814_pp0_iter5_reg <= data_56_V_read_3_reg_8814_pp0_iter4_reg;
        data_56_V_read_3_reg_8814_pp0_iter6_reg <= data_56_V_read_3_reg_8814_pp0_iter5_reg;
        data_56_V_read_3_reg_8814_pp0_iter7_reg <= data_56_V_read_3_reg_8814_pp0_iter6_reg;
        data_56_V_read_3_reg_8814_pp0_iter8_reg <= data_56_V_read_3_reg_8814_pp0_iter7_reg;
        data_56_V_read_3_reg_8814_pp0_iter9_reg <= data_56_V_read_3_reg_8814_pp0_iter8_reg;
        data_57_V_read_3_reg_8786 <= data_57_V_read_int_reg;
        data_57_V_read_3_reg_8786_pp0_iter10_reg <= data_57_V_read_3_reg_8786_pp0_iter9_reg;
        data_57_V_read_3_reg_8786_pp0_iter11_reg <= data_57_V_read_3_reg_8786_pp0_iter10_reg;
        data_57_V_read_3_reg_8786_pp0_iter12_reg <= data_57_V_read_3_reg_8786_pp0_iter11_reg;
        data_57_V_read_3_reg_8786_pp0_iter13_reg <= data_57_V_read_3_reg_8786_pp0_iter12_reg;
        data_57_V_read_3_reg_8786_pp0_iter14_reg <= data_57_V_read_3_reg_8786_pp0_iter13_reg;
        data_57_V_read_3_reg_8786_pp0_iter15_reg <= data_57_V_read_3_reg_8786_pp0_iter14_reg;
        data_57_V_read_3_reg_8786_pp0_iter1_reg <= data_57_V_read_3_reg_8786;
        data_57_V_read_3_reg_8786_pp0_iter2_reg <= data_57_V_read_3_reg_8786_pp0_iter1_reg;
        data_57_V_read_3_reg_8786_pp0_iter3_reg <= data_57_V_read_3_reg_8786_pp0_iter2_reg;
        data_57_V_read_3_reg_8786_pp0_iter4_reg <= data_57_V_read_3_reg_8786_pp0_iter3_reg;
        data_57_V_read_3_reg_8786_pp0_iter5_reg <= data_57_V_read_3_reg_8786_pp0_iter4_reg;
        data_57_V_read_3_reg_8786_pp0_iter6_reg <= data_57_V_read_3_reg_8786_pp0_iter5_reg;
        data_57_V_read_3_reg_8786_pp0_iter7_reg <= data_57_V_read_3_reg_8786_pp0_iter6_reg;
        data_57_V_read_3_reg_8786_pp0_iter8_reg <= data_57_V_read_3_reg_8786_pp0_iter7_reg;
        data_57_V_read_3_reg_8786_pp0_iter9_reg <= data_57_V_read_3_reg_8786_pp0_iter8_reg;
        data_58_V_read_3_reg_8756 <= data_58_V_read_int_reg;
        data_58_V_read_3_reg_8756_pp0_iter10_reg <= data_58_V_read_3_reg_8756_pp0_iter9_reg;
        data_58_V_read_3_reg_8756_pp0_iter11_reg <= data_58_V_read_3_reg_8756_pp0_iter10_reg;
        data_58_V_read_3_reg_8756_pp0_iter12_reg <= data_58_V_read_3_reg_8756_pp0_iter11_reg;
        data_58_V_read_3_reg_8756_pp0_iter13_reg <= data_58_V_read_3_reg_8756_pp0_iter12_reg;
        data_58_V_read_3_reg_8756_pp0_iter14_reg <= data_58_V_read_3_reg_8756_pp0_iter13_reg;
        data_58_V_read_3_reg_8756_pp0_iter15_reg <= data_58_V_read_3_reg_8756_pp0_iter14_reg;
        data_58_V_read_3_reg_8756_pp0_iter1_reg <= data_58_V_read_3_reg_8756;
        data_58_V_read_3_reg_8756_pp0_iter2_reg <= data_58_V_read_3_reg_8756_pp0_iter1_reg;
        data_58_V_read_3_reg_8756_pp0_iter3_reg <= data_58_V_read_3_reg_8756_pp0_iter2_reg;
        data_58_V_read_3_reg_8756_pp0_iter4_reg <= data_58_V_read_3_reg_8756_pp0_iter3_reg;
        data_58_V_read_3_reg_8756_pp0_iter5_reg <= data_58_V_read_3_reg_8756_pp0_iter4_reg;
        data_58_V_read_3_reg_8756_pp0_iter6_reg <= data_58_V_read_3_reg_8756_pp0_iter5_reg;
        data_58_V_read_3_reg_8756_pp0_iter7_reg <= data_58_V_read_3_reg_8756_pp0_iter6_reg;
        data_58_V_read_3_reg_8756_pp0_iter8_reg <= data_58_V_read_3_reg_8756_pp0_iter7_reg;
        data_58_V_read_3_reg_8756_pp0_iter9_reg <= data_58_V_read_3_reg_8756_pp0_iter8_reg;
        data_59_V_read_3_reg_8724 <= data_59_V_read_int_reg;
        data_59_V_read_3_reg_8724_pp0_iter10_reg <= data_59_V_read_3_reg_8724_pp0_iter9_reg;
        data_59_V_read_3_reg_8724_pp0_iter11_reg <= data_59_V_read_3_reg_8724_pp0_iter10_reg;
        data_59_V_read_3_reg_8724_pp0_iter12_reg <= data_59_V_read_3_reg_8724_pp0_iter11_reg;
        data_59_V_read_3_reg_8724_pp0_iter13_reg <= data_59_V_read_3_reg_8724_pp0_iter12_reg;
        data_59_V_read_3_reg_8724_pp0_iter14_reg <= data_59_V_read_3_reg_8724_pp0_iter13_reg;
        data_59_V_read_3_reg_8724_pp0_iter15_reg <= data_59_V_read_3_reg_8724_pp0_iter14_reg;
        data_59_V_read_3_reg_8724_pp0_iter16_reg <= data_59_V_read_3_reg_8724_pp0_iter15_reg;
        data_59_V_read_3_reg_8724_pp0_iter1_reg <= data_59_V_read_3_reg_8724;
        data_59_V_read_3_reg_8724_pp0_iter2_reg <= data_59_V_read_3_reg_8724_pp0_iter1_reg;
        data_59_V_read_3_reg_8724_pp0_iter3_reg <= data_59_V_read_3_reg_8724_pp0_iter2_reg;
        data_59_V_read_3_reg_8724_pp0_iter4_reg <= data_59_V_read_3_reg_8724_pp0_iter3_reg;
        data_59_V_read_3_reg_8724_pp0_iter5_reg <= data_59_V_read_3_reg_8724_pp0_iter4_reg;
        data_59_V_read_3_reg_8724_pp0_iter6_reg <= data_59_V_read_3_reg_8724_pp0_iter5_reg;
        data_59_V_read_3_reg_8724_pp0_iter7_reg <= data_59_V_read_3_reg_8724_pp0_iter6_reg;
        data_59_V_read_3_reg_8724_pp0_iter8_reg <= data_59_V_read_3_reg_8724_pp0_iter7_reg;
        data_59_V_read_3_reg_8724_pp0_iter9_reg <= data_59_V_read_3_reg_8724_pp0_iter8_reg;
        data_5_V_read_9_reg_10245 <= data_5_V_read_int_reg;
        data_5_V_read_9_reg_10245_pp0_iter1_reg <= data_5_V_read_9_reg_10245;
        data_5_V_read_9_reg_10245_pp0_iter2_reg <= data_5_V_read_9_reg_10245_pp0_iter1_reg;
        data_5_V_read_9_reg_10245_pp0_iter3_reg <= data_5_V_read_9_reg_10245_pp0_iter2_reg;
        data_60_V_read61_reg_8691 <= data_60_V_read_int_reg;
        data_60_V_read61_reg_8691_pp0_iter10_reg <= data_60_V_read61_reg_8691_pp0_iter9_reg;
        data_60_V_read61_reg_8691_pp0_iter11_reg <= data_60_V_read61_reg_8691_pp0_iter10_reg;
        data_60_V_read61_reg_8691_pp0_iter12_reg <= data_60_V_read61_reg_8691_pp0_iter11_reg;
        data_60_V_read61_reg_8691_pp0_iter13_reg <= data_60_V_read61_reg_8691_pp0_iter12_reg;
        data_60_V_read61_reg_8691_pp0_iter14_reg <= data_60_V_read61_reg_8691_pp0_iter13_reg;
        data_60_V_read61_reg_8691_pp0_iter15_reg <= data_60_V_read61_reg_8691_pp0_iter14_reg;
        data_60_V_read61_reg_8691_pp0_iter16_reg <= data_60_V_read61_reg_8691_pp0_iter15_reg;
        data_60_V_read61_reg_8691_pp0_iter1_reg <= data_60_V_read61_reg_8691;
        data_60_V_read61_reg_8691_pp0_iter2_reg <= data_60_V_read61_reg_8691_pp0_iter1_reg;
        data_60_V_read61_reg_8691_pp0_iter3_reg <= data_60_V_read61_reg_8691_pp0_iter2_reg;
        data_60_V_read61_reg_8691_pp0_iter4_reg <= data_60_V_read61_reg_8691_pp0_iter3_reg;
        data_60_V_read61_reg_8691_pp0_iter5_reg <= data_60_V_read61_reg_8691_pp0_iter4_reg;
        data_60_V_read61_reg_8691_pp0_iter6_reg <= data_60_V_read61_reg_8691_pp0_iter5_reg;
        data_60_V_read61_reg_8691_pp0_iter7_reg <= data_60_V_read61_reg_8691_pp0_iter6_reg;
        data_60_V_read61_reg_8691_pp0_iter8_reg <= data_60_V_read61_reg_8691_pp0_iter7_reg;
        data_60_V_read61_reg_8691_pp0_iter9_reg <= data_60_V_read61_reg_8691_pp0_iter8_reg;
        data_61_V_read62_reg_8663 <= data_61_V_read_int_reg;
        data_61_V_read62_reg_8663_pp0_iter10_reg <= data_61_V_read62_reg_8663_pp0_iter9_reg;
        data_61_V_read62_reg_8663_pp0_iter11_reg <= data_61_V_read62_reg_8663_pp0_iter10_reg;
        data_61_V_read62_reg_8663_pp0_iter12_reg <= data_61_V_read62_reg_8663_pp0_iter11_reg;
        data_61_V_read62_reg_8663_pp0_iter13_reg <= data_61_V_read62_reg_8663_pp0_iter12_reg;
        data_61_V_read62_reg_8663_pp0_iter14_reg <= data_61_V_read62_reg_8663_pp0_iter13_reg;
        data_61_V_read62_reg_8663_pp0_iter15_reg <= data_61_V_read62_reg_8663_pp0_iter14_reg;
        data_61_V_read62_reg_8663_pp0_iter16_reg <= data_61_V_read62_reg_8663_pp0_iter15_reg;
        data_61_V_read62_reg_8663_pp0_iter1_reg <= data_61_V_read62_reg_8663;
        data_61_V_read62_reg_8663_pp0_iter2_reg <= data_61_V_read62_reg_8663_pp0_iter1_reg;
        data_61_V_read62_reg_8663_pp0_iter3_reg <= data_61_V_read62_reg_8663_pp0_iter2_reg;
        data_61_V_read62_reg_8663_pp0_iter4_reg <= data_61_V_read62_reg_8663_pp0_iter3_reg;
        data_61_V_read62_reg_8663_pp0_iter5_reg <= data_61_V_read62_reg_8663_pp0_iter4_reg;
        data_61_V_read62_reg_8663_pp0_iter6_reg <= data_61_V_read62_reg_8663_pp0_iter5_reg;
        data_61_V_read62_reg_8663_pp0_iter7_reg <= data_61_V_read62_reg_8663_pp0_iter6_reg;
        data_61_V_read62_reg_8663_pp0_iter8_reg <= data_61_V_read62_reg_8663_pp0_iter7_reg;
        data_61_V_read62_reg_8663_pp0_iter9_reg <= data_61_V_read62_reg_8663_pp0_iter8_reg;
        data_62_V_read_3_reg_8645 <= data_62_V_read_int_reg;
        data_62_V_read_3_reg_8645_pp0_iter10_reg <= data_62_V_read_3_reg_8645_pp0_iter9_reg;
        data_62_V_read_3_reg_8645_pp0_iter11_reg <= data_62_V_read_3_reg_8645_pp0_iter10_reg;
        data_62_V_read_3_reg_8645_pp0_iter12_reg <= data_62_V_read_3_reg_8645_pp0_iter11_reg;
        data_62_V_read_3_reg_8645_pp0_iter13_reg <= data_62_V_read_3_reg_8645_pp0_iter12_reg;
        data_62_V_read_3_reg_8645_pp0_iter14_reg <= data_62_V_read_3_reg_8645_pp0_iter13_reg;
        data_62_V_read_3_reg_8645_pp0_iter15_reg <= data_62_V_read_3_reg_8645_pp0_iter14_reg;
        data_62_V_read_3_reg_8645_pp0_iter16_reg <= data_62_V_read_3_reg_8645_pp0_iter15_reg;
        data_62_V_read_3_reg_8645_pp0_iter1_reg <= data_62_V_read_3_reg_8645;
        data_62_V_read_3_reg_8645_pp0_iter2_reg <= data_62_V_read_3_reg_8645_pp0_iter1_reg;
        data_62_V_read_3_reg_8645_pp0_iter3_reg <= data_62_V_read_3_reg_8645_pp0_iter2_reg;
        data_62_V_read_3_reg_8645_pp0_iter4_reg <= data_62_V_read_3_reg_8645_pp0_iter3_reg;
        data_62_V_read_3_reg_8645_pp0_iter5_reg <= data_62_V_read_3_reg_8645_pp0_iter4_reg;
        data_62_V_read_3_reg_8645_pp0_iter6_reg <= data_62_V_read_3_reg_8645_pp0_iter5_reg;
        data_62_V_read_3_reg_8645_pp0_iter7_reg <= data_62_V_read_3_reg_8645_pp0_iter6_reg;
        data_62_V_read_3_reg_8645_pp0_iter8_reg <= data_62_V_read_3_reg_8645_pp0_iter7_reg;
        data_62_V_read_3_reg_8645_pp0_iter9_reg <= data_62_V_read_3_reg_8645_pp0_iter8_reg;
        data_63_V_read_3_reg_8620 <= data_63_V_read_int_reg;
        data_63_V_read_3_reg_8620_pp0_iter10_reg <= data_63_V_read_3_reg_8620_pp0_iter9_reg;
        data_63_V_read_3_reg_8620_pp0_iter11_reg <= data_63_V_read_3_reg_8620_pp0_iter10_reg;
        data_63_V_read_3_reg_8620_pp0_iter12_reg <= data_63_V_read_3_reg_8620_pp0_iter11_reg;
        data_63_V_read_3_reg_8620_pp0_iter13_reg <= data_63_V_read_3_reg_8620_pp0_iter12_reg;
        data_63_V_read_3_reg_8620_pp0_iter14_reg <= data_63_V_read_3_reg_8620_pp0_iter13_reg;
        data_63_V_read_3_reg_8620_pp0_iter15_reg <= data_63_V_read_3_reg_8620_pp0_iter14_reg;
        data_63_V_read_3_reg_8620_pp0_iter16_reg <= data_63_V_read_3_reg_8620_pp0_iter15_reg;
        data_63_V_read_3_reg_8620_pp0_iter1_reg <= data_63_V_read_3_reg_8620;
        data_63_V_read_3_reg_8620_pp0_iter2_reg <= data_63_V_read_3_reg_8620_pp0_iter1_reg;
        data_63_V_read_3_reg_8620_pp0_iter3_reg <= data_63_V_read_3_reg_8620_pp0_iter2_reg;
        data_63_V_read_3_reg_8620_pp0_iter4_reg <= data_63_V_read_3_reg_8620_pp0_iter3_reg;
        data_63_V_read_3_reg_8620_pp0_iter5_reg <= data_63_V_read_3_reg_8620_pp0_iter4_reg;
        data_63_V_read_3_reg_8620_pp0_iter6_reg <= data_63_V_read_3_reg_8620_pp0_iter5_reg;
        data_63_V_read_3_reg_8620_pp0_iter7_reg <= data_63_V_read_3_reg_8620_pp0_iter6_reg;
        data_63_V_read_3_reg_8620_pp0_iter8_reg <= data_63_V_read_3_reg_8620_pp0_iter7_reg;
        data_63_V_read_3_reg_8620_pp0_iter9_reg <= data_63_V_read_3_reg_8620_pp0_iter8_reg;
        data_6_V_read_9_reg_10218 <= data_6_V_read_int_reg;
        data_6_V_read_9_reg_10218_pp0_iter1_reg <= data_6_V_read_9_reg_10218;
        data_6_V_read_9_reg_10218_pp0_iter2_reg <= data_6_V_read_9_reg_10218_pp0_iter1_reg;
        data_6_V_read_9_reg_10218_pp0_iter3_reg <= data_6_V_read_9_reg_10218_pp0_iter2_reg;
        data_7_V_read_9_reg_10191 <= data_7_V_read_int_reg;
        data_7_V_read_9_reg_10191_pp0_iter1_reg <= data_7_V_read_9_reg_10191;
        data_7_V_read_9_reg_10191_pp0_iter2_reg <= data_7_V_read_9_reg_10191_pp0_iter1_reg;
        data_7_V_read_9_reg_10191_pp0_iter3_reg <= data_7_V_read_9_reg_10191_pp0_iter2_reg;
        data_7_V_read_9_reg_10191_pp0_iter4_reg <= data_7_V_read_9_reg_10191_pp0_iter3_reg;
        data_8_V_read_8_reg_10164 <= data_8_V_read_int_reg;
        data_8_V_read_8_reg_10164_pp0_iter1_reg <= data_8_V_read_8_reg_10164;
        data_8_V_read_8_reg_10164_pp0_iter2_reg <= data_8_V_read_8_reg_10164_pp0_iter1_reg;
        data_8_V_read_8_reg_10164_pp0_iter3_reg <= data_8_V_read_8_reg_10164_pp0_iter2_reg;
        data_8_V_read_8_reg_10164_pp0_iter4_reg <= data_8_V_read_8_reg_10164_pp0_iter3_reg;
        data_9_V_read_8_reg_10136 <= data_9_V_read_int_reg;
        data_9_V_read_8_reg_10136_pp0_iter1_reg <= data_9_V_read_8_reg_10136;
        data_9_V_read_8_reg_10136_pp0_iter2_reg <= data_9_V_read_8_reg_10136_pp0_iter1_reg;
        data_9_V_read_8_reg_10136_pp0_iter3_reg <= data_9_V_read_8_reg_10136_pp0_iter2_reg;
        data_9_V_read_8_reg_10136_pp0_iter4_reg <= data_9_V_read_8_reg_10136_pp0_iter3_reg;
        sub_ln703_106_reg_10707 <= sub_ln703_106_fu_1378_p2;
        sub_ln703_107_reg_10712 <= sub_ln703_107_fu_1383_p2;
        sub_ln703_108_reg_10717 <= sub_ln703_108_fu_1388_p2;
        sub_ln703_109_reg_10722 <= sub_ln703_109_fu_1407_p2;
        sub_ln703_10_reg_10420 <= sub_ln703_10_fu_615_p2;
        sub_ln703_115_reg_10727 <= sub_ln703_115_fu_1432_p2;
        sub_ln703_11_reg_10398 <= sub_ln703_11_fu_576_p2;
        sub_ln703_11_reg_10398_pp0_iter3_reg <= sub_ln703_11_reg_10398;
        sub_ln703_122_reg_10742 <= sub_ln703_122_fu_1462_p2;
        sub_ln703_123_reg_10747 <= sub_ln703_123_fu_1467_p2;
        sub_ln703_125_reg_10757 <= sub_ln703_125_fu_1482_p2;
        sub_ln703_128_reg_10762 <= sub_ln703_128_fu_1496_p2;
        sub_ln703_133_reg_10782 <= sub_ln703_133_fu_1532_p2;
        sub_ln703_137_reg_10787 <= sub_ln703_137_fu_1548_p2;
        sub_ln703_141_reg_10792 <= sub_ln703_141_fu_1553_p2;
        sub_ln703_142_reg_10797 <= sub_ln703_142_fu_1558_p2;
        sub_ln703_146_reg_10812 <= sub_ln703_146_fu_1580_p2;
        sub_ln703_152_reg_10822 <= sub_ln703_152_fu_1599_p2;
        sub_ln703_154_reg_10832 <= sub_ln703_154_fu_1609_p2;
        sub_ln703_15_reg_10430 <= sub_ln703_15_fu_631_p2;
        sub_ln703_166_reg_10863 <= sub_ln703_166_fu_1834_p2;
        sub_ln703_16_reg_10436 <= sub_ln703_16_fu_640_p2;
        sub_ln703_17_reg_10453 <= sub_ln703_17_fu_653_p2;
        sub_ln703_183_reg_10868 <= sub_ln703_183_fu_1959_p2;
        sub_ln703_184_reg_10878 <= sub_ln703_184_fu_1984_p2;
        sub_ln703_186_reg_10883 <= sub_ln703_186_fu_1994_p2;
        sub_ln703_18_reg_10459 <= sub_ln703_18_fu_658_p2;
        sub_ln703_191_reg_10893 <= sub_ln703_191_fu_2029_p2;
        sub_ln703_194_reg_10908 <= sub_ln703_194_fu_2054_p2;
        sub_ln703_196_reg_10913 <= sub_ln703_196_fu_2074_p2;
        sub_ln703_198_reg_10935 <= sub_ln703_198_fu_2099_p2;
        sub_ln703_1_reg_10348 <= sub_ln703_1_fu_540_p2;
        sub_ln703_200_reg_10950 <= sub_ln703_200_fu_2115_p2;
        sub_ln703_202_reg_10955 <= sub_ln703_202_fu_2120_p2;
        sub_ln703_203_reg_10965 <= sub_ln703_203_fu_2131_p2;
        sub_ln703_204_reg_10975 <= sub_ln703_204_fu_2142_p2;
        sub_ln703_208_reg_10985 <= sub_ln703_208_fu_2152_p2;
        sub_ln703_209_reg_10990 <= sub_ln703_209_fu_2157_p2;
        sub_ln703_20_reg_10465 <= sub_ln703_20_fu_662_p2;
        sub_ln703_210_reg_10995 <= sub_ln703_210_fu_2162_p2;
        sub_ln703_212_reg_11000 <= sub_ln703_212_fu_2173_p2;
        sub_ln703_230_reg_11010 <= sub_ln703_230_fu_2194_p2;
        sub_ln703_234_reg_11046 <= sub_ln703_234_fu_2395_p2;
        sub_ln703_237_reg_11020 <= sub_ln703_237_fu_2214_p2;
        sub_ln703_23_reg_10471 <= sub_ln703_23_fu_666_p2;
        sub_ln703_246_reg_11051 <= sub_ln703_246_fu_2477_p2;
        sub_ln703_249_reg_11056 <= sub_ln703_249_fu_2496_p2;
        sub_ln703_250_reg_11061 <= sub_ln703_250_fu_2501_p2;
        sub_ln703_251_reg_11066 <= sub_ln703_251_fu_2506_p2;
        sub_ln703_254_reg_11076 <= sub_ln703_254_fu_2525_p2;
        sub_ln703_256_reg_11081 <= sub_ln703_256_fu_2534_p2;
        sub_ln703_257_reg_11086 <= sub_ln703_257_fu_2539_p2;
        sub_ln703_261_reg_11091 <= sub_ln703_261_fu_2569_p2;
        sub_ln703_262_reg_11096 <= sub_ln703_262_fu_2574_p2;
        sub_ln703_263_reg_11101 <= sub_ln703_263_fu_2579_p2;
        sub_ln703_265_reg_11116 <= sub_ln703_265_fu_2613_p2;
        sub_ln703_270_reg_11121 <= sub_ln703_270_fu_2628_p2;
        sub_ln703_272_reg_11138 <= sub_ln703_272_fu_2647_p2;
        sub_ln703_274_reg_11143 <= sub_ln703_274_fu_2652_p2;
        sub_ln703_275_reg_11153 <= sub_ln703_275_fu_2662_p2;
        sub_ln703_281_reg_11163 <= sub_ln703_281_fu_2688_p2;
        sub_ln703_284_reg_11168 <= sub_ln703_284_fu_2698_p2;
        sub_ln703_289_reg_11173 <= sub_ln703_289_fu_2703_p2;
        sub_ln703_28_reg_10476 <= sub_ln703_28_fu_671_p2;
        sub_ln703_293_reg_11178 <= sub_ln703_293_fu_2708_p2;
        sub_ln703_296_reg_11183 <= sub_ln703_296_fu_2713_p2;
        sub_ln703_2_reg_10367 <= sub_ln703_2_fu_552_p2;
        sub_ln703_301_reg_11188 <= sub_ln703_301_fu_2718_p2;
        sub_ln703_313_reg_11257 <= sub_ln703_313_fu_2998_p2;
        sub_ln703_315_reg_11267 <= sub_ln703_315_fu_3021_p2;
        sub_ln703_326_reg_11277 <= sub_ln703_326_fu_3101_p2;
        sub_ln703_328_reg_11282 <= sub_ln703_328_fu_3111_p2;
        sub_ln703_333_reg_11292 <= sub_ln703_333_fu_3155_p2;
        sub_ln703_334_reg_11302 <= sub_ln703_334_fu_3175_p2;
        sub_ln703_336_reg_11307 <= sub_ln703_336_fu_3180_p2;
        sub_ln703_339_reg_11317 <= sub_ln703_339_fu_3200_p2;
        sub_ln703_340_reg_11322 <= sub_ln703_340_fu_3205_p2;
        sub_ln703_342_reg_11327 <= sub_ln703_342_fu_3215_p2;
        sub_ln703_344_reg_11332 <= sub_ln703_344_fu_3220_p2;
        sub_ln703_345_reg_11337 <= sub_ln703_345_fu_3234_p2;
        sub_ln703_350_reg_11342 <= sub_ln703_350_fu_3244_p2;
        sub_ln703_353_reg_11352 <= sub_ln703_353_fu_3269_p2;
        sub_ln703_356_reg_11367 <= sub_ln703_356_fu_3290_p2;
        sub_ln703_358_reg_11372 <= sub_ln703_358_fu_3300_p2;
        sub_ln703_362_reg_11377 <= sub_ln703_362_fu_3305_p2;
        sub_ln703_371_reg_11397 <= sub_ln703_371_fu_3324_p2;
        sub_ln703_384_reg_11474 <= sub_ln703_384_fu_3645_p2;
        sub_ln703_386_reg_11484 <= sub_ln703_386_fu_3660_p2;
        sub_ln703_387_reg_11489 <= sub_ln703_387_fu_3665_p2;
        sub_ln703_38_reg_10508 <= sub_ln703_38_fu_814_p2;
        sub_ln703_390_reg_11499 <= sub_ln703_390_fu_3690_p2;
        sub_ln703_393_reg_11504 <= sub_ln703_393_fu_3705_p2;
        sub_ln703_394_reg_11509 <= sub_ln703_394_fu_3710_p2;
        sub_ln703_395_reg_11514 <= sub_ln703_395_fu_3720_p2;
        sub_ln703_399_reg_11524 <= sub_ln703_399_fu_3761_p2;
        sub_ln703_39_reg_10513 <= sub_ln703_39_fu_819_p2;
        sub_ln703_3_reg_10379 <= sub_ln703_3_fu_560_p2;
        sub_ln703_401_reg_11529 <= sub_ln703_401_fu_3781_p2;
        sub_ln703_402_reg_11534 <= sub_ln703_402_fu_3786_p2;
        sub_ln703_403_reg_11539 <= sub_ln703_403_fu_3791_p2;
        sub_ln703_405_reg_11554 <= sub_ln703_405_fu_3816_p2;
        sub_ln703_408_reg_11564 <= sub_ln703_408_fu_3845_p2;
        sub_ln703_40_reg_10519 <= sub_ln703_40_fu_824_p2;
        sub_ln703_411_reg_11569 <= sub_ln703_411_fu_3850_p2;
        sub_ln703_412_reg_11574 <= sub_ln703_412_fu_3855_p2;
        sub_ln703_414_reg_11579 <= sub_ln703_414_fu_3860_p2;
        sub_ln703_416_reg_11584 <= sub_ln703_416_fu_3865_p2;
        sub_ln703_419_reg_11594 <= sub_ln703_419_fu_3884_p2;
        sub_ln703_43_reg_10524 <= sub_ln703_43_fu_838_p2;
        sub_ln703_440_reg_11624 <= sub_ln703_440_fu_3938_p2;
        sub_ln703_448_reg_11673 <= sub_ln703_448_fu_4206_p2;
        sub_ln703_452_reg_11678 <= sub_ln703_452_fu_4231_p2;
        sub_ln703_453_reg_11683 <= sub_ln703_453_fu_4236_p2;
        sub_ln703_458_reg_11688 <= sub_ln703_458_fu_4270_p2;
        sub_ln703_461_reg_11693 <= sub_ln703_461_fu_4303_p2;
        sub_ln703_462_reg_11703 <= sub_ln703_462_fu_4313_p2;
        sub_ln703_467_reg_11713 <= sub_ln703_467_fu_4333_p2;
        sub_ln703_468_reg_11718 <= sub_ln703_468_fu_4353_p2;
        sub_ln703_469_reg_11733 <= sub_ln703_469_fu_4368_p2;
        sub_ln703_470_reg_11738 <= sub_ln703_470_fu_4373_p2;
        sub_ln703_475_reg_11753 <= sub_ln703_475_fu_4418_p2;
        sub_ln703_482_reg_11773 <= sub_ln703_482_fu_4447_p2;
        sub_ln703_483_reg_11778 <= sub_ln703_483_fu_4452_p2;
        sub_ln703_488_reg_11783 <= sub_ln703_488_fu_4457_p2;
        sub_ln703_490_reg_11788 <= sub_ln703_490_fu_4462_p2;
        sub_ln703_491_reg_11793 <= sub_ln703_491_fu_4467_p2;
        sub_ln703_4_reg_10361 <= sub_ln703_4_fu_548_p2;
        sub_ln703_4_reg_10361_pp0_iter2_reg <= sub_ln703_4_reg_10361;
        sub_ln703_503_reg_11813 <= sub_ln703_503_fu_4516_p2;
        sub_ln703_505_reg_11818 <= sub_ln703_505_fu_4521_p2;
        sub_ln703_526_reg_11864 <= sub_ln703_526_fu_4860_p2;
        sub_ln703_527_reg_11869 <= sub_ln703_527_fu_4865_p2;
        sub_ln703_529_reg_11879 <= sub_ln703_529_fu_4880_p2;
        sub_ln703_532_reg_11884 <= sub_ln703_532_fu_4894_p2;
        sub_ln703_533_reg_11894 <= sub_ln703_533_fu_4904_p2;
        sub_ln703_535_reg_11899 <= sub_ln703_535_fu_4919_p2;
        sub_ln703_538_reg_11904 <= sub_ln703_538_fu_4934_p2;
        sub_ln703_539_reg_11909 <= sub_ln703_539_fu_4939_p2;
        sub_ln703_53_reg_10534 <= sub_ln703_53_fu_912_p2;
        sub_ln703_540_reg_11914 <= sub_ln703_540_fu_4944_p2;
        sub_ln703_541_reg_11919 <= sub_ln703_541_fu_4949_p2;
        sub_ln703_542_reg_11924 <= sub_ln703_542_fu_4954_p2;
        sub_ln703_544_reg_11934 <= sub_ln703_544_fu_4984_p2;
        sub_ln703_551_reg_11949 <= sub_ln703_551_fu_5004_p2;
        sub_ln703_556_reg_11964 <= sub_ln703_556_fu_5024_p2;
        sub_ln703_557_reg_11969 <= sub_ln703_557_fu_5029_p2;
        sub_ln703_558_reg_11974 <= sub_ln703_558_fu_5034_p2;
        sub_ln703_573_reg_12007 <= sub_ln703_573_fu_5101_p2;
        sub_ln703_582_reg_12012 <= sub_ln703_582_fu_5106_p2;
        sub_ln703_583_reg_12017 <= sub_ln703_583_fu_5111_p2;
        sub_ln703_586_reg_12061 <= sub_ln703_586_fu_5351_p2;
        sub_ln703_589_reg_12066 <= sub_ln703_589_fu_5375_p2;
        sub_ln703_58_reg_10545 <= sub_ln703_58_fu_922_p2;
        sub_ln703_593_reg_12071 <= sub_ln703_593_fu_5410_p2;
        sub_ln703_594_reg_12076 <= sub_ln703_594_fu_5415_p2;
        sub_ln703_595_reg_12081 <= sub_ln703_595_fu_5420_p2;
        sub_ln703_598_reg_12091 <= sub_ln703_598_fu_5454_p2;
        sub_ln703_603_reg_12101 <= sub_ln703_603_fu_5491_p2;
        sub_ln703_604_reg_12106 <= sub_ln703_604_fu_5496_p2;
        sub_ln703_605_reg_12111 <= sub_ln703_605_fu_5501_p2;
        sub_ln703_608_reg_12116 <= sub_ln703_608_fu_5511_p2;
        sub_ln703_609_reg_12121 <= sub_ln703_609_fu_5516_p2;
        sub_ln703_610_reg_12126 <= sub_ln703_610_fu_5521_p2;
        sub_ln703_612_reg_12131 <= sub_ln703_612_fu_5526_p2;
        sub_ln703_613_reg_12136 <= sub_ln703_613_fu_5531_p2;
        sub_ln703_614_reg_12141 <= sub_ln703_614_fu_5536_p2;
        sub_ln703_618_reg_12156 <= sub_ln703_618_fu_5566_p2;
        sub_ln703_624_reg_12166 <= sub_ln703_624_fu_5596_p2;
        sub_ln703_62_reg_10550 <= sub_ln703_62_fu_942_p2;
        sub_ln703_630_reg_12171 <= sub_ln703_630_fu_5627_p2;
        sub_ln703_631_reg_12176 <= sub_ln703_631_fu_5632_p2;
        sub_ln703_634_reg_12181 <= sub_ln703_634_fu_5637_p2;
        sub_ln703_637_reg_12186 <= sub_ln703_637_fu_5642_p2;
        sub_ln703_638_reg_12191 <= sub_ln703_638_fu_5647_p2;
        sub_ln703_63_reg_10555 <= sub_ln703_63_fu_947_p2;
        sub_ln703_644_reg_12204 <= sub_ln703_644_fu_5656_p2;
        sub_ln703_648_reg_12209 <= sub_ln703_648_fu_5661_p2;
        sub_ln703_64_reg_10560 <= sub_ln703_64_fu_957_p2;
        sub_ln703_650_reg_12214 <= sub_ln703_650_fu_5666_p2;
        sub_ln703_662_reg_12248 <= sub_ln703_662_fu_5918_p2;
        sub_ln703_665_reg_12253 <= sub_ln703_665_fu_5932_p2;
        sub_ln703_667_reg_12263 <= sub_ln703_667_fu_5956_p2;
        sub_ln703_669_reg_12268 <= sub_ln703_669_fu_5975_p2;
        sub_ln703_66_reg_10581 <= sub_ln703_66_fu_987_p2;
        sub_ln703_676_reg_12278 <= sub_ln703_676_fu_6033_p2;
        sub_ln703_678_reg_12283 <= sub_ln703_678_fu_6052_p2;
        sub_ln703_679_reg_12288 <= sub_ln703_679_fu_6057_p2;
        sub_ln703_680_reg_12293 <= sub_ln703_680_fu_6062_p2;
        sub_ln703_682_reg_12298 <= sub_ln703_682_fu_6067_p2;
        sub_ln703_684_reg_12303 <= sub_ln703_684_fu_6072_p2;
        sub_ln703_686_reg_12308 <= sub_ln703_686_fu_6077_p2;
        sub_ln703_687_reg_12313 <= sub_ln703_687_fu_6086_p2;
        sub_ln703_688_reg_12318 <= sub_ln703_688_fu_6091_p2;
        sub_ln703_690_reg_12323 <= sub_ln703_690_fu_6101_p2;
        sub_ln703_691_reg_12328 <= sub_ln703_691_fu_6106_p2;
        sub_ln703_692_reg_12333 <= sub_ln703_692_fu_6111_p2;
        sub_ln703_693_reg_12338 <= sub_ln703_693_fu_6116_p2;
        sub_ln703_694_reg_12343 <= sub_ln703_694_fu_6126_p2;
        sub_ln703_696_reg_12353 <= sub_ln703_696_fu_6136_p2;
        sub_ln703_697_reg_12358 <= sub_ln703_697_fu_6141_p2;
        sub_ln703_6_reg_10408 <= sub_ln703_6_fu_595_p2;
        sub_ln703_700_reg_12378 <= sub_ln703_700_fu_6172_p2;
        sub_ln703_704_reg_12383 <= sub_ln703_704_fu_6177_p2;
        sub_ln703_707_reg_12388 <= sub_ln703_707_fu_6182_p2;
        sub_ln703_70_reg_10586 <= sub_ln703_70_fu_992_p2;
        sub_ln703_71_reg_10596 <= sub_ln703_71_fu_1002_p2;
        sub_ln703_724_reg_12450 <= sub_ln703_724_fu_6432_p2;
        sub_ln703_727_reg_12460 <= sub_ln703_727_fu_6452_p2;
        sub_ln703_728_reg_12465 <= sub_ln703_728_fu_6457_p2;
        sub_ln703_733_reg_12470 <= sub_ln703_733_fu_6487_p2;
        sub_ln703_736_reg_12475 <= sub_ln703_736_fu_6502_p2;
        sub_ln703_73_reg_10611 <= sub_ln703_73_fu_1026_p2;
        sub_ln703_746_reg_12500 <= sub_ln703_746_fu_6579_p2;
        sub_ln703_749_reg_12510 <= sub_ln703_749_fu_6599_p2;
        sub_ln703_757_reg_12515 <= sub_ln703_757_fu_6629_p2;
        sub_ln703_759_reg_12525 <= sub_ln703_759_fu_6639_p2;
        sub_ln703_75_reg_10616 <= sub_ln703_75_fu_1031_p2;
        sub_ln703_761_reg_12530 <= sub_ln703_761_fu_6644_p2;
        sub_ln703_763_reg_12540 <= sub_ln703_763_fu_6654_p2;
        sub_ln703_767_reg_12545 <= sub_ln703_767_fu_6659_p2;
        sub_ln703_769_reg_12555 <= sub_ln703_769_fu_6684_p2;
        sub_ln703_770_reg_12570 <= sub_ln703_770_fu_6708_p2;
        sub_ln703_781_reg_12580 <= sub_ln703_781_fu_6739_p2;
        sub_ln703_787_reg_12590 <= sub_ln703_787_fu_6759_p2;
        sub_ln703_797_reg_12645 <= sub_ln703_797_fu_7030_p2;
        sub_ln703_799_reg_12595 <= sub_ln703_799_fu_6764_p2;
        sub_ln703_801_reg_12660 <= sub_ln703_801_fu_7060_p2;
        sub_ln703_802_reg_12665 <= sub_ln703_802_fu_7065_p2;
        sub_ln703_805_reg_12670 <= sub_ln703_805_fu_7079_p2;
        sub_ln703_807_reg_12685 <= sub_ln703_807_fu_7099_p2;
        sub_ln703_808_reg_12700 <= sub_ln703_808_fu_7137_p2;
        sub_ln703_814_reg_12735 <= sub_ln703_814_fu_7200_p2;
        sub_ln703_816_reg_12740 <= sub_ln703_816_fu_7205_p2;
        sub_ln703_818_reg_12745 <= sub_ln703_818_fu_7210_p2;
        sub_ln703_820_reg_12750 <= sub_ln703_820_fu_7215_p2;
        sub_ln703_821_reg_12755 <= sub_ln703_821_fu_7220_p2;
        sub_ln703_823_reg_12760 <= sub_ln703_823_fu_7225_p2;
        sub_ln703_824_reg_12765 <= sub_ln703_824_fu_7230_p2;
        sub_ln703_825_reg_12770 <= sub_ln703_825_fu_7235_p2;
        sub_ln703_852_reg_12790 <= sub_ln703_852_fu_7319_p2;
        sub_ln703_857_reg_12835 <= sub_ln703_857_fu_7600_p2;
        sub_ln703_858_reg_12840 <= sub_ln703_858_fu_7605_p2;
        sub_ln703_859_reg_12850 <= sub_ln703_859_fu_7615_p2;
        sub_ln703_862_reg_12795 <= sub_ln703_862_fu_7324_p2;
        sub_ln703_863_reg_12860 <= sub_ln703_863_fu_7639_p2;
        sub_ln703_865_reg_12865 <= sub_ln703_865_fu_7649_p2;
        sub_ln703_866_reg_12870 <= sub_ln703_866_fu_7654_p2;
        sub_ln703_867_reg_12880 <= sub_ln703_867_fu_7669_p2;
        sub_ln703_868_reg_12885 <= sub_ln703_868_fu_7674_p2;
        sub_ln703_869_reg_12800 <= sub_ln703_869_fu_7329_p2;
        sub_ln703_869_reg_12800_pp0_iter16_reg <= sub_ln703_869_reg_12800;
        sub_ln703_870_reg_12895 <= sub_ln703_870_fu_7685_p2;
        sub_ln703_873_reg_12900 <= sub_ln703_873_fu_7710_p2;
        sub_ln703_875_reg_12910 <= sub_ln703_875_fu_7730_p2;
        sub_ln703_879_reg_12915 <= sub_ln703_879_fu_7735_p2;
        sub_ln703_880_reg_12920 <= sub_ln703_880_fu_7750_p2;
        sub_ln703_881_reg_12925 <= sub_ln703_881_fu_7755_p2;
        sub_ln703_892_reg_12935 <= sub_ln703_892_fu_7780_p2;
        sub_ln703_893_reg_12940 <= sub_ln703_893_fu_7785_p2;
        sub_ln703_894_reg_12945 <= sub_ln703_894_fu_7790_p2;
        sub_ln703_895_reg_12950 <= sub_ln703_895_fu_7795_p2;
        sub_ln703_898_reg_12955 <= sub_ln703_898_fu_7805_p2;
        sub_ln703_8_reg_10392 <= sub_ln703_8_fu_572_p2;
        sub_ln703_904_reg_12960 <= sub_ln703_904_fu_7810_p2;
        sub_ln703_911_reg_12970 <= sub_ln703_911_fu_7833_p2;
        sub_ln703_917_reg_12975 <= sub_ln703_917_fu_7838_p2;
        sub_ln703_922_reg_12980 <= sub_ln703_922_fu_7843_p2;
        sub_ln703_92_reg_10636 <= sub_ln703_92_fu_1054_p2;
        sub_ln703_96_reg_10677 <= sub_ln703_96_fu_1294_p2;
        sub_ln703_98_reg_10697 <= sub_ln703_98_fu_1319_p2;
        sub_ln703_reg_10342 <= sub_ln703_fu_536_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_ce_reg)) begin
        ap_return_0_int_reg <= add_ln703_986_fu_8255_p2;
        ap_return_10_int_reg <= acc_10_V_fu_8310_p2;
        ap_return_11_int_reg <= acc_11_V_fu_8315_p2;
        ap_return_12_int_reg <= acc_12_V_fu_8320_p2;
        ap_return_13_int_reg <= acc_13_V_fu_8330_p2;
        ap_return_14_int_reg <= acc_14_V_fu_8335_p2;
        ap_return_15_int_reg <= acc_15_V_fu_8340_p2;
        ap_return_16_int_reg <= acc_16_V_fu_8345_p2;
        ap_return_17_int_reg <= acc_17_V_fu_8350_p2;
        ap_return_18_int_reg <= acc_18_V_fu_8355_p2;
        ap_return_19_int_reg <= acc_19_V_fu_8360_p2;
        ap_return_1_int_reg <= acc_1_V_fu_8265_p2;
        ap_return_20_int_reg <= acc_20_V_fu_8365_p2;
        ap_return_21_int_reg <= acc_21_V_reg_12991;
        ap_return_22_int_reg <= acc_22_V_fu_8370_p2;
        ap_return_23_int_reg <= acc_23_V_fu_8375_p2;
        ap_return_24_int_reg <= acc_24_V_fu_8380_p2;
        ap_return_25_int_reg <= acc_25_V_fu_8385_p2;
        ap_return_26_int_reg <= acc_26_V_fu_8390_p2;
        ap_return_27_int_reg <= acc_27_V_fu_8400_p2;
        ap_return_28_int_reg <= acc_28_V_fu_8405_p2;
        ap_return_29_int_reg <= acc_29_V_fu_8414_p2;
        ap_return_2_int_reg <= acc_2_V_fu_8270_p2;
        ap_return_30_int_reg <= acc_30_V_fu_8419_p2;
        ap_return_31_int_reg <= acc_31_V_fu_8424_p2;
        ap_return_3_int_reg <= acc_3_V_fu_8275_p2;
        ap_return_4_int_reg <= acc_4_V_fu_8280_p2;
        ap_return_5_int_reg <= acc_5_V_fu_8285_p2;
        ap_return_6_int_reg <= acc_6_V_fu_8290_p2;
        ap_return_7_int_reg <= acc_7_V_fu_8295_p2;
        ap_return_8_int_reg <= acc_8_V_fu_8300_p2;
        ap_return_9_int_reg <= acc_9_V_fu_8305_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_ce)) begin
        data_0_V_read_int_reg <= data_0_V_read;
        data_10_V_read_int_reg <= data_10_V_read;
        data_11_V_read_int_reg <= data_11_V_read;
        data_12_V_read_int_reg <= data_12_V_read;
        data_13_V_read_int_reg <= data_13_V_read;
        data_14_V_read_int_reg <= data_14_V_read;
        data_15_V_read_int_reg <= data_15_V_read;
        data_16_V_read_int_reg <= data_16_V_read;
        data_17_V_read_int_reg <= data_17_V_read;
        data_18_V_read_int_reg <= data_18_V_read;
        data_19_V_read_int_reg <= data_19_V_read;
        data_1_V_read_int_reg <= data_1_V_read;
        data_20_V_read_int_reg <= data_20_V_read;
        data_21_V_read_int_reg <= data_21_V_read;
        data_22_V_read_int_reg <= data_22_V_read;
        data_23_V_read_int_reg <= data_23_V_read;
        data_24_V_read_int_reg <= data_24_V_read;
        data_25_V_read_int_reg <= data_25_V_read;
        data_26_V_read_int_reg <= data_26_V_read;
        data_27_V_read_int_reg <= data_27_V_read;
        data_28_V_read_int_reg <= data_28_V_read;
        data_29_V_read_int_reg <= data_29_V_read;
        data_2_V_read_int_reg <= data_2_V_read;
        data_30_V_read_int_reg <= data_30_V_read;
        data_31_V_read_int_reg <= data_31_V_read;
        data_32_V_read_int_reg <= data_32_V_read;
        data_33_V_read_int_reg <= data_33_V_read;
        data_34_V_read_int_reg <= data_34_V_read;
        data_35_V_read_int_reg <= data_35_V_read;
        data_36_V_read_int_reg <= data_36_V_read;
        data_37_V_read_int_reg <= data_37_V_read;
        data_38_V_read_int_reg <= data_38_V_read;
        data_39_V_read_int_reg <= data_39_V_read;
        data_3_V_read_int_reg <= data_3_V_read;
        data_40_V_read_int_reg <= data_40_V_read;
        data_41_V_read_int_reg <= data_41_V_read;
        data_42_V_read_int_reg <= data_42_V_read;
        data_43_V_read_int_reg <= data_43_V_read;
        data_44_V_read_int_reg <= data_44_V_read;
        data_45_V_read_int_reg <= data_45_V_read;
        data_46_V_read_int_reg <= data_46_V_read;
        data_47_V_read_int_reg <= data_47_V_read;
        data_48_V_read_int_reg <= data_48_V_read;
        data_49_V_read_int_reg <= data_49_V_read;
        data_4_V_read_int_reg <= data_4_V_read;
        data_50_V_read_int_reg <= data_50_V_read;
        data_51_V_read_int_reg <= data_51_V_read;
        data_52_V_read_int_reg <= data_52_V_read;
        data_53_V_read_int_reg <= data_53_V_read;
        data_54_V_read_int_reg <= data_54_V_read;
        data_55_V_read_int_reg <= data_55_V_read;
        data_56_V_read_int_reg <= data_56_V_read;
        data_57_V_read_int_reg <= data_57_V_read;
        data_58_V_read_int_reg <= data_58_V_read;
        data_59_V_read_int_reg <= data_59_V_read;
        data_5_V_read_int_reg <= data_5_V_read;
        data_60_V_read_int_reg <= data_60_V_read;
        data_61_V_read_int_reg <= data_61_V_read;
        data_62_V_read_int_reg <= data_62_V_read;
        data_63_V_read_int_reg <= data_63_V_read;
        data_6_V_read_int_reg <= data_6_V_read;
        data_7_V_read_int_reg <= data_7_V_read;
        data_8_V_read_int_reg <= data_8_V_read;
        data_9_V_read_int_reg <= data_9_V_read;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_0 = ap_return_0_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_0 = add_ln703_986_fu_8255_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_1 = ap_return_1_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_1 = acc_1_V_fu_8265_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_10 = ap_return_10_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_10 = acc_10_V_fu_8310_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_11 = ap_return_11_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_11 = acc_11_V_fu_8315_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_12 = ap_return_12_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_12 = acc_12_V_fu_8320_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_13 = ap_return_13_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_13 = acc_13_V_fu_8330_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_14 = ap_return_14_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_14 = acc_14_V_fu_8335_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_15 = ap_return_15_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_15 = acc_15_V_fu_8340_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_16 = ap_return_16_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_16 = acc_16_V_fu_8345_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_17 = ap_return_17_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_17 = acc_17_V_fu_8350_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_18 = ap_return_18_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_18 = acc_18_V_fu_8355_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_19 = ap_return_19_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_19 = acc_19_V_fu_8360_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_2 = ap_return_2_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_2 = acc_2_V_fu_8270_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_20 = ap_return_20_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_20 = acc_20_V_fu_8365_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_21 = ap_return_21_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_21 = acc_21_V_reg_12991;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_22 = ap_return_22_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_22 = acc_22_V_fu_8370_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_23 = ap_return_23_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_23 = acc_23_V_fu_8375_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_24 = ap_return_24_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_24 = acc_24_V_fu_8380_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_25 = ap_return_25_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_25 = acc_25_V_fu_8385_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_26 = ap_return_26_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_26 = acc_26_V_fu_8390_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_27 = ap_return_27_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_27 = acc_27_V_fu_8400_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_28 = ap_return_28_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_28 = acc_28_V_fu_8405_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_29 = ap_return_29_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_29 = acc_29_V_fu_8414_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_3 = ap_return_3_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_3 = acc_3_V_fu_8275_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_30 = ap_return_30_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_30 = acc_30_V_fu_8419_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_31 = ap_return_31_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_31 = acc_31_V_fu_8424_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_4 = ap_return_4_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_4 = acc_4_V_fu_8280_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_5 = ap_return_5_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_5 = acc_5_V_fu_8285_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_6 = ap_return_6_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_6 = acc_6_V_fu_8290_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_7 = ap_return_7_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_7 = acc_7_V_fu_8295_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_8 = ap_return_8_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_8 = acc_8_V_fu_8300_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_9 = ap_return_9_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_9 = acc_9_V_fu_8305_p2;
    end
end

assign acc_10_V_fu_8310_p2 = (add_ln703_974_fu_8159_p2 - data_63_V_read_3_reg_8620_pp0_iter16_reg);

assign acc_11_V_fu_8315_p2 = (sub_ln703_934_fu_8165_p2 - data_63_V_read_3_reg_8620_pp0_iter16_reg);

assign acc_12_V_fu_8320_p2 = (add_ln703_976_fu_8175_p2 - data_63_V_read_3_reg_8620_pp0_iter16_reg);

assign acc_13_V_fu_8330_p2 = (add_ln703_985_reg_12819_pp0_iter16_reg + add_ln703_994_fu_8325_p2);

assign acc_14_V_fu_8335_p2 = (sub_ln703_935_fu_8181_p2 + data_63_V_read_3_reg_8620_pp0_iter16_reg);

assign acc_15_V_fu_8340_p2 = (add_ln703_978_fu_8191_p2 - data_63_V_read_3_reg_8620_pp0_iter16_reg);

assign acc_16_V_fu_8345_p2 = (add_ln703_979_fu_8197_p2 - data_63_V_read_3_reg_8620_pp0_iter16_reg);

assign acc_17_V_fu_8350_p2 = (add_ln703_985_reg_12819_pp0_iter16_reg + sub_ln703_924_fu_8072_p2);

assign acc_18_V_fu_8355_p2 = (add_ln703_985_reg_12819_pp0_iter16_reg + sub_ln703_925_fu_8076_p2);

assign acc_19_V_fu_8360_p2 = (add_ln703_985_reg_12819_pp0_iter16_reg + sub_ln703_926_fu_8080_p2);

assign acc_1_V_fu_8265_p2 = (add_ln703_985_reg_12819_pp0_iter16_reg + add_ln703_987_fu_8260_p2);

assign acc_20_V_fu_8365_p2 = (add_ln703_980_fu_8203_p2 - data_63_V_read_3_reg_8620_pp0_iter16_reg);

assign acc_21_V_fu_7872_p2 = (add_ln703_1003_fu_7867_p2 + add_ln703_1001_fu_7857_p2);

assign acc_22_V_fu_8370_p2 = (add_ln703_985_reg_12819_pp0_iter16_reg + sub_ln703_927_fu_8085_p2);

assign acc_23_V_fu_8375_p2 = (sub_ln703_936_fu_8209_p2 + data_63_V_read_3_reg_8620_pp0_iter16_reg);

assign acc_24_V_fu_8380_p2 = (add_ln703_981_fu_8214_p2 - data_63_V_read_3_reg_8620_pp0_iter16_reg);

assign acc_25_V_fu_8385_p2 = (sub_ln703_937_fu_8219_p2 - data_63_V_read_3_reg_8620_pp0_iter16_reg);

assign acc_26_V_fu_8390_p2 = (sub_ln703_938_fu_8224_p2 - data_63_V_read_3_reg_8620_pp0_iter16_reg);

assign acc_27_V_fu_8400_p2 = (add_ln703_985_reg_12819_pp0_iter16_reg + add_ln703_1007_fu_8395_p2);

assign acc_28_V_fu_8405_p2 = (sub_ln703_939_fu_8229_p2 - data_63_V_read_3_reg_8620_pp0_iter16_reg);

assign acc_29_V_fu_8414_p2 = (add_ln703_985_reg_12819_pp0_iter16_reg + add_ln703_1009_fu_8410_p2);

assign acc_2_V_fu_8270_p2 = (add_ln703_985_reg_12819_pp0_iter16_reg + sub_ln703_919_fu_8037_p2);

assign acc_30_V_fu_8419_p2 = (sub_ln703_940_fu_8234_p2 - data_63_V_read_3_reg_8620_pp0_iter16_reg);

assign acc_31_V_fu_8424_p2 = (add_ln703_983_fu_8244_p2 - data_63_V_read_3_reg_8620_pp0_iter16_reg);

assign acc_3_V_fu_8275_p2 = (add_ln703_985_reg_12819_pp0_iter16_reg + sub_ln703_920_fu_8042_p2);

assign acc_4_V_fu_8280_p2 = (sub_ln703_930_fu_8120_p2 + data_63_V_read_3_reg_8620_pp0_iter16_reg);

assign acc_5_V_fu_8285_p2 = (add_ln703_971_fu_8129_p2 - data_63_V_read_3_reg_8620_pp0_iter16_reg);

assign acc_6_V_fu_8290_p2 = (sub_ln703_931_fu_8134_p2 - data_63_V_read_3_reg_8620_pp0_iter16_reg);

assign acc_7_V_fu_8295_p2 = (sub_ln703_932_fu_8139_p2 + data_63_V_read_3_reg_8620_pp0_iter16_reg);

assign acc_8_V_fu_8300_p2 = (sub_ln703_933_fu_8143_p2 + data_63_V_read_3_reg_8620_pp0_iter16_reg);

assign acc_9_V_fu_8305_p2 = (add_ln703_973_fu_8153_p2 - data_63_V_read_3_reg_8620_pp0_iter16_reg);

assign add_ln703_1000_fu_7852_p2 = (sub_ln703_819_fu_7386_p2 + data_56_V_read_3_reg_8814_pp0_iter15_reg);

assign add_ln703_1001_fu_7857_p2 = (add_ln703_937_fu_7659_p2 + add_ln703_1000_fu_7852_p2);

assign add_ln703_1002_fu_7863_p2 = (add_ln703_985_reg_12819 + data_61_V_read62_reg_8663_pp0_iter15_reg);

assign add_ln703_1003_fu_7867_p2 = (add_ln703_1002_fu_7863_p2 + add_ln703_954_reg_12812);

assign add_ln703_1007_fu_8395_p2 = (sub_ln703_916_fu_8028_p2 + data_61_V_read62_reg_8663_pp0_iter16_reg);

assign add_ln703_1009_fu_8410_p2 = (sub_ln703_917_reg_12975 + data_61_V_read62_reg_8663_pp0_iter16_reg);

assign add_ln703_130_fu_556_p2 = (sub_ln703_1_reg_10348 + data_2_V_read_10_reg_10312_pp0_iter1_reg);

assign add_ln703_131_fu_544_p2 = (add_ln703_reg_10335 + data_2_V_read_10_reg_10312);

assign add_ln703_132_fu_599_p2 = (add_ln703_130_reg_10373 + data_3_V_read_10_reg_10295_pp0_iter2_reg);

assign add_ln703_133_fu_603_p2 = (sub_ln703_3_reg_10379 + data_3_V_read_10_reg_10295_pp0_iter2_reg);

assign add_ln703_134_fu_568_p2 = (add_ln703_131_reg_10354 + data_3_V_read_10_reg_10295_pp0_iter1_reg);

assign add_ln703_135_fu_619_p2 = (sub_ln703_2_reg_10367 + data_3_V_read_10_reg_10295_pp0_iter2_reg);

assign add_ln703_136_fu_623_p2 = (sub_ln703_4_reg_10361_pp0_iter2_reg + data_3_V_read_10_reg_10295_pp0_iter2_reg);

assign add_ln703_137_fu_697_p2 = (sub_ln703_6_reg_10408 + data_4_V_read_10_reg_10273_pp0_iter3_reg);

assign add_ln703_138_fu_701_p2 = (add_ln703_132_reg_10414 + data_4_V_read_10_reg_10273_pp0_iter3_reg);

assign add_ln703_139_fu_636_p2 = (add_ln703_134_reg_10385 + data_4_V_read_10_reg_10273_pp0_iter2_reg);

assign add_ln703_140_fu_644_p2 = (sub_ln703_7_fu_607_p2 + data_4_V_read_10_reg_10273_pp0_iter2_reg);

assign add_ln703_141_fu_649_p2 = (sub_ln703_8_reg_10392 + data_4_V_read_10_reg_10273_pp0_iter2_reg);

assign add_ln703_142_fu_581_p2 = (sub_ln703_reg_10342 + data_2_V_read_10_reg_10312_pp0_iter1_reg);

assign add_ln703_143_fu_585_p2 = (data_3_V_read_10_reg_10295_pp0_iter1_reg + data_4_V_read_10_reg_10273_pp0_iter1_reg);

assign add_ln703_144_fu_589_p2 = (add_ln703_143_fu_585_p2 + add_ln703_142_fu_581_p2);

assign add_ln703_145_fu_736_p2 = (add_ln703_138_fu_701_p2 + data_5_V_read_9_reg_10245_pp0_iter3_reg);

assign add_ln703_146_fu_741_p2 = (sub_ln703_15_reg_10430 + data_5_V_read_9_reg_10245_pp0_iter3_reg);

assign add_ln703_147_fu_745_p2 = (sub_ln703_16_reg_10436 + data_5_V_read_9_reg_10245_pp0_iter3_reg);

assign add_ln703_148_fu_757_p2 = (add_ln703_141_reg_10447 + data_5_V_read_9_reg_10245_pp0_iter3_reg);

assign add_ln703_149_fu_773_p2 = (sub_ln703_19_fu_705_p2 + data_5_V_read_9_reg_10245_pp0_iter3_reg);

assign add_ln703_150_fu_782_p2 = (sub_ln703_22_fu_713_p2 + data_5_V_read_9_reg_10245_pp0_iter3_reg);

assign add_ln703_151_fu_791_p2 = (sub_ln703_20_reg_10465 + data_5_V_read_9_reg_10245_pp0_iter3_reg);

assign add_ln703_152_fu_804_p2 = (sub_ln703_24_fu_717_p2 + data_6_V_read_9_reg_10218_pp0_iter3_reg);

assign add_ln703_153_fu_809_p2 = (sub_ln703_25_fu_722_p2 + data_6_V_read_9_reg_10218_pp0_iter3_reg);

assign add_ln703_154_fu_843_p2 = (sub_ln703_30_fu_753_p2 + data_6_V_read_9_reg_10218_pp0_iter3_reg);

assign add_ln703_155_fu_868_p2 = (data_5_V_read_9_reg_10245_pp0_iter3_reg + data_6_V_read_9_reg_10218_pp0_iter3_reg);

assign add_ln703_156_fu_872_p2 = (add_ln703_155_fu_868_p2 + sub_ln703_18_reg_10459);

assign add_ln703_157_fu_892_p2 = (sub_ln703_35_fu_787_p2 + data_6_V_read_9_reg_10218_pp0_iter3_reg);

assign add_ln703_158_fu_676_p2 = (sub_ln703_12_fu_627_p2 + data_4_V_read_10_reg_10273_pp0_iter2_reg);

assign add_ln703_160_fu_902_p2 = (add_ln703_155_fu_868_p2 + add_ln703_158_reg_10482);

assign add_ln703_161_fu_681_p2 = (data_6_V_read_9_reg_10218_pp0_iter2_reg + data_7_V_read_9_reg_10191_pp0_iter2_reg);

assign add_ln703_162_fu_917_p2 = (add_ln703_161_reg_10487 + sub_ln703_26_fu_727_p2);

assign add_ln703_163_fu_1098_p2 = (sub_ln703_39_reg_10513 + data_7_V_read_9_reg_10191_pp0_iter4_reg);

assign add_ln703_164_fu_937_p2 = (sub_ln703_45_fu_853_p2 + data_7_V_read_9_reg_10191_pp0_iter3_reg);

assign add_ln703_165_fu_952_p2 = (sub_ln703_38_fu_814_p2 + data_7_V_read_9_reg_10191_pp0_iter3_reg);

assign add_ln703_166_fu_962_p2 = (sub_ln703_21_fu_709_p2 + data_5_V_read_9_reg_10245_pp0_iter3_reg);

assign add_ln703_168_fu_967_p2 = (add_ln703_161_reg_10487 + add_ln703_166_fu_962_p2);

assign add_ln703_170_fu_972_p2 = (add_ln703_161_reg_10487 + add_ln703_149_fu_773_p2);

assign add_ln703_171_fu_977_p2 = (sub_ln703_51_fu_897_p2 + data_7_V_read_9_reg_10191_pp0_iter3_reg);

assign add_ln703_173_fu_982_p2 = (add_ln703_161_reg_10487 + sub_ln703_36_fu_795_p2);

assign add_ln703_174_fu_1114_p2 = (sub_ln703_54_fu_1086_p2 + data_8_V_read_8_reg_10164_pp0_iter4_reg);

assign add_ln703_175_fu_1123_p2 = (sub_ln703_55_fu_1090_p2 + data_8_V_read_8_reg_10164_pp0_iter4_reg);

assign add_ln703_176_fu_1128_p2 = (sub_ln703_56_fu_1094_p2 + data_8_V_read_8_reg_10164_pp0_iter4_reg);

assign add_ln703_177_fu_997_p2 = (sub_ln703_61_fu_932_p2 + data_8_V_read_8_reg_10164_pp0_iter3_reg);

assign add_ln703_178_fu_1007_p2 = (sub_ln703_17_reg_10453 + data_5_V_read_9_reg_10245_pp0_iter3_reg);

assign add_ln703_179_fu_685_p2 = (data_7_V_read_9_reg_10191_pp0_iter2_reg + data_8_V_read_8_reg_10164_pp0_iter2_reg);

assign add_ln703_180_fu_1011_p2 = (add_ln703_179_reg_10495 + data_6_V_read_9_reg_10218_pp0_iter3_reg);

assign add_ln703_181_fu_1015_p2 = (add_ln703_180_fu_1011_p2 + add_ln703_178_fu_1007_p2);

assign add_ln703_183_fu_1021_p2 = (add_ln703_179_reg_10495 + sub_ln703_47_fu_863_p2);

assign add_ln703_184_fu_1143_p2 = (sub_ln703_62_reg_10550 + data_8_V_read_8_reg_10164_pp0_iter4_reg);

assign add_ln703_186_fu_1036_p2 = (add_ln703_179_reg_10495 + sub_ln703_50_fu_887_p2);

assign add_ln703_187_fu_1041_p2 = (sub_ln703_28_reg_10476 + data_6_V_read_9_reg_10218_pp0_iter3_reg);

assign add_ln703_189_fu_1045_p2 = (add_ln703_179_reg_10495 + add_ln703_187_fu_1041_p2);

assign add_ln703_190_fu_1172_p2 = (sub_ln703_64_reg_10560 + data_8_V_read_8_reg_10164_pp0_iter4_reg);

assign add_ln703_191_fu_1176_p2 = (sub_ln703_66_reg_10581 + data_8_V_read_8_reg_10164_pp0_iter4_reg);

assign add_ln703_192_fu_1050_p2 = (data_8_V_read_8_reg_10164_pp0_iter3_reg + data_9_V_read_8_reg_10136_pp0_iter3_reg);

assign add_ln703_193_fu_1180_p2 = (add_ln703_192_reg_10626 + sub_ln703_53_reg_10534);

assign add_ln703_194_fu_1189_p2 = (sub_ln703_67_fu_1119_p2 + data_9_V_read_8_reg_10136_pp0_iter4_reg);

assign add_ln703_195_fu_1204_p2 = (sub_ln703_69_fu_1138_p2 + data_9_V_read_8_reg_10136_pp0_iter4_reg);

assign add_ln703_197_fu_1209_p2 = (add_ln703_192_reg_10626 + sub_ln703_58_reg_10545);

assign add_ln703_199_fu_1213_p2 = (add_ln703_192_reg_10626 + sub_ln703_59_fu_1106_p2);

assign add_ln703_200_fu_1226_p2 = (sub_ln703_71_reg_10596 + data_9_V_read_8_reg_10136_pp0_iter4_reg);

assign add_ln703_201_fu_1243_p2 = (sub_ln703_72_fu_1147_p2 + data_9_V_read_8_reg_10136_pp0_iter4_reg);

assign add_ln703_202_fu_1265_p2 = (sub_ln703_77_fu_1159_p2 + data_9_V_read_8_reg_10136_pp0_iter4_reg);

assign add_ln703_203_fu_1270_p2 = (sub_ln703_78_fu_1164_p2 + data_9_V_read_8_reg_10136_pp0_iter4_reg);

assign add_ln703_204_fu_1059_p2 = (sub_ln703_52_fu_907_p2 + data_7_V_read_9_reg_10191_pp0_iter3_reg);

assign add_ln703_206_fu_1290_p2 = (add_ln703_192_reg_10626 + add_ln703_204_reg_10641);

assign add_ln703_207_fu_1299_p2 = (sub_ln703_80_fu_1184_p2 + data_10_V_read11_reg_10105_pp0_iter4_reg);

assign add_ln703_208_fu_1309_p2 = (sub_ln703_82_fu_1199_p2 + data_10_V_read11_reg_10105_pp0_iter4_reg);

assign add_ln703_209_fu_1064_p2 = (data_9_V_read_8_reg_10136_pp0_iter3_reg + data_10_V_read11_reg_10105_pp0_iter3_reg);

assign add_ln703_210_fu_1314_p2 = (add_ln703_209_reg_10646 + sub_ln703_68_fu_1133_p2);

assign add_ln703_211_fu_1339_p2 = (sub_ln703_84_fu_1222_p2 + data_10_V_read11_reg_10105_pp0_iter4_reg);

assign add_ln703_213_fu_1068_p2 = (sub_ln703_46_fu_858_p2 + data_10_V_read11_reg_10105_pp0_iter3_reg);

assign add_ln703_214_fu_1349_p2 = (add_ln703_213_reg_10653 + data_7_V_read_9_reg_10191_pp0_iter4_reg);

assign add_ln703_215_fu_1353_p2 = (add_ln703_214_fu_1349_p2 + add_ln703_192_reg_10626);

assign add_ln703_216_fu_1358_p2 = (sub_ln703_85_fu_1230_p2 + data_10_V_read11_reg_10105_pp0_iter4_reg);

assign add_ln703_217_fu_1393_p2 = (add_ln703_162_reg_10539 + data_8_V_read_8_reg_10164_pp0_iter4_reg);

assign add_ln703_219_fu_1397_p2 = (add_ln703_209_reg_10646 + add_ln703_217_fu_1393_p2);

assign add_ln703_221_fu_1402_p2 = (add_ln703_209_reg_10646 + sub_ln703_76_fu_1155_p2);

assign add_ln703_222_fu_1626_p2 = (sub_ln703_96_reg_10677 + data_11_V_read12_reg_10075_pp0_iter5_reg);

assign add_ln703_223_fu_1073_p2 = (data_10_V_read11_reg_10105_pp0_iter3_reg + data_11_V_read12_reg_10075_pp0_iter3_reg);

assign add_ln703_224_fu_1437_p2 = (add_ln703_223_reg_10658 + sub_ln703_81_fu_1194_p2);

assign add_ln703_225_fu_1452_p2 = (sub_ln703_102_fu_1344_p2 + data_11_V_read12_reg_10075_pp0_iter4_reg);

assign add_ln703_226_fu_1457_p2 = (add_ln703_215_fu_1353_p2 + data_11_V_read12_reg_10075_pp0_iter4_reg);

assign add_ln703_227_fu_1472_p2 = (sub_ln703_104_fu_1368_p2 + data_11_V_read12_reg_10075_pp0_iter4_reg);

assign add_ln703_228_fu_1477_p2 = (sub_ln703_105_fu_1373_p2 + data_11_V_read12_reg_10075_pp0_iter4_reg);

assign add_ln703_229_fu_1654_p2 = (sub_ln703_107_reg_10712 + data_11_V_read12_reg_10075_pp0_iter5_reg);

assign add_ln703_230_fu_1658_p2 = (sub_ln703_108_reg_10717 + data_11_V_read12_reg_10075_pp0_iter5_reg);

assign add_ln703_232_fu_1492_p2 = (add_ln703_223_reg_10658 + sub_ln703_92_reg_10636);

assign add_ln703_233_fu_1501_p2 = (sub_ln703_112_fu_1422_p2 + data_11_V_read12_reg_10075_pp0_iter4_reg);

assign add_ln703_234_fu_1671_p2 = (sub_ln703_114_fu_1630_p2 + data_12_V_read13_reg_10045_pp0_iter5_reg);

assign add_ln703_235_fu_1676_p2 = (sub_ln703_115_reg_10727 + data_12_V_read13_reg_10045_pp0_iter5_reg);

assign add_ln703_236_fu_1511_p2 = (sub_ln703_119_fu_1442_p2 + data_12_V_read13_reg_10045_pp0_iter4_reg);

assign add_ln703_237_fu_1516_p2 = (data_11_V_read12_reg_10075_pp0_iter4_reg + data_12_V_read13_reg_10045_pp0_iter4_reg);

assign add_ln703_238_fu_1520_p2 = (add_ln703_237_fu_1516_p2 + sub_ln703_100_fu_1329_p2);

assign add_ln703_240_fu_1526_p2 = (add_ln703_237_fu_1516_p2 + sub_ln703_101_fu_1334_p2);

assign add_ln703_241_fu_1693_p2 = (sub_ln703_121_fu_1646_p2 + data_12_V_read13_reg_10045_pp0_iter5_reg);

assign add_ln703_242_fu_1537_p2 = (sub_ln703_86_fu_1234_p2 + data_10_V_read11_reg_10105_pp0_iter4_reg);

assign add_ln703_244_fu_1542_p2 = (add_ln703_237_fu_1516_p2 + add_ln703_242_fu_1537_p2);

assign add_ln703_245_fu_1721_p2 = (sub_ln703_125_reg_10757 + data_12_V_read13_reg_10045_pp0_iter5_reg);

assign add_ln703_247_fu_1563_p2 = (add_ln703_237_fu_1516_p2 + sub_ln703_110_fu_1412_p2);

assign add_ln703_248_fu_1569_p2 = (sub_ln703_95_fu_1285_p2 + data_10_V_read11_reg_10105_pp0_iter4_reg);

assign add_ln703_250_fu_1574_p2 = (add_ln703_237_fu_1516_p2 + add_ln703_248_fu_1569_p2);

assign add_ln703_251_fu_1753_p2 = (sub_ln703_131_fu_1680_p2 + data_13_V_read14_reg_10015_pp0_iter5_reg);

assign add_ln703_252_fu_1077_p2 = (data_12_V_read13_reg_10045_pp0_iter3_reg + data_13_V_read14_reg_10015_pp0_iter3_reg);

assign add_ln703_253_fu_1758_p2 = (add_ln703_252_reg_10665_pp0_iter5_reg + sub_ln703_117_fu_1638_p2);

assign add_ln703_254_fu_1081_p2 = (sub_ln703_42_fu_833_p2 + data_7_V_read_9_reg_10191_pp0_iter3_reg);

assign add_ln703_256_fu_1585_p2 = (add_ln703_192_reg_10626 + add_ln703_254_reg_10672);

assign add_ln703_259_fu_1589_p2 = (add_ln703_252_reg_10665 + add_ln703_223_reg_10658);

assign add_ln703_260_fu_1593_p2 = (add_ln703_259_fu_1589_p2 + add_ln703_256_fu_1585_p2);

assign add_ln703_262_fu_1604_p2 = (add_ln703_252_reg_10665 + sub_ln703_120_fu_1447_p2);

assign add_ln703_263_fu_1771_p2 = (sub_ln703_133_reg_10782 + data_13_V_read14_reg_10015_pp0_iter5_reg);

assign add_ln703_264_fu_1821_p2 = (sub_ln703_145_fu_1734_p2 + data_13_V_read14_reg_10015_pp0_iter5_reg);

assign add_ln703_265_fu_1614_p2 = (data_13_V_read14_reg_10015_pp0_iter4_reg + data_14_V_read15_reg_9987_pp0_iter4_reg);

assign add_ln703_266_fu_1854_p2 = (add_ln703_265_reg_10837 + sub_ln703_132_fu_1684_p2);

assign add_ln703_268_fu_1886_p2 = (add_ln703_265_reg_10837 + sub_ln703_134_fu_1689_p2);

assign add_ln703_269_fu_1891_p2 = (sub_ln703_122_reg_10742 + data_12_V_read13_reg_10045_pp0_iter5_reg);

assign add_ln703_271_fu_1895_p2 = (add_ln703_265_reg_10837 + add_ln703_269_fu_1891_p2);

assign add_ln703_273_fu_1914_p2 = (add_ln703_265_reg_10837 + sub_ln703_138_fu_1706_p2);

assign add_ln703_274_fu_1924_p2 = (sub_ln703_161_fu_1809_p2 + data_14_V_read15_reg_9987_pp0_iter5_reg);

assign add_ln703_276_fu_1934_p2 = (add_ln703_265_reg_10837 + sub_ln703_143_fu_1725_p2);

assign add_ln703_277_fu_1939_p2 = (sub_ln703_163_fu_1817_p2 + data_14_V_read15_reg_9987_pp0_iter5_reg);

assign add_ln703_278_fu_1954_p2 = (sub_ln703_165_fu_1830_p2 + data_14_V_read15_reg_9987_pp0_iter5_reg);

assign add_ln703_279_fu_1964_p2 = (sub_ln703_116_fu_1634_p2 + data_12_V_read13_reg_10045_pp0_iter5_reg);

assign add_ln703_280_fu_1618_p2 = (data_14_V_read15_reg_9987_pp0_iter4_reg + data_15_V_read16_reg_9962_pp0_iter4_reg);

assign add_ln703_281_fu_1969_p2 = (add_ln703_280_reg_10846 + data_13_V_read14_reg_10015_pp0_iter5_reg);

assign add_ln703_282_fu_1973_p2 = (add_ln703_281_fu_1969_p2 + add_ln703_279_fu_1964_p2);

assign add_ln703_283_fu_1979_p2 = (sub_ln703_169_fu_1849_p2 + data_15_V_read16_reg_9962_pp0_iter5_reg);

assign add_ln703_285_fu_2009_p2 = (add_ln703_280_reg_10846 + sub_ln703_153_fu_1775_p2);

assign add_ln703_287_fu_2019_p2 = (add_ln703_280_reg_10846 + sub_ln703_155_fu_1780_p2);

assign add_ln703_289_fu_2034_p2 = (add_ln703_280_reg_10846 + sub_ln703_158_fu_1794_p2);

assign add_ln703_290_fu_2039_p2 = (sub_ln703_179_fu_1919_p2 + data_15_V_read16_reg_9962_pp0_iter5_reg);

assign add_ln703_291_fu_2064_p2 = (sub_ln703_144_fu_1730_p2 + data_13_V_read14_reg_10015_pp0_iter5_reg);

assign add_ln703_293_fu_2069_p2 = (add_ln703_280_reg_10846 + add_ln703_291_fu_2064_p2);

assign add_ln703_294_fu_2084_p2 = (sub_ln703_147_fu_1738_p2 + data_14_V_read15_reg_9987_pp0_iter5_reg);

assign add_ln703_295_fu_2089_p2 = (data_15_V_read16_reg_9962_pp0_iter5_reg + data_16_V_read17_reg_9935_pp0_iter5_reg);

assign add_ln703_296_fu_2238_p2 = (add_ln703_295_reg_10923 + add_ln703_294_reg_10918);

assign add_ln703_298_fu_2242_p2 = (add_ln703_295_reg_10923 + sub_ln703_166_reg_10863);

assign add_ln703_300_fu_2093_p2 = (add_ln703_295_fu_2089_p2 + sub_ln703_167_fu_1839_p2);

assign add_ln703_301_fu_2250_p2 = (sub_ln703_184_reg_10878 + data_16_V_read17_reg_9935_pp0_iter6_reg);

assign add_ln703_303_fu_2104_p2 = (add_ln703_295_fu_2089_p2 + sub_ln703_171_fu_1864_p2);

assign add_ln703_304_fu_2110_p2 = (sub_ln703_185_fu_1989_p2 + data_16_V_read17_reg_9935_pp0_iter5_reg);

assign add_ln703_305_fu_2254_p2 = (sub_ln703_186_reg_10883 + data_16_V_read17_reg_9935_pp0_iter6_reg);

assign add_ln703_307_fu_2125_p2 = (add_ln703_295_fu_2089_p2 + sub_ln703_176_fu_1900_p2);

assign add_ln703_309_fu_2136_p2 = (add_ln703_295_fu_2089_p2 + sub_ln703_177_fu_1904_p2);

assign add_ln703_310_fu_2147_p2 = (sub_ln703_159_fu_1799_p2 + data_14_V_read15_reg_9987_pp0_iter5_reg);

assign add_ln703_312_fu_2270_p2 = (add_ln703_295_reg_10923 + add_ln703_310_reg_10980);

assign add_ln703_314_fu_2167_p2 = (add_ln703_295_fu_2089_p2 + sub_ln703_182_fu_1949_p2);

assign add_ln703_315_fu_2300_p2 = (sub_ln703_199_fu_2246_p2 + data_17_V_read18_reg_9904_pp0_iter6_reg);

assign add_ln703_316_fu_2178_p2 = (data_16_V_read17_reg_9935_pp0_iter5_reg + data_17_V_read18_reg_9904_pp0_iter5_reg);

assign add_ln703_317_fu_2182_p2 = (add_ln703_316_fu_2178_p2 + sub_ln703_187_fu_1999_p2);

assign add_ln703_318_fu_2323_p2 = (sub_ln703_201_fu_2258_p2 + data_17_V_read18_reg_9904_pp0_iter6_reg);

assign add_ln703_319_fu_2328_p2 = (sub_ln703_202_reg_10955 + data_17_V_read18_reg_9904_pp0_iter6_reg);

assign add_ln703_320_fu_2336_p2 = (sub_ln703_203_reg_10965 + data_17_V_read18_reg_9904_pp0_iter6_reg);

assign add_ln703_321_fu_2353_p2 = (sub_ln703_206_fu_2266_p2 + data_17_V_read18_reg_9904_pp0_iter6_reg);

assign add_ln703_323_fu_2188_p2 = (add_ln703_316_fu_2178_p2 + sub_ln703_193_fu_2049_p2);

assign add_ln703_324_fu_2405_p2 = (sub_ln703_217_fu_2305_p2 + data_18_V_read_8_reg_9874_pp0_iter6_reg);

assign add_ln703_325_fu_2199_p2 = (sub_ln703_170_fu_1859_p2 + data_15_V_read16_reg_9962_pp0_iter5_reg);

assign add_ln703_326_fu_1622_p2 = (data_17_V_read18_reg_9904_pp0_iter4_reg + data_18_V_read_8_reg_9874_pp0_iter4_reg);

assign add_ln703_327_fu_2204_p2 = (add_ln703_326_reg_10855 + data_16_V_read17_reg_9935_pp0_iter5_reg);

assign add_ln703_328_fu_2208_p2 = (add_ln703_327_fu_2204_p2 + add_ln703_325_fu_2199_p2);

assign add_ln703_329_fu_2410_p2 = (sub_ln703_218_fu_2310_p2 + data_18_V_read_8_reg_9874_pp0_iter6_reg);

assign add_ln703_330_fu_2219_p2 = (sub_ln703_175_fu_1881_p2 + data_15_V_read16_reg_9962_pp0_iter5_reg);

assign add_ln703_333_fu_2224_p2 = (add_ln703_327_fu_2204_p2 + add_ln703_330_fu_2219_p2);

assign add_ln703_335_fu_2420_p2 = (add_ln703_326_reg_10855_pp0_iter6_reg + sub_ln703_200_reg_10950);

assign add_ln703_336_fu_2449_p2 = (sub_ln703_224_fu_2348_p2 + data_18_V_read_8_reg_9874_pp0_iter6_reg);

assign add_ln703_337_fu_2459_p2 = (sub_ln703_225_fu_2358_p2 + data_18_V_read_8_reg_9874_pp0_iter6_reg);

assign add_ln703_339_fu_2464_p2 = (add_ln703_326_reg_10855_pp0_iter6_reg + sub_ln703_208_reg_10985);

assign add_ln703_340_fu_2491_p2 = (sub_ln703_231_fu_2381_p2 + data_18_V_read_8_reg_9874_pp0_iter6_reg);

assign add_ln703_341_fu_2230_p2 = (data_18_V_read_8_reg_9874_pp0_iter5_reg + data_19_V_read_8_reg_9845_pp0_iter5_reg);

assign add_ln703_342_fu_2520_p2 = (add_ln703_341_reg_11030 + sub_ln703_219_fu_2314_p2);

assign add_ln703_343_fu_2554_p2 = (sub_ln703_241_fu_2439_p2 + data_19_V_read_8_reg_9845_pp0_iter6_reg);

assign add_ln703_345_fu_2564_p2 = (add_ln703_341_reg_11030 + sub_ln703_223_fu_2344_p2);

assign add_ln703_346_fu_2589_p2 = (sub_ln703_244_fu_2468_p2 + data_19_V_read_8_reg_9845_pp0_iter6_reg);

assign add_ln703_347_fu_2594_p2 = (sub_ln703_194_reg_10908 + data_16_V_read17_reg_9935_pp0_iter6_reg);

assign add_ln703_349_fu_2598_p2 = (add_ln703_341_reg_11030 + data_17_V_read18_reg_9904_pp0_iter6_reg);

assign add_ln703_350_fu_2602_p2 = (add_ln703_349_fu_2598_p2 + add_ln703_347_fu_2594_p2);

assign add_ln703_351_fu_2608_p2 = (sub_ln703_245_fu_2472_p2 + data_19_V_read_8_reg_9845_pp0_iter6_reg);

assign add_ln703_352_fu_2633_p2 = (sub_ln703_253_fu_2515_p2 + data_20_V_read21_reg_9814_pp0_iter6_reg);

assign add_ln703_353_fu_2795_p2 = (sub_ln703_254_reg_11076 + data_20_V_read21_reg_9814_pp0_iter7_reg);

assign add_ln703_354_fu_2638_p2 = (data_19_V_read_8_reg_9845_pp0_iter6_reg + data_20_V_read21_reg_9814_pp0_iter6_reg);

assign add_ln703_355_fu_2642_p2 = (add_ln703_354_fu_2638_p2 + sub_ln703_237_reg_11020);

assign add_ln703_356_fu_2657_p2 = (sub_ln703_259_fu_2549_p2 + data_20_V_read21_reg_9814_pp0_iter6_reg);

assign add_ln703_357_fu_2811_p2 = (sub_ln703_263_reg_11101 + data_20_V_read21_reg_9814_pp0_iter7_reg);

assign add_ln703_358_fu_2672_p2 = (sub_ln703_226_fu_2363_p2 + data_18_V_read_8_reg_9874_pp0_iter6_reg);

assign add_ln703_360_fu_2677_p2 = (add_ln703_354_fu_2638_p2 + add_ln703_358_fu_2672_p2);

assign add_ln703_361_fu_2683_p2 = (sub_ln703_264_fu_2584_p2 + data_20_V_read21_reg_9814_pp0_iter6_reg);

assign add_ln703_363_fu_2823_p2 = (add_ln703_354_reg_11131 + sub_ln703_246_reg_11051);

assign add_ln703_364_fu_2831_p2 = (sub_ln703_268_fu_2783_p2 + data_21_V_read22_reg_9784_pp0_iter7_reg);

assign add_ln703_365_fu_2841_p2 = (sub_ln703_270_reg_11121 + data_21_V_read22_reg_9784_pp0_iter7_reg);

assign add_ln703_366_fu_2871_p2 = (sub_ln703_275_reg_11153 + data_21_V_read22_reg_9784_pp0_iter7_reg);

assign add_ln703_367_fu_2903_p2 = (sub_ln703_284_reg_11168 + data_21_V_read22_reg_9784_pp0_iter7_reg);

assign add_ln703_368_fu_2723_p2 = (sub_ln703_233_fu_2390_p2 + data_19_V_read_8_reg_9845_pp0_iter6_reg);

assign add_ln703_369_fu_2234_p2 = (data_21_V_read22_reg_9784_pp0_iter5_reg + data_22_V_read23_reg_9756_pp0_iter5_reg);

assign add_ln703_370_fu_2728_p2 = (add_ln703_369_reg_11037 + data_20_V_read21_reg_9814_pp0_iter6_reg);

assign add_ln703_371_fu_2732_p2 = (add_ln703_370_fu_2728_p2 + add_ln703_368_fu_2723_p2);

assign add_ln703_372_fu_2927_p2 = (sub_ln703_289_reg_11173 + data_22_V_read23_reg_9756_pp0_iter7_reg);

assign add_ln703_374_fu_2936_p2 = (add_ln703_369_reg_11037_pp0_iter7_reg + sub_ln703_273_fu_2799_p2);

assign add_ln703_375_fu_2738_p2 = (sub_ln703_260_fu_2559_p2 + data_20_V_read21_reg_9814_pp0_iter6_reg);

assign add_ln703_377_fu_2956_p2 = (add_ln703_369_reg_11037_pp0_iter7_reg + add_ln703_375_reg_11198);

assign add_ln703_378_fu_2960_p2 = (sub_ln703_293_reg_11178 + data_22_V_read23_reg_9756_pp0_iter7_reg);

assign add_ln703_379_fu_2964_p2 = (sub_ln703_295_fu_2880_p2 + data_22_V_read23_reg_9756_pp0_iter7_reg);

assign add_ln703_380_fu_2969_p2 = (sub_ln703_296_reg_11183 + data_22_V_read23_reg_9756_pp0_iter7_reg);

assign add_ln703_381_fu_2973_p2 = (sub_ln703_297_fu_2884_p2 + data_22_V_read23_reg_9756_pp0_iter7_reg);

assign add_ln703_382_fu_2983_p2 = (sub_ln703_299_fu_2894_p2 + data_22_V_read23_reg_9756_pp0_iter7_reg);

assign add_ln703_383_fu_3007_p2 = (sub_ln703_250_reg_11061 + data_20_V_read21_reg_9814_pp0_iter7_reg);

assign add_ln703_384_fu_2743_p2 = (data_22_V_read23_reg_9756_pp0_iter6_reg + data_23_V_read24_reg_9730_pp0_iter6_reg);

assign add_ln703_385_fu_3011_p2 = (add_ln703_384_reg_11203 + data_21_V_read22_reg_9784_pp0_iter7_reg);

assign add_ln703_386_fu_3015_p2 = (add_ln703_385_fu_3011_p2 + add_ln703_383_fu_3007_p2);

assign add_ln703_387_fu_3046_p2 = (sub_ln703_257_reg_11086 + data_20_V_read21_reg_9814_pp0_iter7_reg);

assign add_ln703_390_fu_3050_p2 = (add_ln703_385_fu_3011_p2 + add_ln703_387_fu_3046_p2);

assign add_ln703_391_fu_3061_p2 = (sub_ln703_308_fu_2946_p2 + data_23_V_read24_reg_9730_pp0_iter7_reg);

assign add_ln703_392_fu_3081_p2 = (sub_ln703_277_fu_2803_p2 + data_21_V_read22_reg_9784_pp0_iter7_reg);

assign add_ln703_394_fu_3086_p2 = (add_ln703_384_reg_11203 + add_ln703_392_fu_3081_p2);

assign add_ln703_395_fu_3116_p2 = (sub_ln703_282_fu_2827_p2 + data_21_V_read22_reg_9784_pp0_iter7_reg);

assign add_ln703_397_fu_3121_p2 = (add_ln703_384_reg_11203 + add_ln703_395_fu_3116_p2);

assign add_ln703_398_fu_2747_p2 = (sub_ln703_214_fu_2287_p2 + data_18_V_read_8_reg_9874_pp0_iter6_reg);

assign add_ln703_400_fu_2752_p2 = (add_ln703_354_fu_2638_p2 + add_ln703_398_fu_2747_p2);

assign add_ln703_402_fu_2758_p2 = (data_23_V_read24_reg_9730_pp0_iter6_reg + data_24_V_read25_reg_9704_pp0_iter6_reg);

assign add_ln703_403_fu_3131_p2 = (add_ln703_402_reg_11215 + add_ln703_369_reg_11037_pp0_iter7_reg);

assign add_ln703_404_fu_3135_p2 = (add_ln703_403_fu_3131_p2 + add_ln703_400_reg_11210);

assign add_ln703_406_fu_3145_p2 = (add_ln703_354_reg_11131 + sub_ln703_234_reg_11046);

assign add_ln703_410_fu_3149_p2 = (add_ln703_403_fu_3131_p2 + add_ln703_406_fu_3145_p2);

assign add_ln703_411_fu_3380_p2 = (sub_ln703_315_reg_11267 + data_24_V_read25_reg_9704_pp0_iter8_reg);

assign add_ln703_413_fu_3160_p2 = (add_ln703_402_reg_11215 + sub_ln703_305_fu_2922_p2);

assign add_ln703_414_fu_3165_p2 = (sub_ln703_288_fu_2854_p2 + data_22_V_read23_reg_9756_pp0_iter7_reg);

assign add_ln703_416_fu_3170_p2 = (add_ln703_402_reg_11215 + add_ln703_414_fu_3165_p2);

assign add_ln703_417_fu_3185_p2 = (sub_ln703_321_fu_3066_p2 + data_24_V_read25_reg_9704_pp0_iter7_reg);

assign add_ln703_418_fu_3210_p2 = (sub_ln703_325_fu_3096_p2 + data_24_V_read25_reg_9704_pp0_iter7_reg);

assign add_ln703_419_fu_3225_p2 = (sub_ln703_301_reg_11188 + data_22_V_read23_reg_9756_pp0_iter7_reg);

assign add_ln703_421_fu_3229_p2 = (add_ln703_402_reg_11215 + add_ln703_419_fu_3225_p2);

assign add_ln703_422_fu_3239_p2 = (sub_ln703_331_fu_3140_p2 + data_25_V_read26_reg_9677_pp0_iter7_reg);

assign add_ln703_423_fu_3249_p2 = (sub_ln703_287_fu_2849_p2 + data_22_V_read23_reg_9756_pp0_iter7_reg);

assign add_ln703_424_fu_2762_p2 = (data_24_V_read25_reg_9704_pp0_iter6_reg + data_25_V_read26_reg_9677_pp0_iter6_reg);

assign add_ln703_425_fu_3254_p2 = (add_ln703_424_reg_11225 + data_23_V_read24_reg_9730_pp0_iter7_reg);

assign add_ln703_426_fu_3258_p2 = (add_ln703_425_fu_3254_p2 + add_ln703_423_fu_3249_p2);

assign add_ln703_428_fu_3264_p2 = (add_ln703_424_reg_11225 + sub_ln703_317_fu_3031_p2);

assign add_ln703_429_fu_3418_p2 = (sub_ln703_335_fu_3384_p2 + data_25_V_read26_reg_9677_pp0_iter8_reg);

assign add_ln703_430_fu_3423_p2 = (sub_ln703_336_reg_11307 + data_25_V_read26_reg_9677_pp0_iter8_reg);

assign add_ln703_431_fu_3274_p2 = (sub_ln703_338_fu_3195_p2 + data_25_V_read26_reg_9677_pp0_iter7_reg);

assign add_ln703_432_fu_3279_p2 = (sub_ln703_294_fu_2875_p2 + data_22_V_read23_reg_9756_pp0_iter7_reg);

assign add_ln703_435_fu_3284_p2 = (add_ln703_425_fu_3254_p2 + add_ln703_432_fu_3279_p2);

assign add_ln703_436_fu_3439_p2 = (sub_ln703_342_reg_11327 + data_25_V_read26_reg_9677_pp0_iter8_reg);

assign add_ln703_437_fu_3443_p2 = (sub_ln703_346_fu_3396_p2 + data_26_V_read27_reg_9652_pp0_iter8_reg);

assign add_ln703_438_fu_3310_p2 = (sub_ln703_320_fu_3056_p2 + data_24_V_read25_reg_9704_pp0_iter7_reg);

assign add_ln703_439_fu_2766_p2 = (data_25_V_read26_reg_9677_pp0_iter6_reg + data_26_V_read27_reg_9652_pp0_iter6_reg);

assign add_ln703_440_fu_3466_p2 = (add_ln703_439_reg_11233_pp0_iter8_reg + add_ln703_438_reg_11382);

assign add_ln703_441_fu_3480_p2 = (sub_ln703_353_reg_11352 + data_26_V_read27_reg_9652_pp0_iter8_reg);

assign add_ln703_442_fu_3502_p2 = (sub_ln703_356_reg_11367 + data_26_V_read27_reg_9652_pp0_iter8_reg);

assign add_ln703_444_fu_3506_p2 = (add_ln703_439_reg_11233_pp0_iter8_reg + sub_ln703_341_fu_3388_p2);

assign add_ln703_445_fu_3315_p2 = (sub_ln703_310_fu_2978_p2 + data_23_V_read24_reg_9730_pp0_iter7_reg);

assign add_ln703_447_fu_3320_p2 = (add_ln703_439_reg_11233 + data_24_V_read25_reg_9704_pp0_iter7_reg);

assign add_ln703_448_fu_3511_p2 = (add_ln703_447_reg_11392 + add_ln703_445_reg_11387);

assign add_ln703_450_fu_3520_p2 = (add_ln703_439_reg_11233_pp0_iter8_reg + sub_ln703_344_reg_11332);

assign add_ln703_451_fu_3329_p2 = (data_26_V_read27_reg_9652_pp0_iter7_reg + data_27_V_read28_reg_9625_pp0_iter7_reg);

assign add_ln703_452_fu_3524_p2 = (add_ln703_451_reg_11402 + sub_ln703_345_reg_11337);

assign add_ln703_453_fu_3528_p2 = (sub_ln703_358_reg_11372 + data_27_V_read28_reg_9625_pp0_iter8_reg);

assign add_ln703_455_fu_3537_p2 = (add_ln703_451_reg_11402 + sub_ln703_348_fu_3405_p2);

assign add_ln703_456_fu_3542_p2 = (sub_ln703_359_fu_3448_p2 + data_27_V_read28_reg_9625_pp0_iter8_reg);

assign add_ln703_458_fu_3552_p2 = (add_ln703_451_reg_11402 + sub_ln703_351_fu_3414_p2);

assign add_ln703_459_fu_3557_p2 = (sub_ln703_334_reg_11302 + data_25_V_read26_reg_9677_pp0_iter8_reg);

assign add_ln703_461_fu_3561_p2 = (add_ln703_451_reg_11402 + add_ln703_459_fu_3557_p2);

assign add_ln703_462_fu_3571_p2 = (sub_ln703_364_fu_3470_p2 + data_27_V_read28_reg_9625_pp0_iter8_reg);

assign add_ln703_463_fu_3581_p2 = (sub_ln703_366_fu_3484_p2 + data_27_V_read28_reg_9625_pp0_iter8_reg);

assign add_ln703_464_fu_3586_p2 = (sub_ln703_367_fu_3488_p2 + data_27_V_read28_reg_9625_pp0_iter8_reg);

assign add_ln703_465_fu_3630_p2 = (sub_ln703_330_fu_3372_p2 + data_25_V_read26_reg_9677_pp0_iter8_reg);

assign add_ln703_466_fu_3333_p2 = (data_27_V_read28_reg_9625_pp0_iter7_reg + data_28_V_read_8_reg_9598_pp0_iter7_reg);

assign add_ln703_467_fu_3635_p2 = (add_ln703_466_reg_11410 + data_26_V_read27_reg_9652_pp0_iter8_reg);

assign add_ln703_468_fu_3639_p2 = (add_ln703_467_fu_3635_p2 + add_ln703_465_fu_3630_p2);

assign add_ln703_469_fu_3655_p2 = (sub_ln703_372_fu_3532_p2 + data_28_V_read_8_reg_9598_pp0_iter8_reg);

assign add_ln703_471_fu_3337_p2 = (add_ln703_424_reg_11225 + sub_ln703_319_fu_3041_p2);

assign add_ln703_474_fu_3680_p2 = (add_ln703_467_fu_3635_p2 + add_ln703_471_reg_11418);

assign add_ln703_476_fu_3685_p2 = (add_ln703_466_reg_11410 + sub_ln703_363_fu_3461_p2);

assign add_ln703_477_fu_3715_p2 = (sub_ln703_378_fu_3601_p2 + data_28_V_read_8_reg_9598_pp0_iter8_reg);

assign add_ln703_478_fu_3730_p2 = (sub_ln703_381_fu_3616_p2 + data_28_V_read_8_reg_9598_pp0_iter8_reg);

assign add_ln703_479_fu_3735_p2 = (sub_ln703_343_fu_3392_p2 + data_25_V_read26_reg_9677_pp0_iter8_reg);

assign add_ln703_482_fu_3740_p2 = (add_ln703_467_fu_3635_p2 + add_ln703_479_fu_3735_p2);

assign add_ln703_484_fu_3342_p2 = (add_ln703_424_reg_11225 + sub_ln703_329_fu_3126_p2);

assign add_ln703_487_fu_3756_p2 = (add_ln703_467_fu_3635_p2 + add_ln703_484_reg_11423);

assign add_ln703_488_fu_3766_p2 = (sub_ln703_385_fu_3650_p2 + data_29_V_read_8_reg_9573_pp0_iter8_reg);

assign add_ln703_489_fu_3771_p2 = (sub_ln703_361_fu_3457_p2 + data_27_V_read28_reg_9625_pp0_iter8_reg);

assign add_ln703_490_fu_3347_p2 = (data_28_V_read_8_reg_9598_pp0_iter7_reg + data_29_V_read_8_reg_9573_pp0_iter7_reg);

assign add_ln703_491_fu_3776_p2 = (add_ln703_490_reg_11428 + add_ln703_489_fu_3771_p2);

assign add_ln703_493_fu_3796_p2 = (add_ln703_490_reg_11428 + sub_ln703_374_fu_3566_p2);

assign add_ln703_494_fu_3801_p2 = (sub_ln703_365_fu_3475_p2 + data_27_V_read28_reg_9625_pp0_iter8_reg);

assign add_ln703_496_fu_3806_p2 = (add_ln703_490_reg_11428 + add_ln703_494_fu_3801_p2);

assign add_ln703_497_fu_3811_p2 = (sub_ln703_391_fu_3695_p2 + data_29_V_read_8_reg_9573_pp0_iter8_reg);

assign add_ln703_498_fu_3351_p2 = (sub_ln703_278_fu_2807_p2 + data_21_V_read22_reg_9784_pp0_iter7_reg);

assign add_ln703_500_fu_3821_p2 = (add_ln703_402_reg_11215_pp0_iter8_reg + data_22_V_read23_reg_9756_pp0_iter8_reg);

assign add_ln703_501_fu_3825_p2 = (add_ln703_500_fu_3821_p2 + add_ln703_498_reg_11436);

assign add_ln703_504_fu_3830_p2 = (add_ln703_490_reg_11428 + data_27_V_read28_reg_9625_pp0_iter8_reg);

assign add_ln703_505_fu_3834_p2 = (add_ln703_504_fu_3830_p2 + add_ln703_439_reg_11233_pp0_iter8_reg);

assign add_ln703_506_fu_3839_p2 = (add_ln703_505_fu_3834_p2 + add_ln703_501_fu_3825_p2);

assign add_ln703_507_fu_3356_p2 = (data_29_V_read_8_reg_9573_pp0_iter7_reg + data_30_V_read31_reg_9549_pp0_iter7_reg);

assign add_ln703_508_fu_4006_p2 = (add_ln703_507_reg_11441_pp0_iter9_reg + sub_ln703_386_reg_11484);

assign add_ln703_509_fu_3870_p2 = (sub_ln703_362_reg_11377 + data_27_V_read28_reg_9625_pp0_iter8_reg);

assign add_ln703_511_fu_3874_p2 = (add_ln703_507_reg_11441 + data_28_V_read_8_reg_9598_pp0_iter8_reg);

assign add_ln703_512_fu_3878_p2 = (add_ln703_511_fu_3874_p2 + add_ln703_509_fu_3870_p2);

assign add_ln703_513_fu_4035_p2 = (sub_ln703_407_fu_3985_p2 + data_30_V_read31_reg_9549_pp0_iter9_reg);

assign add_ln703_515_fu_3889_p2 = (add_ln703_507_reg_11441 + sub_ln703_396_fu_3725_p2);

assign add_ln703_517_fu_3894_p2 = (add_ln703_507_reg_11441 + sub_ln703_397_fu_3746_p2);

assign add_ln703_519_fu_3899_p2 = (add_ln703_507_reg_11441 + sub_ln703_398_fu_3751_p2);

assign add_ln703_520_fu_4058_p2 = (sub_ln703_412_reg_11574 + data_30_V_read31_reg_9549_pp0_iter9_reg);

assign add_ln703_521_fu_4062_p2 = (sub_ln703_413_fu_3997_p2 + data_31_V_read32_reg_9521_pp0_iter9_reg);

assign add_ln703_522_fu_4067_p2 = (sub_ln703_414_reg_11579 + data_31_V_read32_reg_9521_pp0_iter9_reg);

assign add_ln703_523_fu_2770_p2 = (sub_ln703_183_reg_10868 + data_16_V_read17_reg_9935_pp0_iter6_reg);

assign add_ln703_525_fu_2774_p2 = (add_ln703_326_reg_10855_pp0_iter6_reg + add_ln703_523_fu_2770_p2);

assign add_ln703_528_fu_3360_p2 = (add_ln703_369_reg_11037_pp0_iter7_reg + add_ln703_354_reg_11131);

assign add_ln703_529_fu_4071_p2 = (add_ln703_528_reg_11452_pp0_iter9_reg + add_ln703_525_reg_11243_pp0_iter9_reg);

assign add_ln703_532_fu_3904_p2 = (add_ln703_439_reg_11233_pp0_iter8_reg + add_ln703_402_reg_11215_pp0_iter8_reg);

assign add_ln703_534_fu_2779_p2 = (data_30_V_read31_reg_9549_pp0_iter6_reg + data_31_V_read32_reg_9521_pp0_iter6_reg);

assign add_ln703_535_fu_3364_p2 = (add_ln703_534_reg_11248 + data_29_V_read_8_reg_9573_pp0_iter7_reg);

assign add_ln703_536_fu_3908_p2 = (add_ln703_535_reg_11457 + add_ln703_466_reg_11410);

assign add_ln703_537_fu_3912_p2 = (add_ln703_536_fu_3908_p2 + add_ln703_532_fu_3904_p2);

assign add_ln703_538_fu_4075_p2 = (add_ln703_537_reg_11609 + add_ln703_529_fu_4071_p2);

assign add_ln703_539_fu_4085_p2 = (sub_ln703_387_reg_11489 + data_29_V_read_8_reg_9573_pp0_iter9_reg);

assign add_ln703_541_fu_4089_p2 = (add_ln703_534_reg_11248_pp0_iter9_reg + add_ln703_539_fu_4085_p2);

assign add_ln703_542_fu_3918_p2 = (sub_ln703_373_fu_3547_p2 + data_28_V_read_8_reg_9598_pp0_iter8_reg);

assign add_ln703_545_fu_3923_p2 = (add_ln703_535_reg_11457 + add_ln703_542_fu_3918_p2);

assign add_ln703_546_fu_4094_p2 = (sub_ln703_416_reg_11584 + data_31_V_read32_reg_9521_pp0_iter9_reg);

assign add_ln703_548_fu_4098_p2 = (add_ln703_534_reg_11248_pp0_iter9_reg + sub_ln703_401_reg_11529);

assign add_ln703_550_fu_4111_p2 = (add_ln703_534_reg_11248_pp0_iter9_reg + sub_ln703_403_reg_11539);

assign add_ln703_551_fu_4115_p2 = (sub_ln703_418_fu_4014_p2 + data_31_V_read32_reg_9521_pp0_iter9_reg);

assign add_ln703_552_fu_4139_p2 = (sub_ln703_423_fu_4031_p2 + data_31_V_read32_reg_9521_pp0_iter9_reg);

assign add_ln703_553_fu_3928_p2 = (sub_ln703_376_fu_3591_p2 + data_28_V_read_8_reg_9598_pp0_iter8_reg);

assign add_ln703_556_fu_3933_p2 = (add_ln703_535_reg_11457 + add_ln703_553_fu_3928_p2);

assign add_ln703_557_fu_4158_p2 = (sub_ln703_426_fu_4049_p2 + data_31_V_read32_reg_9521_pp0_iter9_reg);

assign add_ln703_558_fu_4216_p2 = (sub_ln703_429_fu_4102_p2 + data_32_V_read_3_reg_9492_pp0_iter9_reg);

assign add_ln703_559_fu_4241_p2 = (sub_ln703_432_fu_4124_p2 + data_32_V_read_3_reg_9492_pp0_iter9_reg);

assign add_ln703_560_fu_3943_p2 = (data_31_V_read32_reg_9521_pp0_iter8_reg + data_32_V_read_3_reg_9492_pp0_iter8_reg);

assign add_ln703_561_fu_4260_p2 = (add_ln703_560_reg_11629 + sub_ln703_425_fu_4044_p2);

assign add_ln703_562_fu_4275_p2 = (sub_ln703_439_fu_4168_p2 + data_32_V_read_3_reg_9492_pp0_iter9_reg);

assign add_ln703_563_fu_4280_p2 = (sub_ln703_440_reg_11624 + data_32_V_read_3_reg_9492_pp0_iter9_reg);

assign add_ln703_564_fu_3947_p2 = (sub_ln703_347_fu_3400_p2 + data_26_V_read27_reg_9652_pp0_iter8_reg);

assign add_ln703_566_fu_3952_p2 = (add_ln703_466_reg_11410 + add_ln703_564_fu_3947_p2);

assign add_ln703_568_fu_3368_p2 = (data_32_V_read_3_reg_9492_pp0_iter7_reg + data_33_V_read_3_reg_9463_pp0_iter7_reg);

assign add_ln703_569_fu_3957_p2 = (add_ln703_568_reg_11464 + data_31_V_read32_reg_9521_pp0_iter8_reg);

assign add_ln703_570_fu_4294_p2 = (add_ln703_569_reg_11640 + add_ln703_507_reg_11441_pp0_iter9_reg);

assign add_ln703_571_fu_4298_p2 = (add_ln703_570_fu_4294_p2 + add_ln703_566_reg_11635);

assign add_ln703_572_fu_4308_p2 = (sub_ln703_446_fu_4197_p2 + data_33_V_read_3_reg_9463_pp0_iter9_reg);

assign add_ln703_573_fu_4323_p2 = (sub_ln703_450_fu_4221_p2 + data_33_V_read_3_reg_9463_pp0_iter9_reg);

assign add_ln703_574_fu_4566_p2 = (sub_ln703_453_reg_11683 + data_33_V_read_3_reg_9463_pp0_iter10_reg);

assign add_ln703_576_fu_4338_p2 = (add_ln703_568_reg_11464_pp0_iter9_reg + sub_ln703_433_fu_4129_p2);

assign add_ln703_577_fu_4343_p2 = (sub_ln703_406_fu_3981_p2 + data_30_V_read31_reg_9549_pp0_iter9_reg);

assign add_ln703_580_fu_4348_p2 = (add_ln703_569_reg_11640 + add_ln703_577_fu_4343_p2);

assign add_ln703_581_fu_4358_p2 = (sub_ln703_455_fu_4251_p2 + data_33_V_read_3_reg_9463_pp0_iter9_reg);

assign add_ln703_583_fu_4363_p2 = (add_ln703_568_reg_11464_pp0_iter9_reg + sub_ln703_435_fu_4144_p2);

assign add_ln703_585_fu_4383_p2 = (add_ln703_568_reg_11464_pp0_iter9_reg + sub_ln703_438_fu_4163_p2);

assign add_ln703_586_fu_4398_p2 = (sub_ln703_460_fu_4289_p2 + data_34_V_read_3_reg_9434_pp0_iter9_reg);

assign add_ln703_587_fu_4403_p2 = (sub_ln703_415_fu_4001_p2 + data_31_V_read32_reg_9521_pp0_iter9_reg);

assign add_ln703_588_fu_3961_p2 = (data_33_V_read_3_reg_9463_pp0_iter8_reg + data_34_V_read_3_reg_9434_pp0_iter8_reg);

assign add_ln703_589_fu_4408_p2 = (add_ln703_588_reg_11646 + data_32_V_read_3_reg_9492_pp0_iter9_reg);

assign add_ln703_590_fu_4412_p2 = (add_ln703_589_fu_4408_p2 + add_ln703_587_fu_4403_p2);

assign add_ln703_591_fu_4423_p2 = (sub_ln703_464_fu_4318_p2 + data_34_V_read_3_reg_9434_pp0_iter9_reg);

assign add_ln703_592_fu_4428_p2 = (sub_ln703_465_fu_4328_p2 + data_34_V_read_3_reg_9434_pp0_iter9_reg);

assign add_ln703_594_fu_4433_p2 = (add_ln703_507_reg_11441_pp0_iter9_reg + sub_ln703_390_reg_11499);

assign add_ln703_597_fu_4437_p2 = (add_ln703_588_reg_11646 + add_ln703_560_reg_11629);

assign add_ln703_598_fu_4441_p2 = (add_ln703_597_fu_4437_p2 + add_ln703_594_fu_4433_p2);

assign add_ln703_599_fu_4477_p2 = (sub_ln703_442_fu_4177_p2 + data_33_V_read_3_reg_9463_pp0_iter9_reg);

assign add_ln703_600_fu_3965_p2 = (data_34_V_read_3_reg_9434_pp0_iter8_reg + data_35_V_read_3_reg_9410_pp0_iter8_reg);

assign add_ln703_601_fu_4620_p2 = (add_ln703_600_reg_11652_pp0_iter10_reg + add_ln703_599_reg_11798);

assign add_ln703_602_fu_4482_p2 = (sub_ln703_384_reg_11474 + data_29_V_read_8_reg_9573_pp0_iter9_reg);

assign add_ln703_604_fu_4486_p2 = (add_ln703_534_reg_11248_pp0_iter9_reg + add_ln703_602_fu_4482_p2);

assign add_ln703_607_fu_4491_p2 = (add_ln703_600_reg_11652 + add_ln703_568_reg_11464_pp0_iter9_reg);

assign add_ln703_608_fu_4495_p2 = (add_ln703_607_fu_4491_p2 + add_ln703_604_fu_4486_p2);

assign add_ln703_609_fu_4501_p2 = (sub_ln703_444_fu_4187_p2 + data_33_V_read_3_reg_9463_pp0_iter9_reg);

assign add_ln703_611_fu_4628_p2 = (add_ln703_600_reg_11652_pp0_iter10_reg + add_ln703_609_reg_11803);

assign add_ln703_612_fu_4640_p2 = (sub_ln703_477_fu_4578_p2 + data_35_V_read_3_reg_9410_pp0_iter10_reg);

assign add_ln703_613_fu_4645_p2 = (sub_ln703_478_fu_4582_p2 + data_35_V_read_3_reg_9410_pp0_iter10_reg);

assign add_ln703_614_fu_4506_p2 = (sub_ln703_449_fu_4211_p2 + data_33_V_read_3_reg_9463_pp0_iter9_reg);

assign add_ln703_616_fu_4511_p2 = (add_ln703_600_reg_11652 + add_ln703_614_fu_4506_p2);

assign add_ln703_617_fu_4677_p2 = (sub_ln703_484_fu_4599_p2 + data_35_V_read_3_reg_9410_pp0_iter10_reg);

assign add_ln703_618_fu_4687_p2 = (sub_ln703_486_fu_4607_p2 + data_35_V_read_3_reg_9410_pp0_iter10_reg);

assign add_ln703_619_fu_4692_p2 = (sub_ln703_488_reg_11783 + data_35_V_read_3_reg_9410_pp0_iter10_reg);

assign add_ln703_620_fu_4696_p2 = (sub_ln703_491_reg_11793 + data_35_V_read_3_reg_9410_pp0_iter10_reg);

assign add_ln703_621_fu_3969_p2 = (data_35_V_read_3_reg_9410_pp0_iter8_reg + data_36_V_read_3_reg_9383_pp0_iter8_reg);

assign add_ln703_622_fu_4720_p2 = (add_ln703_621_reg_11662_pp0_iter10_reg + sub_ln703_476_fu_4574_p2);

assign add_ln703_623_fu_4739_p2 = (sub_ln703_496_fu_4650_p2 + data_36_V_read_3_reg_9383_pp0_iter10_reg);

assign add_ln703_624_fu_4754_p2 = (sub_ln703_466_fu_4562_p2 + data_34_V_read_3_reg_9434_pp0_iter10_reg);

assign add_ln703_626_fu_4759_p2 = (add_ln703_621_reg_11662_pp0_iter10_reg + add_ln703_624_fu_4754_p2);

assign add_ln703_627_fu_4769_p2 = (sub_ln703_501_fu_4672_p2 + data_36_V_read_3_reg_9383_pp0_iter10_reg);

assign add_ln703_629_fu_4774_p2 = (add_ln703_621_reg_11662_pp0_iter10_reg + sub_ln703_482_reg_11773);

assign add_ln703_631_fu_4526_p2 = (add_ln703_568_reg_11464_pp0_iter9_reg + sub_ln703_434_fu_4134_p2);

assign add_ln703_633_fu_4531_p2 = (add_ln703_621_reg_11662 + data_34_V_read_3_reg_9434_pp0_iter9_reg);

assign add_ln703_634_fu_4535_p2 = (add_ln703_633_fu_4531_p2 + add_ln703_631_fu_4526_p2);

assign add_ln703_636_fu_4793_p2 = (add_ln703_621_reg_11662_pp0_iter10_reg + sub_ln703_487_fu_4611_p2);

assign add_ln703_638_fu_4803_p2 = (add_ln703_621_reg_11662_pp0_iter10_reg + sub_ln703_489_fu_4615_p2);

assign add_ln703_639_fu_4541_p2 = (sub_ln703_459_fu_4284_p2 + data_33_V_read_3_reg_9463_pp0_iter9_reg);

assign add_ln703_642_fu_4817_p2 = (add_ln703_633_reg_11823 + add_ln703_639_reg_11833);

assign add_ln703_643_fu_4821_p2 = (sub_ln703_504_fu_4700_p2 + data_37_V_read_3_reg_9353_pp0_iter10_reg);

assign add_ln703_644_fu_4826_p2 = (sub_ln703_505_reg_11818 + data_37_V_read_3_reg_9353_pp0_iter10_reg);

assign add_ln703_645_fu_4835_p2 = (sub_ln703_507_fu_4710_p2 + data_37_V_read_3_reg_9353_pp0_iter10_reg);

assign add_ln703_646_fu_4546_p2 = (data_36_V_read_3_reg_9383_pp0_iter9_reg + data_37_V_read_3_reg_9353_pp0_iter9_reg);

assign add_ln703_647_fu_4870_p2 = (add_ln703_646_reg_11838 + sub_ln703_499_fu_4663_p2);

assign add_ln703_648_fu_4899_p2 = (sub_ln703_516_fu_4783_p2 + data_37_V_read_3_reg_9353_pp0_iter10_reg);

assign add_ln703_649_fu_4914_p2 = (sub_ln703_518_fu_4798_p2 + data_37_V_read_3_reg_9353_pp0_iter10_reg);

assign add_ln703_650_fu_4550_p2 = (data_37_V_read_3_reg_9353_pp0_iter9_reg + data_38_V_read_3_reg_9328_pp0_iter9_reg);

assign add_ln703_651_fu_4959_p2 = (add_ln703_650_reg_11844 + sub_ln703_510_fu_4730_p2);

assign add_ln703_653_fu_4964_p2 = (add_ln703_600_reg_11652_pp0_iter10_reg + sub_ln703_463_fu_4558_p2);

assign add_ln703_655_fu_4969_p2 = (add_ln703_650_reg_11844 + data_36_V_read_3_reg_9383_pp0_iter10_reg);

assign add_ln703_656_fu_4973_p2 = (add_ln703_655_fu_4969_p2 + add_ln703_653_fu_4964_p2);

assign add_ln703_658_fu_4989_p2 = (add_ln703_650_reg_11844 + sub_ln703_513_fu_4749_p2);

assign add_ln703_659_fu_5150_p2 = (sub_ln703_529_reg_11879 + data_38_V_read_3_reg_9328_pp0_iter11_reg);

assign add_ln703_660_fu_4994_p2 = (sub_ln703_531_fu_4890_p2 + data_38_V_read_3_reg_9328_pp0_iter10_reg);

assign add_ln703_661_fu_4999_p2 = (sub_ln703_534_fu_4909_p2 + data_38_V_read_3_reg_9328_pp0_iter10_reg);

assign add_ln703_662_fu_5166_p2 = (sub_ln703_535_reg_11899 + data_38_V_read_3_reg_9328_pp0_iter11_reg);

assign add_ln703_663_fu_5009_p2 = (sub_ln703_490_reg_11788 + data_35_V_read_3_reg_9410_pp0_iter10_reg);

assign add_ln703_666_fu_5013_p2 = (add_ln703_655_fu_4969_p2 + add_ln703_663_fu_5009_p2);

assign add_ln703_667_fu_4554_p2 = (data_38_V_read_3_reg_9328_pp0_iter9_reg + data_39_V_read_3_reg_9301_pp0_iter9_reg);

assign add_ln703_668_fu_5019_p2 = (add_ln703_667_reg_11853 + sub_ln703_521_fu_4830_p2);

assign add_ln703_669_fu_5186_p2 = (sub_ln703_544_reg_11934 + data_39_V_read_3_reg_9301_pp0_iter11_reg);

assign add_ln703_671_fu_5039_p2 = (add_ln703_667_reg_11853 + sub_ln703_530_fu_4885_p2);

assign add_ln703_673_fu_5044_p2 = (add_ln703_621_reg_11662_pp0_iter10_reg + sub_ln703_483_reg_11778);

assign add_ln703_675_fu_5048_p2 = (add_ln703_667_reg_11853 + data_37_V_read_3_reg_9353_pp0_iter10_reg);

assign add_ln703_676_fu_5052_p2 = (add_ln703_675_fu_5048_p2 + add_ln703_673_fu_5044_p2);

assign add_ln703_678_fu_5058_p2 = (add_ln703_600_reg_11652_pp0_iter10_reg + sub_ln703_469_reg_11733);

assign add_ln703_681_fu_5062_p2 = (add_ln703_667_reg_11853 + add_ln703_646_reg_11838);

assign add_ln703_682_fu_5066_p2 = (add_ln703_681_fu_5062_p2 + add_ln703_678_fu_5058_p2);

assign add_ln703_683_fu_5072_p2 = (sub_ln703_519_fu_4808_p2 + data_37_V_read_3_reg_9353_pp0_iter10_reg);

assign add_ln703_685_fu_5077_p2 = (add_ln703_667_reg_11853 + add_ln703_683_fu_5072_p2);

assign add_ln703_687_fu_5082_p2 = (add_ln703_667_reg_11853 + sub_ln703_536_fu_4924_p2);

assign add_ln703_689_fu_5087_p2 = (add_ln703_667_reg_11853 + sub_ln703_537_fu_4929_p2);

assign add_ln703_690_fu_5240_p2 = (sub_ln703_553_fu_5174_p2 + data_40_V_read41_reg_9272_pp0_iter11_reg);

assign add_ln703_691_fu_5092_p2 = (data_39_V_read_3_reg_9301_pp0_iter10_reg + data_40_V_read41_reg_9272_pp0_iter10_reg);

assign add_ln703_692_fu_5245_p2 = (add_ln703_691_reg_11994 + sub_ln703_541_reg_11919);

assign add_ln703_693_fu_5249_p2 = (sub_ln703_554_fu_5178_p2 + data_40_V_read41_reg_9272_pp0_iter11_reg);

assign add_ln703_694_fu_5254_p2 = (sub_ln703_555_fu_5182_p2 + data_40_V_read41_reg_9272_pp0_iter11_reg);

assign add_ln703_695_fu_5259_p2 = (sub_ln703_556_reg_11964 + data_40_V_read41_reg_9272_pp0_iter11_reg);

assign add_ln703_696_fu_5272_p2 = (sub_ln703_558_reg_11974 + data_40_V_read41_reg_9272_pp0_iter11_reg);

assign add_ln703_697_fu_5096_p2 = (sub_ln703_528_fu_4875_p2 + data_38_V_read_3_reg_9328_pp0_iter10_reg);

assign add_ln703_699_fu_5281_p2 = (add_ln703_691_reg_11994 + add_ln703_697_reg_12002);

assign add_ln703_700_fu_5285_p2 = (sub_ln703_561_fu_5200_p2 + data_40_V_read41_reg_9272_pp0_iter11_reg);

assign add_ln703_701_fu_5313_p2 = (sub_ln703_566_fu_5223_p2 + data_40_V_read41_reg_9272_pp0_iter11_reg);

assign add_ln703_702_fu_5332_p2 = (sub_ln703_538_reg_11904 + data_39_V_read_3_reg_9301_pp0_iter11_reg);

assign add_ln703_703_fu_5116_p2 = (data_40_V_read41_reg_9272_pp0_iter10_reg + data_41_V_read42_reg_9242_pp0_iter10_reg);

assign add_ln703_704_fu_5336_p2 = (add_ln703_703_reg_12022 + add_ln703_702_fu_5332_p2);

assign add_ln703_706_fu_5120_p2 = (add_ln703_650_reg_11844 + sub_ln703_509_fu_4725_p2);

assign add_ln703_708_fu_5361_p2 = (add_ln703_703_reg_12022 + data_39_V_read_3_reg_9301_pp0_iter11_reg);

assign add_ln703_709_fu_5365_p2 = (add_ln703_708_fu_5361_p2 + add_ln703_706_reg_12031);

assign add_ln703_710_fu_5390_p2 = (sub_ln703_545_fu_5138_p2 + data_39_V_read_3_reg_9301_pp0_iter11_reg);

assign add_ln703_712_fu_5395_p2 = (add_ln703_703_reg_12022 + add_ln703_710_fu_5390_p2);

assign add_ln703_714_fu_5405_p2 = (add_ln703_703_reg_12022 + sub_ln703_559_fu_5190_p2);

assign add_ln703_715_fu_5425_p2 = (sub_ln703_573_reg_12007 + data_41_V_read42_reg_9242_pp0_iter11_reg);

assign add_ln703_716_fu_5429_p2 = (sub_ln703_574_fu_5290_p2 + data_41_V_read42_reg_9242_pp0_iter11_reg);

assign add_ln703_718_fu_5434_p2 = (add_ln703_703_reg_12022 + sub_ln703_563_fu_5209_p2);

assign add_ln703_719_fu_5439_p2 = (sub_ln703_576_fu_5299_p2 + data_41_V_read42_reg_9242_pp0_iter11_reg);

assign add_ln703_720_fu_5469_p2 = (sub_ln703_582_reg_12012 + data_41_V_read42_reg_9242_pp0_iter11_reg);

assign add_ln703_721_fu_5692_p2 = (sub_ln703_586_reg_12061 + data_42_V_read_3_reg_9212_pp0_iter12_reg);

assign add_ln703_722_fu_5125_p2 = (sub_ln703_495_fu_4636_p2 + data_36_V_read_3_reg_9383_pp0_iter10_reg);

assign add_ln703_724_fu_5477_p2 = (add_ln703_650_reg_11844_pp0_iter11_reg + add_ln703_722_reg_12036);

assign add_ln703_726_fu_5130_p2 = (data_41_V_read42_reg_9242_pp0_iter10_reg + data_42_V_read_3_reg_9212_pp0_iter10_reg);

assign add_ln703_727_fu_5481_p2 = (add_ln703_726_reg_12041 + add_ln703_691_reg_11994);

assign add_ln703_728_fu_5485_p2 = (add_ln703_727_fu_5481_p2 + add_ln703_724_fu_5477_p2);

assign add_ln703_729_fu_5700_p2 = (sub_ln703_593_reg_12071 + data_42_V_read_3_reg_9212_pp0_iter12_reg);

assign add_ln703_730_fu_5541_p2 = (sub_ln703_596_fu_5444_p2 + data_42_V_read_3_reg_9212_pp0_iter11_reg);

assign add_ln703_732_fu_5546_p2 = (add_ln703_726_reg_12041 + sub_ln703_578_fu_5308_p2);

assign add_ln703_733_fu_5551_p2 = (sub_ln703_597_fu_5449_p2 + data_42_V_read_3_reg_9212_pp0_iter11_reg);

assign add_ln703_734_fu_5556_p2 = (sub_ln703_599_fu_5459_p2 + data_42_V_read_3_reg_9212_pp0_iter11_reg);

assign add_ln703_735_fu_5571_p2 = (sub_ln703_601_fu_5473_p2 + data_42_V_read_3_reg_9212_pp0_iter11_reg);

assign add_ln703_736_fu_5576_p2 = (sub_ln703_552_fu_5170_p2 + data_40_V_read41_reg_9272_pp0_iter11_reg);

assign add_ln703_737_fu_5134_p2 = (data_42_V_read_3_reg_9212_pp0_iter10_reg + data_43_V_read_3_reg_9184_pp0_iter10_reg);

assign add_ln703_738_fu_5581_p2 = (add_ln703_737_reg_12047 + data_41_V_read42_reg_9242_pp0_iter11_reg);

assign add_ln703_739_fu_5585_p2 = (add_ln703_738_fu_5581_p2 + add_ln703_736_fu_5576_p2);

assign add_ln703_741_fu_5591_p2 = (add_ln703_737_reg_12047 + sub_ln703_584_fu_5341_p2);

assign add_ln703_742_fu_5738_p2 = (sub_ln703_605_reg_12111 + data_43_V_read_3_reg_9184_pp0_iter12_reg);

assign add_ln703_744_fu_5601_p2 = (add_ln703_737_reg_12047 + sub_ln703_592_fu_5400_p2);

assign add_ln703_745_fu_5606_p2 = (sub_ln703_575_fu_5295_p2 + data_41_V_read42_reg_9242_pp0_iter11_reg);

assign add_ln703_747_fu_5611_p2 = (add_ln703_737_reg_12047 + add_ln703_745_fu_5606_p2);

assign add_ln703_748_fu_5759_p2 = (sub_ln703_614_reg_12141 + data_43_V_read_3_reg_9184_pp0_iter12_reg);

assign add_ln703_750_fu_5616_p2 = (add_ln703_691_reg_11994 + sub_ln703_549_fu_5158_p2);

assign add_ln703_753_fu_5621_p2 = (add_ln703_738_fu_5581_p2 + add_ln703_750_fu_5616_p2);

assign add_ln703_754_fu_5776_p2 = (sub_ln703_618_reg_12156 + data_43_V_read_3_reg_9184_pp0_iter12_reg);

assign add_ln703_755_fu_5652_p2 = (data_43_V_read_3_reg_9184_pp0_iter11_reg + data_44_V_read_3_reg_9154_pp0_iter11_reg);

assign add_ln703_756_fu_5809_p2 = (add_ln703_755_reg_12196 + sub_ln703_606_fu_5696_p2);

assign add_ln703_757_fu_5814_p2 = (sub_ln703_624_reg_12166 + data_44_V_read_3_reg_9154_pp0_iter12_reg);

assign add_ln703_759_fu_5818_p2 = (add_ln703_755_reg_12196 + sub_ln703_608_reg_12116);

assign add_ln703_761_fu_5837_p2 = (add_ln703_755_reg_12196 + sub_ln703_611_fu_5704_p2);

assign add_ln703_763_fu_5842_p2 = (add_ln703_755_reg_12196 + sub_ln703_612_reg_12131);

assign add_ln703_764_fu_5861_p2 = (sub_ln703_630_reg_12171 + data_44_V_read_3_reg_9154_pp0_iter12_reg);

assign add_ln703_765_fu_5671_p2 = (data_44_V_read_3_reg_9154_pp0_iter11_reg + data_45_V_read_3_reg_9125_pp0_iter11_reg);

assign add_ln703_766_fu_5893_p2 = (add_ln703_765_reg_12219 + sub_ln703_621_fu_5726_p2);

assign add_ln703_767_fu_5942_p2 = (sub_ln703_595_reg_12081 + data_42_V_read_3_reg_9212_pp0_iter12_reg);

assign add_ln703_769_fu_5946_p2 = (add_ln703_765_reg_12219 + data_43_V_read_3_reg_9184_pp0_iter12_reg);

assign add_ln703_770_fu_5950_p2 = (add_ln703_769_fu_5946_p2 + add_ln703_767_fu_5942_p2);

assign add_ln703_771_fu_5961_p2 = (sub_ln703_647_fu_5846_p2 + data_45_V_read_3_reg_9125_pp0_iter12_reg);

assign add_ln703_772_fu_5966_p2 = (sub_ln703_649_fu_5851_p2 + data_45_V_read_3_reg_9125_pp0_iter12_reg);

assign add_ln703_774_fu_5985_p2 = (add_ln703_765_reg_12219 + sub_ln703_631_reg_12176);

assign add_ln703_775_fu_5994_p2 = (sub_ln703_616_fu_5712_p2 + data_43_V_read_3_reg_9184_pp0_iter12_reg);

assign add_ln703_777_fu_5999_p2 = (add_ln703_765_reg_12219 + add_ln703_775_fu_5994_p2);

assign add_ln703_778_fu_5675_p2 = (data_45_V_read_3_reg_9125_pp0_iter11_reg + data_46_V_read_3_reg_9094_pp0_iter11_reg);

assign add_ln703_779_fu_6024_p2 = (add_ln703_778_reg_12227 + sub_ln703_636_fu_5784_p2);

assign add_ln703_781_fu_6029_p2 = (add_ln703_778_reg_12227 + sub_ln703_637_reg_12186);

assign add_ln703_783_fu_5679_p2 = (add_ln703_737_reg_12047 + sub_ln703_585_fu_5346_p2);

assign add_ln703_785_fu_6038_p2 = (add_ln703_778_reg_12227 + data_44_V_read_3_reg_9154_pp0_iter12_reg);

assign add_ln703_786_fu_6042_p2 = (add_ln703_785_fu_6038_p2 + add_ln703_783_reg_12236);

assign add_ln703_788_fu_6082_p2 = (add_ln703_778_reg_12227 + sub_ln703_648_reg_12209);

assign add_ln703_789_fu_6250_p2 = (sub_ln703_669_reg_12268 + data_46_V_read_3_reg_9094_pp0_iter13_reg);

assign add_ln703_790_fu_6121_p2 = (sub_ln703_673_fu_6009_p2 + data_46_V_read_3_reg_9094_pp0_iter12_reg);

assign add_ln703_791_fu_6131_p2 = (sub_ln703_675_fu_6019_p2 + data_46_V_read_3_reg_9094_pp0_iter12_reg);

assign add_ln703_792_fu_6146_p2 = (sub_ln703_677_fu_6047_p2 + data_47_V_read_3_reg_9066_pp0_iter12_reg);

assign add_ln703_793_fu_6258_p2 = (sub_ln703_678_reg_12283 + data_47_V_read_3_reg_9066_pp0_iter13_reg);

assign add_ln703_794_fu_6151_p2 = (sub_ln703_641_fu_5799_p2 + data_45_V_read_3_reg_9125_pp0_iter12_reg);

assign add_ln703_795_fu_6156_p2 = (data_46_V_read_3_reg_9094_pp0_iter12_reg + data_47_V_read_3_reg_9066_pp0_iter12_reg);

assign add_ln703_796_fu_6160_p2 = (add_ln703_795_fu_6156_p2 + add_ln703_794_fu_6151_p2);

assign add_ln703_797_fu_6262_p2 = (sub_ln703_681_fu_6238_p2 + data_47_V_read_3_reg_9066_pp0_iter13_reg);

assign add_ln703_798_fu_6166_p2 = (add_ln703_795_fu_6156_p2 + sub_ln703_663_fu_5923_p2);

assign add_ln703_799_fu_6276_p2 = (sub_ln703_685_fu_6246_p2 + data_47_V_read_3_reg_9066_pp0_iter13_reg);

assign add_ln703_800_fu_6315_p2 = (sub_ln703_697_reg_12358 + data_48_V_read_3_reg_9040_pp0_iter13_reg);

assign add_ln703_801_fu_6187_p2 = (sub_ln703_639_fu_5789_p2 + data_45_V_read_3_reg_9125_pp0_iter12_reg);

assign add_ln703_802_fu_6192_p2 = (data_47_V_read_3_reg_9066_pp0_iter12_reg + data_48_V_read_3_reg_9040_pp0_iter12_reg);

assign add_ln703_803_fu_6319_p2 = (add_ln703_802_reg_12398 + data_46_V_read_3_reg_9094_pp0_iter13_reg);

assign add_ln703_804_fu_6323_p2 = (add_ln703_803_fu_6319_p2 + add_ln703_801_reg_12393);

assign add_ln703_805_fu_6341_p2 = (add_ln703_802_reg_12398 + sub_ln703_680_reg_12293);

assign add_ln703_806_fu_6359_p2 = (sub_ln703_699_fu_6271_p2 + data_48_V_read_3_reg_9040_pp0_iter13_reg);

assign add_ln703_807_fu_6369_p2 = (sub_ln703_667_reg_12263 + data_46_V_read_3_reg_9094_pp0_iter13_reg);

assign add_ln703_808_fu_6373_p2 = (add_ln703_802_reg_12398 + add_ln703_807_fu_6369_p2);

assign add_ln703_809_fu_6378_p2 = (add_ln703_802_reg_12398 + sub_ln703_686_reg_12308);

assign add_ln703_810_fu_6396_p2 = (sub_ln703_703_fu_6289_p2 + data_48_V_read_3_reg_9040_pp0_iter13_reg);

assign add_ln703_811_fu_6401_p2 = (sub_ln703_704_reg_12383 + data_48_V_read_3_reg_9040_pp0_iter13_reg);

assign add_ln703_812_fu_6405_p2 = (add_ln703_802_reg_12398 + sub_ln703_690_reg_12323);

assign add_ln703_813_fu_6409_p2 = (add_ln703_802_reg_12398 + sub_ln703_692_reg_12333);

assign add_ln703_814_fu_6417_p2 = (sub_ln703_708_fu_6302_p2 + data_48_V_read_3_reg_9040_pp0_iter13_reg);

assign add_ln703_815_fu_6196_p2 = (sub_ln703_661_fu_5913_p2 + data_46_V_read_3_reg_9094_pp0_iter12_reg);

assign add_ln703_816_fu_5684_p2 = (data_48_V_read_3_reg_9040_pp0_iter11_reg + data_49_V_read_3_reg_9012_pp0_iter11_reg);

assign add_ln703_817_fu_6201_p2 = (add_ln703_816_reg_12241 + data_47_V_read_3_reg_9066_pp0_iter12_reg);

assign add_ln703_818_fu_6205_p2 = (add_ln703_817_fu_6201_p2 + add_ln703_815_fu_6196_p2);

assign add_ln703_819_fu_6447_p2 = (sub_ln703_714_fu_6345_p2 + data_49_V_read_3_reg_9012_pp0_iter13_reg);

assign add_ln703_820_fu_6211_p2 = (add_ln703_778_reg_12227 + sub_ln703_645_fu_5827_p2);

assign add_ln703_821_fu_6216_p2 = (add_ln703_817_fu_6201_p2 + add_ln703_820_fu_6211_p2);

assign add_ln703_822_fu_6482_p2 = (sub_ln703_720_fu_6391_p2 + data_49_V_read_3_reg_9012_pp0_iter13_reg);

assign add_ln703_823_fu_6512_p2 = (sub_ln703_694_reg_12343 + data_47_V_read_3_reg_9066_pp0_iter13_reg);

assign add_ln703_824_fu_6516_p2 = (add_ln703_816_reg_12241_pp0_iter13_reg + add_ln703_823_fu_6512_p2);

assign add_ln703_825_fu_6526_p2 = (sub_ln703_722_fu_6422_p2 + data_50_V_read51_reg_8984_pp0_iter13_reg);

assign add_ln703_826_fu_6222_p2 = (data_49_V_read_3_reg_9012_pp0_iter12_reg + data_50_V_read51_reg_8984_pp0_iter12_reg);

assign add_ln703_827_fu_6531_p2 = (add_ln703_826_reg_12419 + sub_ln703_710_fu_6311_p2);

assign add_ln703_828_fu_6536_p2 = (add_ln703_826_reg_12419 + sub_ln703_712_fu_6332_p2);

assign add_ln703_829_fu_6546_p2 = (sub_ln703_679_reg_12288 + data_47_V_read_3_reg_9066_pp0_iter13_reg);

assign add_ln703_830_fu_6550_p2 = (add_ln703_826_reg_12419 + data_48_V_read_3_reg_9040_pp0_iter13_reg);

assign add_ln703_831_fu_6554_p2 = (add_ln703_830_fu_6550_p2 + add_ln703_829_fu_6546_p2);

assign add_ln703_832_fu_6569_p2 = (sub_ln703_684_reg_12303 + data_47_V_read_3_reg_9066_pp0_iter13_reg);

assign add_ln703_833_fu_6573_p2 = (add_ln703_830_fu_6550_p2 + add_ln703_832_fu_6569_p2);

assign add_ln703_834_fu_6594_p2 = (sub_ln703_732_fu_6477_p2 + data_50_V_read51_reg_8984_pp0_iter13_reg);

assign add_ln703_835_fu_6815_p2 = (sub_ln703_736_reg_12475 + data_50_V_read51_reg_8984_pp0_iter14_reg);

assign add_ln703_836_fu_6226_p2 = (data_50_V_read51_reg_8984_pp0_iter12_reg + data_51_V_read52_reg_8956_pp0_iter12_reg);

assign add_ln703_837_fu_6624_p2 = (add_ln703_836_reg_12428 + sub_ln703_723_fu_6427_p2);

assign add_ln703_838_fu_6634_p2 = (sub_ln703_739_fu_6541_p2 + data_51_V_read52_reg_8956_pp0_iter13_reg);

assign add_ln703_839_fu_6836_p2 = (sub_ln703_743_fu_6803_p2 + data_51_V_read52_reg_8956_pp0_iter14_reg);

assign add_ln703_840_fu_6649_p2 = (sub_ln703_747_fu_6584_p2 + data_51_V_read52_reg_8956_pp0_iter13_reg);

assign add_ln703_841_fu_6664_p2 = (sub_ln703_752_fu_6609_p2 + data_51_V_read52_reg_8956_pp0_iter13_reg);

assign add_ln703_842_fu_6669_p2 = (sub_ln703_705_fu_6294_p2 + data_48_V_read_3_reg_9040_pp0_iter13_reg);

assign add_ln703_843_fu_6674_p2 = (add_ln703_836_reg_12428 + data_49_V_read_3_reg_9012_pp0_iter13_reg);

assign add_ln703_844_fu_6678_p2 = (add_ln703_843_fu_6674_p2 + add_ln703_842_fu_6669_p2);

assign add_ln703_845_fu_6689_p2 = (sub_ln703_754_fu_6619_p2 + data_51_V_read52_reg_8956_pp0_iter13_reg);

assign add_ln703_846_fu_6863_p2 = (sub_ln703_755_fu_6819_p2 + data_52_V_read_3_reg_8928_pp0_iter14_reg);

assign add_ln703_847_fu_6868_p2 = (sub_ln703_756_fu_6823_p2 + data_52_V_read_3_reg_8928_pp0_iter14_reg);

assign add_ln703_848_fu_6694_p2 = (add_ln703_802_reg_12398 + sub_ln703_676_reg_12278);

assign add_ln703_849_fu_6230_p2 = (data_51_V_read52_reg_8956_pp0_iter12_reg + data_52_V_read_3_reg_8928_pp0_iter12_reg);

assign add_ln703_850_fu_6698_p2 = (add_ln703_849_reg_12434 + add_ln703_826_reg_12419);

assign add_ln703_851_fu_6702_p2 = (add_ln703_850_fu_6698_p2 + add_ln703_848_fu_6694_p2);

assign add_ln703_852_fu_6713_p2 = (sub_ln703_711_fu_6328_p2 + data_49_V_read_3_reg_9012_pp0_iter13_reg);

assign add_ln703_853_fu_6718_p2 = (add_ln703_849_reg_12434 + data_50_V_read51_reg_8984_pp0_iter13_reg);

assign add_ln703_854_fu_6722_p2 = (add_ln703_853_fu_6718_p2 + add_ln703_852_fu_6713_p2);

assign add_ln703_855_fu_6882_p2 = (sub_ln703_759_reg_12525 + data_52_V_read_3_reg_8928_pp0_iter14_reg);

assign add_ln703_856_fu_6891_p2 = (add_ln703_849_reg_12434_pp0_iter14_reg + sub_ln703_742_fu_6799_p2);

assign add_ln703_857_fu_6728_p2 = (sub_ln703_716_fu_6354_p2 + data_49_V_read_3_reg_9012_pp0_iter13_reg);

assign add_ln703_858_fu_6733_p2 = (add_ln703_853_fu_6718_p2 + add_ln703_857_fu_6728_p2);

assign add_ln703_859_fu_6901_p2 = (sub_ln703_761_reg_12530 + data_52_V_read_3_reg_8928_pp0_iter14_reg);

assign add_ln703_860_fu_6905_p2 = (add_ln703_849_reg_12434_pp0_iter14_reg + sub_ln703_745_fu_6807_p2);

assign add_ln703_861_fu_6919_p2 = (sub_ln703_763_reg_12540 + data_52_V_read_3_reg_8928_pp0_iter14_reg);

assign add_ln703_862_fu_6923_p2 = (sub_ln703_764_fu_6845_p2 + data_52_V_read_3_reg_8928_pp0_iter14_reg);

assign add_ln703_863_fu_6744_p2 = (add_ln703_816_reg_12241_pp0_iter13_reg + sub_ln703_706_fu_6298_p2);

assign add_ln703_864_fu_6749_p2 = (add_ln703_853_fu_6718_p2 + add_ln703_863_fu_6744_p2);

assign add_ln703_865_fu_6968_p2 = (sub_ln703_770_reg_12570 + data_53_V_read_3_reg_8899_pp0_iter14_reg);

assign add_ln703_866_fu_6972_p2 = (sub_ln703_724_reg_12450 + data_50_V_read51_reg_8984_pp0_iter14_reg);

assign add_ln703_867_fu_6234_p2 = (data_52_V_read_3_reg_8928_pp0_iter12_reg + data_53_V_read_3_reg_8899_pp0_iter12_reg);

assign add_ln703_868_fu_6755_p2 = (add_ln703_867_reg_12444 + data_51_V_read52_reg_8956_pp0_iter13_reg);

assign add_ln703_869_fu_6976_p2 = (add_ln703_868_reg_12585 + add_ln703_866_fu_6972_p2);

assign add_ln703_870_fu_7025_p2 = (sub_ln703_777_fu_6928_p2 + data_53_V_read_3_reg_8899_pp0_iter14_reg);

assign add_ln703_871_fu_7040_p2 = (sub_ln703_782_fu_6946_p2 + data_53_V_read_3_reg_8899_pp0_iter14_reg);

assign add_ln703_872_fu_7050_p2 = (sub_ln703_784_fu_6954_p2 + data_54_V_read_3_reg_8873_pp0_iter14_reg);

assign add_ln703_873_fu_7055_p2 = (sub_ln703_785_fu_6959_p2 + data_54_V_read_3_reg_8873_pp0_iter14_reg);

assign add_ln703_874_fu_7084_p2 = (sub_ln703_791_fu_6996_p2 + data_54_V_read_3_reg_8873_pp0_iter14_reg);

assign add_ln703_875_fu_7094_p2 = (sub_ln703_793_fu_7005_p2 + data_54_V_read_3_reg_8873_pp0_iter14_reg);

assign add_ln703_876_fu_6769_p2 = (add_ln703_826_reg_12419 + sub_ln703_717_fu_6364_p2);

assign add_ln703_877_fu_6774_p2 = (data_53_V_read_3_reg_8899_pp0_iter13_reg + data_54_V_read_3_reg_8873_pp0_iter13_reg);

assign add_ln703_878_fu_7104_p2 = (add_ln703_877_reg_12605 + add_ln703_849_reg_12434_pp0_iter14_reg);

assign add_ln703_879_fu_7108_p2 = (add_ln703_878_fu_7104_p2 + add_ln703_876_reg_12600);

assign add_ln703_880_fu_7113_p2 = (sub_ln703_746_reg_12500 + data_51_V_read52_reg_8956_pp0_iter14_reg);

assign add_ln703_881_fu_7117_p2 = (add_ln703_877_reg_12605 + data_52_V_read_3_reg_8928_pp0_iter14_reg);

assign add_ln703_882_fu_7121_p2 = (add_ln703_881_fu_7117_p2 + add_ln703_880_fu_7113_p2);

assign add_ln703_883_fu_7127_p2 = (sub_ln703_795_fu_7015_p2 + data_54_V_read_3_reg_8873_pp0_iter14_reg);

assign add_ln703_884_fu_7132_p2 = (sub_ln703_796_fu_7020_p2 + data_54_V_read_3_reg_8873_pp0_iter14_reg);

assign add_ln703_885_fu_7142_p2 = (sub_ln703_798_fu_7035_p2 + data_54_V_read_3_reg_8873_pp0_iter14_reg);

assign add_ln703_886_fu_7147_p2 = (add_ln703_877_reg_12605 + sub_ln703_781_reg_12580);

assign add_ln703_887_fu_7151_p2 = (sub_ln703_768_fu_6858_p2 + data_52_V_read_3_reg_8928_pp0_iter14_reg);

assign add_ln703_888_fu_7156_p2 = (add_ln703_877_reg_12605 + add_ln703_887_fu_7151_p2);

assign add_ln703_889_fu_7161_p2 = (sub_ln703_799_reg_12595 + data_54_V_read_3_reg_8873_pp0_iter14_reg);

assign add_ln703_890_fu_7354_p2 = (sub_ln703_801_reg_12660 + data_55_V_read_3_reg_8844_pp0_iter15_reg);

assign add_ln703_891_fu_7358_p2 = (sub_ln703_802_reg_12665 + data_55_V_read_3_reg_8844_pp0_iter15_reg);

assign add_ln703_892_fu_7175_p2 = (sub_ln703_803_fu_7070_p2 + data_55_V_read_3_reg_8844_pp0_iter14_reg);

assign add_ln703_893_fu_7180_p2 = (sub_ln703_804_fu_7075_p2 + data_55_V_read_3_reg_8844_pp0_iter14_reg);

assign add_ln703_894_fu_6778_p2 = (data_54_V_read_3_reg_8873_pp0_iter13_reg + data_55_V_read_3_reg_8844_pp0_iter13_reg);

assign add_ln703_895_fu_7185_p2 = (add_ln703_894_reg_12616 + sub_ln703_788_fu_6981_p2);

assign add_ln703_896_fu_7190_p2 = (sub_ln703_773_fu_6886_p2 + data_53_V_read_3_reg_8899_pp0_iter14_reg);

assign add_ln703_897_fu_7362_p2 = (add_ln703_894_reg_12616_pp0_iter15_reg + add_ln703_896_reg_12725);

assign add_ln703_898_fu_7195_p2 = (sub_ln703_774_fu_6896_p2 + data_53_V_read_3_reg_8899_pp0_iter14_reg);

assign add_ln703_899_fu_7366_p2 = (add_ln703_894_reg_12616_pp0_iter15_reg + add_ln703_898_reg_12730);

assign add_ln703_900_fu_7378_p2 = (sub_ln703_807_reg_12685 + data_55_V_read_3_reg_8844_pp0_iter15_reg);

assign add_ln703_901_fu_7390_p2 = (sub_ln703_808_reg_12700 + data_55_V_read_3_reg_8844_pp0_iter15_reg);

assign add_ln703_902_fu_7394_p2 = (add_ln703_894_reg_12616_pp0_iter15_reg + sub_ln703_797_reg_12645);

assign add_ln703_903_fu_7402_p2 = (sub_ln703_811_fu_7346_p2 + data_56_V_read_3_reg_8814_pp0_iter15_reg);

assign add_ln703_904_fu_7240_p2 = (sub_ln703_789_fu_6986_p2 + data_54_V_read_3_reg_8873_pp0_iter14_reg);

assign add_ln703_905_fu_6782_p2 = (data_55_V_read_3_reg_8844_pp0_iter13_reg + data_56_V_read_3_reg_8814_pp0_iter13_reg);

assign add_ln703_906_fu_7245_p2 = (add_ln703_905_reg_12625 + add_ln703_904_fu_7240_p2);

assign add_ln703_907_fu_7477_p2 = (sub_ln703_820_reg_12750 + data_56_V_read_3_reg_8814_pp0_iter15_reg);

assign add_ln703_908_fu_7250_p2 = (sub_ln703_780_fu_6942_p2 + data_53_V_read_3_reg_8899_pp0_iter14_reg);

assign add_ln703_909_fu_7255_p2 = (add_ln703_905_reg_12625 + data_54_V_read_3_reg_8873_pp0_iter14_reg);

assign add_ln703_910_fu_7259_p2 = (add_ln703_909_fu_7255_p2 + add_ln703_908_fu_7250_p2);

assign add_ln703_911_fu_7481_p2 = (sub_ln703_821_reg_12755 + data_56_V_read_3_reg_8814_pp0_iter15_reg);

assign add_ln703_912_fu_7490_p2 = (sub_ln703_824_reg_12765 + data_56_V_read_3_reg_8814_pp0_iter15_reg);

assign add_ln703_913_fu_7494_p2 = (sub_ln703_825_reg_12770 + data_56_V_read_3_reg_8814_pp0_iter15_reg);

assign add_ln703_914_fu_6786_p2 = (sub_ln703_738_fu_6521_p2 + data_50_V_read51_reg_8984_pp0_iter13_reg);

assign add_ln703_915_fu_7265_p2 = (add_ln703_849_reg_12434_pp0_iter14_reg + add_ln703_914_reg_12632);

assign add_ln703_916_fu_7269_p2 = (add_ln703_905_reg_12625 + add_ln703_877_reg_12605);

assign add_ln703_917_fu_7273_p2 = (add_ln703_916_fu_7269_p2 + add_ln703_915_fu_7265_p2);

assign add_ln703_918_fu_7513_p2 = (sub_ln703_828_fu_7417_p2 + data_57_V_read_3_reg_8786_pp0_iter15_reg);

assign add_ln703_919_fu_7279_p2 = (add_ln703_867_reg_12444_pp0_iter14_reg + sub_ln703_757_reg_12515);

assign add_ln703_920_fu_6791_p2 = (data_56_V_read_3_reg_8814_pp0_iter13_reg + data_57_V_read_3_reg_8786_pp0_iter13_reg);

assign add_ln703_921_fu_7283_p2 = (add_ln703_920_reg_12637 + add_ln703_894_reg_12616);

assign add_ln703_922_fu_7287_p2 = (add_ln703_921_fu_7283_p2 + add_ln703_919_fu_7279_p2);

assign add_ln703_923_fu_7293_p2 = (add_ln703_877_reg_12605 + sub_ln703_771_fu_6873_p2);

assign add_ln703_924_fu_7298_p2 = (add_ln703_920_reg_12637 + data_55_V_read_3_reg_8844_pp0_iter14_reg);

assign add_ln703_925_fu_7302_p2 = (add_ln703_924_fu_7298_p2 + add_ln703_923_fu_7293_p2);

assign add_ln703_926_fu_7532_p2 = (sub_ln703_832_fu_7434_p2 + data_57_V_read_3_reg_8786_pp0_iter15_reg);

assign add_ln703_927_fu_7537_p2 = (sub_ln703_805_reg_12670 + data_55_V_read_3_reg_8844_pp0_iter15_reg);

assign add_ln703_928_fu_7541_p2 = (add_ln703_920_reg_12637_pp0_iter15_reg + add_ln703_927_fu_7537_p2);

assign add_ln703_929_fu_7546_p2 = (sub_ln703_833_fu_7439_p2 + data_57_V_read_3_reg_8786_pp0_iter15_reg);

assign add_ln703_930_fu_7561_p2 = (sub_ln703_837_fu_7458_p2 + data_57_V_read_3_reg_8786_pp0_iter15_reg);

assign add_ln703_931_fu_7308_p2 = (add_ln703_877_reg_12605 + sub_ln703_776_fu_6915_p2);

assign add_ln703_932_fu_7313_p2 = (add_ln703_924_fu_7298_p2 + add_ln703_931_fu_7308_p2);

assign add_ln703_933_fu_7581_p2 = (sub_ln703_841_fu_7485_p2 + data_57_V_read_3_reg_8786_pp0_iter15_reg);

assign add_ln703_934_fu_7610_p2 = (sub_ln703_844_fu_7508_p2 + data_58_V_read_3_reg_8756_pp0_iter15_reg);

assign add_ln703_935_fu_7629_p2 = (sub_ln703_846_fu_7523_p2 + data_58_V_read_3_reg_8756_pp0_iter15_reg);

assign add_ln703_936_fu_7634_p2 = (sub_ln703_847_fu_7528_p2 + data_58_V_read_3_reg_8756_pp0_iter15_reg);

assign add_ln703_937_fu_7659_p2 = (data_57_V_read_3_reg_8786_pp0_iter15_reg + data_58_V_read_3_reg_8756_pp0_iter15_reg);

assign add_ln703_938_fu_7663_p2 = (add_ln703_937_fu_7659_p2 + sub_ln703_835_fu_7449_p2);

assign add_ln703_939_fu_7679_p2 = (add_ln703_937_fu_7659_p2 + sub_ln703_838_fu_7463_p2);

assign add_ln703_940_fu_7690_p2 = (add_ln703_937_fu_7659_p2 + sub_ln703_840_fu_7472_p2);

assign add_ln703_941_fu_7701_p2 = (sub_ln703_852_reg_12790 + data_58_V_read_3_reg_8756_pp0_iter15_reg);

assign add_ln703_942_fu_7715_p2 = (sub_ln703_823_reg_12760 + data_56_V_read_3_reg_8814_pp0_iter15_reg);

assign add_ln703_943_fu_7719_p2 = (add_ln703_937_fu_7659_p2 + add_ln703_942_fu_7715_p2);

assign add_ln703_944_fu_7882_p2 = (sub_ln703_858_reg_12840 + data_59_V_read_3_reg_8724_pp0_iter16_reg);

assign add_ln703_945_fu_7740_p2 = (sub_ln703_830_fu_7426_p2 + data_57_V_read_3_reg_8786_pp0_iter15_reg);

assign add_ln703_946_fu_7334_p2 = (data_58_V_read_3_reg_8756_pp0_iter14_reg + data_59_V_read_3_reg_8724_pp0_iter14_reg);

assign add_ln703_947_fu_7745_p2 = (add_ln703_946_reg_12805 + add_ln703_945_fu_7740_p2);

assign add_ln703_948_fu_7760_p2 = (sub_ln703_864_fu_7644_p2 + data_59_V_read_3_reg_8724_pp0_iter15_reg);

assign add_ln703_949_fu_7765_p2 = (sub_ln703_817_fu_7382_p2 + data_56_V_read_3_reg_8814_pp0_iter15_reg);

assign add_ln703_950_fu_7770_p2 = (add_ln703_946_reg_12805 + data_57_V_read_3_reg_8786_pp0_iter15_reg);

assign add_ln703_951_fu_7774_p2 = (add_ln703_950_fu_7770_p2 + add_ln703_949_fu_7765_p2);

assign add_ln703_952_fu_7800_p2 = (add_ln703_946_reg_12805 + sub_ln703_854_fu_7586_p2);

assign add_ln703_953_fu_7956_p2 = (sub_ln703_877_fu_7886_p2 + data_60_V_read61_reg_8691_pp0_iter16_reg);

assign add_ln703_954_fu_7338_p2 = (data_59_V_read_3_reg_8724_pp0_iter14_reg + data_60_V_read61_reg_8691_pp0_iter14_reg);

assign add_ln703_955_fu_7815_p2 = (add_ln703_954_reg_12812 + sub_ln703_862_reg_12795);

assign add_ln703_956_fu_7819_p2 = (add_ln703_920_reg_12637_pp0_iter15_reg + sub_ln703_816_reg_12740);

assign add_ln703_957_fu_7823_p2 = (add_ln703_954_reg_12812 + data_58_V_read_3_reg_8756_pp0_iter15_reg);

assign add_ln703_958_fu_7827_p2 = (add_ln703_957_fu_7823_p2 + add_ln703_956_fu_7819_p2);

assign add_ln703_959_fu_7997_p2 = (sub_ln703_889_fu_7922_p2 + data_60_V_read61_reg_8691_pp0_iter16_reg);

assign add_ln703_960_fu_8012_p2 = (sub_ln703_892_reg_12935 + data_60_V_read61_reg_8691_pp0_iter16_reg);

assign add_ln703_961_fu_8016_p2 = (sub_ln703_893_reg_12940 + data_60_V_read61_reg_8691_pp0_iter16_reg);

assign add_ln703_962_fu_8052_p2 = (sub_ln703_905_fu_7970_p2 + data_61_V_read62_reg_8663_pp0_iter16_reg);

assign add_ln703_963_fu_8062_p2 = (sub_ln703_908_fu_7983_p2 + data_61_V_read62_reg_8663_pp0_iter16_reg);

assign add_ln703_964_fu_7848_p2 = (data_60_V_read61_reg_8691_pp0_iter15_reg + data_61_V_read62_reg_8663_pp0_iter15_reg);

assign add_ln703_965_fu_8067_p2 = (add_ln703_964_reg_12985 + sub_ln703_886_fu_7910_p2);

assign add_ln703_966_fu_8100_p2 = (sub_ln703_914_fu_8020_p2 + data_61_V_read62_reg_8663_pp0_iter16_reg);

assign add_ln703_967_fu_8105_p2 = (sub_ln703_915_fu_8024_p2 + data_61_V_read62_reg_8663_pp0_iter16_reg);

assign add_ln703_968_fu_8110_p2 = (add_ln703_964_reg_12985 + sub_ln703_897_fu_7938_p2);

assign add_ln703_969_fu_8115_p2 = (sub_ln703_918_fu_8033_p2 + data_61_V_read62_reg_8663_pp0_iter16_reg);

assign add_ln703_970_fu_8125_p2 = (data_61_V_read62_reg_8663_pp0_iter16_reg + data_62_V_read_3_reg_8645_pp0_iter16_reg);

assign add_ln703_971_fu_8129_p2 = (add_ln703_970_fu_8125_p2 + sub_ln703_904_reg_12960);

assign add_ln703_972_fu_8148_p2 = (sub_ln703_882_fu_7894_p2 + data_60_V_read61_reg_8691_pp0_iter16_reg);

assign add_ln703_973_fu_8153_p2 = (add_ln703_970_fu_8125_p2 + add_ln703_972_fu_8148_p2);

assign add_ln703_974_fu_8159_p2 = (add_ln703_970_fu_8125_p2 + sub_ln703_907_fu_7978_p2);

assign add_ln703_975_fu_8170_p2 = (sub_ln703_884_fu_7902_p2 + data_60_V_read61_reg_8691_pp0_iter16_reg);

assign add_ln703_976_fu_8175_p2 = (add_ln703_970_fu_8125_p2 + add_ln703_975_fu_8170_p2);

assign add_ln703_977_fu_8186_p2 = (sub_ln703_887_fu_7914_p2 + data_60_V_read61_reg_8691_pp0_iter16_reg);

assign add_ln703_978_fu_8191_p2 = (add_ln703_970_fu_8125_p2 + add_ln703_977_fu_8186_p2);

assign add_ln703_979_fu_8197_p2 = (add_ln703_970_fu_8125_p2 + sub_ln703_910_fu_7992_p2);

assign add_ln703_980_fu_8203_p2 = (add_ln703_970_fu_8125_p2 + sub_ln703_912_fu_8002_p2);

assign add_ln703_981_fu_8214_p2 = (sub_ln703_929_fu_8095_p2 + data_62_V_read_3_reg_8645_pp0_iter16_reg);

assign add_ln703_982_fu_8239_p2 = (sub_ln703_899_fu_7942_p2 + data_60_V_read61_reg_8691_pp0_iter16_reg);

assign add_ln703_983_fu_8244_p2 = (add_ln703_970_fu_8125_p2 + add_ln703_982_fu_8239_p2);

assign add_ln703_984_fu_8250_p2 = (sub_ln703_900_fu_7946_p2 + data_61_V_read62_reg_8663_pp0_iter16_reg);

assign add_ln703_985_fu_7342_p2 = (data_62_V_read_3_reg_8645_pp0_iter14_reg + data_63_V_read_3_reg_8620_pp0_iter14_reg);

assign add_ln703_986_fu_8255_p2 = (add_ln703_985_reg_12819_pp0_iter16_reg + add_ln703_984_fu_8250_p2);

assign add_ln703_987_fu_8260_p2 = (sub_ln703_901_fu_7951_p2 + data_61_V_read62_reg_8663_pp0_iter16_reg);

assign add_ln703_994_fu_8325_p2 = (sub_ln703_909_fu_7987_p2 + data_61_V_read62_reg_8663_pp0_iter16_reg);

assign add_ln703_fu_530_p2 = (data_0_V_read_int_reg + data_1_V_read_int_reg);

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_state10_pp0_stage0_iter9 = ~(1'b1 == 1'b1);

assign ap_block_state11_pp0_stage0_iter10 = ~(1'b1 == 1'b1);

assign ap_block_state12_pp0_stage0_iter11 = ~(1'b1 == 1'b1);

assign ap_block_state13_pp0_stage0_iter12 = ~(1'b1 == 1'b1);

assign ap_block_state14_pp0_stage0_iter13 = ~(1'b1 == 1'b1);

assign ap_block_state15_pp0_stage0_iter14 = ~(1'b1 == 1'b1);

assign ap_block_state16_pp0_stage0_iter15 = ~(1'b1 == 1'b1);

assign ap_block_state17_pp0_stage0_iter16 = ~(1'b1 == 1'b1);

assign ap_block_state18_pp0_stage0_iter17 = ~(1'b1 == 1'b1);

assign ap_block_state1_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter4 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter5 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage0_iter6 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage0_iter7 = ~(1'b1 == 1'b1);

assign ap_block_state9_pp0_stage0_iter8 = ~(1'b1 == 1'b1);

assign sub_ln703_100_fu_1329_p2 = (add_ln703_199_fu_1213_p2 - data_10_V_read11_reg_10105_pp0_iter4_reg);

assign sub_ln703_101_fu_1334_p2 = (sub_ln703_83_fu_1218_p2 - data_10_V_read11_reg_10105_pp0_iter4_reg);

assign sub_ln703_102_fu_1344_p2 = (add_ln703_200_fu_1226_p2 - data_10_V_read11_reg_10105_pp0_iter4_reg);

assign sub_ln703_103_fu_1363_p2 = (sub_ln703_87_fu_1238_p2 - data_10_V_read11_reg_10105_pp0_iter4_reg);

assign sub_ln703_104_fu_1368_p2 = (add_ln703_201_fu_1243_p2 - data_10_V_read11_reg_10105_pp0_iter4_reg);

assign sub_ln703_105_fu_1373_p2 = (sub_ln703_88_fu_1248_p2 - data_10_V_read11_reg_10105_pp0_iter4_reg);

assign sub_ln703_106_fu_1378_p2 = (sub_ln703_89_fu_1252_p2 - data_10_V_read11_reg_10105_pp0_iter4_reg);

assign sub_ln703_107_fu_1383_p2 = (sub_ln703_90_fu_1257_p2 - data_10_V_read11_reg_10105_pp0_iter4_reg);

assign sub_ln703_108_fu_1388_p2 = (sub_ln703_91_fu_1261_p2 - data_10_V_read11_reg_10105_pp0_iter4_reg);

assign sub_ln703_109_fu_1407_p2 = (add_ln703_202_fu_1265_p2 - data_10_V_read11_reg_10105_pp0_iter4_reg);

assign sub_ln703_10_fu_615_p2 = (data_3_V_read_10_reg_10295_pp0_iter2_reg - add_ln703_131_reg_10354_pp0_iter2_reg);

assign sub_ln703_110_fu_1412_p2 = (add_ln703_203_fu_1270_p2 - data_10_V_read11_reg_10105_pp0_iter4_reg);

assign sub_ln703_111_fu_1417_p2 = (sub_ln703_93_fu_1275_p2 - data_10_V_read11_reg_10105_pp0_iter4_reg);

assign sub_ln703_112_fu_1422_p2 = (sub_ln703_94_fu_1280_p2 - data_10_V_read11_reg_10105_pp0_iter4_reg);

assign sub_ln703_113_fu_1427_p2 = (add_ln703_206_fu_1290_p2 - data_10_V_read11_reg_10105_pp0_iter4_reg);

assign sub_ln703_114_fu_1630_p2 = (add_ln703_207_reg_10682 - data_11_V_read12_reg_10075_pp0_iter5_reg);

assign sub_ln703_115_fu_1432_p2 = (sub_ln703_97_fu_1304_p2 - data_11_V_read12_reg_10075_pp0_iter4_reg);

assign sub_ln703_116_fu_1634_p2 = (add_ln703_208_reg_10687 - data_11_V_read12_reg_10075_pp0_iter5_reg);

assign sub_ln703_117_fu_1638_p2 = (add_ln703_210_reg_10692 - data_11_V_read12_reg_10075_pp0_iter5_reg);

assign sub_ln703_118_fu_1642_p2 = (sub_ln703_98_reg_10697 - data_11_V_read12_reg_10075_pp0_iter5_reg);

assign sub_ln703_119_fu_1442_p2 = (sub_ln703_99_fu_1324_p2 - data_11_V_read12_reg_10075_pp0_iter4_reg);

assign sub_ln703_11_fu_576_p2 = (sub_ln703_5_fu_564_p2 - data_3_V_read_10_reg_10295_pp0_iter1_reg);

assign sub_ln703_120_fu_1447_p2 = (add_ln703_211_fu_1339_p2 - data_11_V_read12_reg_10075_pp0_iter4_reg);

assign sub_ln703_121_fu_1646_p2 = (add_ln703_216_reg_10702 - data_11_V_read12_reg_10075_pp0_iter5_reg);

assign sub_ln703_122_fu_1462_p2 = (add_ln703_215_fu_1353_p2 - data_11_V_read12_reg_10075_pp0_iter4_reg);

assign sub_ln703_123_fu_1467_p2 = (sub_ln703_103_fu_1363_p2 - data_11_V_read12_reg_10075_pp0_iter4_reg);

assign sub_ln703_124_fu_1650_p2 = (sub_ln703_106_reg_10707 - data_11_V_read12_reg_10075_pp0_iter5_reg);

assign sub_ln703_125_fu_1482_p2 = (add_ln703_219_fu_1397_p2 - data_11_V_read12_reg_10075_pp0_iter4_reg);

assign sub_ln703_126_fu_1487_p2 = (add_ln703_221_fu_1402_p2 - data_11_V_read12_reg_10075_pp0_iter4_reg);

assign sub_ln703_127_fu_1662_p2 = (sub_ln703_109_reg_10722 - data_11_V_read12_reg_10075_pp0_iter5_reg);

assign sub_ln703_128_fu_1496_p2 = (sub_ln703_111_fu_1417_p2 - data_11_V_read12_reg_10075_pp0_iter4_reg);

assign sub_ln703_129_fu_1506_p2 = (sub_ln703_113_fu_1427_p2 - data_11_V_read12_reg_10075_pp0_iter4_reg);

assign sub_ln703_12_fu_627_p2 = (add_ln703_131_reg_10354_pp0_iter2_reg - data_3_V_read_10_reg_10295_pp0_iter2_reg);

assign sub_ln703_130_fu_1666_p2 = (add_ln703_222_fu_1626_p2 - data_12_V_read13_reg_10045_pp0_iter5_reg);

assign sub_ln703_131_fu_1680_p2 = (add_ln703_224_reg_10732 - data_12_V_read13_reg_10045_pp0_iter5_reg);

assign sub_ln703_132_fu_1684_p2 = (sub_ln703_118_fu_1642_p2 - data_12_V_read13_reg_10045_pp0_iter5_reg);

assign sub_ln703_133_fu_1532_p2 = (add_ln703_225_fu_1452_p2 - data_12_V_read13_reg_10045_pp0_iter4_reg);

assign sub_ln703_134_fu_1689_p2 = (add_ln703_226_reg_10737 - data_12_V_read13_reg_10045_pp0_iter5_reg);

assign sub_ln703_135_fu_1698_p2 = (sub_ln703_123_reg_10747 - data_12_V_read13_reg_10045_pp0_iter5_reg);

assign sub_ln703_136_fu_1702_p2 = (add_ln703_227_reg_10752 - data_12_V_read13_reg_10045_pp0_iter5_reg);

assign sub_ln703_137_fu_1548_p2 = (add_ln703_228_fu_1477_p2 - data_12_V_read13_reg_10045_pp0_iter4_reg);

assign sub_ln703_138_fu_1706_p2 = (sub_ln703_124_fu_1650_p2 - data_12_V_read13_reg_10045_pp0_iter5_reg);

assign sub_ln703_139_fu_1711_p2 = (add_ln703_229_fu_1654_p2 - data_12_V_read13_reg_10045_pp0_iter5_reg);

assign sub_ln703_13_fu_689_p2 = (sub_ln703_6_reg_10408 - data_4_V_read_10_reg_10273_pp0_iter3_reg);

assign sub_ln703_140_fu_1716_p2 = (add_ln703_230_fu_1658_p2 - data_12_V_read13_reg_10045_pp0_iter5_reg);

assign sub_ln703_141_fu_1553_p2 = (sub_ln703_126_fu_1487_p2 - data_12_V_read13_reg_10045_pp0_iter4_reg);

assign sub_ln703_142_fu_1558_p2 = (add_ln703_232_fu_1492_p2 - data_12_V_read13_reg_10045_pp0_iter4_reg);

assign sub_ln703_143_fu_1725_p2 = (sub_ln703_127_fu_1662_p2 - data_12_V_read13_reg_10045_pp0_iter5_reg);

assign sub_ln703_144_fu_1730_p2 = (sub_ln703_128_reg_10762 - data_12_V_read13_reg_10045_pp0_iter5_reg);

assign sub_ln703_145_fu_1734_p2 = (add_ln703_233_reg_10767 - data_12_V_read13_reg_10045_pp0_iter5_reg);

assign sub_ln703_146_fu_1580_p2 = (sub_ln703_129_fu_1506_p2 - data_12_V_read13_reg_10045_pp0_iter4_reg);

assign sub_ln703_147_fu_1738_p2 = (sub_ln703_130_fu_1666_p2 - data_13_V_read14_reg_10015_pp0_iter5_reg);

assign sub_ln703_148_fu_1743_p2 = (add_ln703_234_fu_1671_p2 - data_13_V_read14_reg_10015_pp0_iter5_reg);

assign sub_ln703_149_fu_1748_p2 = (add_ln703_235_fu_1676_p2 - data_13_V_read14_reg_10015_pp0_iter5_reg);

assign sub_ln703_14_fu_693_p2 = (add_ln703_132_reg_10414 - data_4_V_read_10_reg_10273_pp0_iter3_reg);

assign sub_ln703_150_fu_1763_p2 = (add_ln703_236_reg_10772 - data_13_V_read14_reg_10015_pp0_iter5_reg);

assign sub_ln703_151_fu_1767_p2 = (add_ln703_238_reg_10777 - data_13_V_read14_reg_10015_pp0_iter5_reg);

assign sub_ln703_152_fu_1599_p2 = (add_ln703_240_fu_1526_p2 - data_13_V_read14_reg_10015_pp0_iter4_reg);

assign sub_ln703_153_fu_1775_p2 = (add_ln703_241_fu_1693_p2 - data_13_V_read14_reg_10015_pp0_iter5_reg);

assign sub_ln703_154_fu_1609_p2 = (add_ln703_244_fu_1542_p2 - data_13_V_read14_reg_10015_pp0_iter4_reg);

assign sub_ln703_155_fu_1780_p2 = (sub_ln703_135_fu_1698_p2 - data_13_V_read14_reg_10015_pp0_iter5_reg);

assign sub_ln703_156_fu_1785_p2 = (sub_ln703_136_fu_1702_p2 - data_13_V_read14_reg_10015_pp0_iter5_reg);

assign sub_ln703_157_fu_1790_p2 = (sub_ln703_137_reg_10787 - data_13_V_read14_reg_10015_pp0_iter5_reg);

assign sub_ln703_158_fu_1794_p2 = (sub_ln703_139_fu_1711_p2 - data_13_V_read14_reg_10015_pp0_iter5_reg);

assign sub_ln703_159_fu_1799_p2 = (sub_ln703_140_fu_1716_p2 - data_13_V_read14_reg_10015_pp0_iter5_reg);

assign sub_ln703_15_fu_631_p2 = (add_ln703_133_fu_603_p2 - data_4_V_read_10_reg_10273_pp0_iter2_reg);

assign sub_ln703_160_fu_1804_p2 = (add_ln703_245_fu_1721_p2 - data_13_V_read14_reg_10015_pp0_iter5_reg);

assign sub_ln703_161_fu_1809_p2 = (sub_ln703_141_reg_10792 - data_13_V_read14_reg_10015_pp0_iter5_reg);

assign sub_ln703_162_fu_1813_p2 = (sub_ln703_142_reg_10797 - data_13_V_read14_reg_10015_pp0_iter5_reg);

assign sub_ln703_163_fu_1817_p2 = (add_ln703_247_reg_10802 - data_13_V_read14_reg_10015_pp0_iter5_reg);

assign sub_ln703_164_fu_1826_p2 = (add_ln703_250_reg_10807 - data_13_V_read14_reg_10015_pp0_iter5_reg);

assign sub_ln703_165_fu_1830_p2 = (sub_ln703_146_reg_10812 - data_13_V_read14_reg_10015_pp0_iter5_reg);

assign sub_ln703_166_fu_1834_p2 = (sub_ln703_148_fu_1743_p2 - data_14_V_read15_reg_9987_pp0_iter5_reg);

assign sub_ln703_167_fu_1839_p2 = (sub_ln703_149_fu_1748_p2 - data_14_V_read15_reg_9987_pp0_iter5_reg);

assign sub_ln703_168_fu_1844_p2 = (add_ln703_251_fu_1753_p2 - data_14_V_read15_reg_9987_pp0_iter5_reg);

assign sub_ln703_169_fu_1849_p2 = (add_ln703_253_fu_1758_p2 - data_14_V_read15_reg_9987_pp0_iter5_reg);

assign sub_ln703_16_fu_640_p2 = (data_4_V_read_10_reg_10273_pp0_iter2_reg - add_ln703_134_reg_10385);

assign sub_ln703_170_fu_1859_p2 = (sub_ln703_150_fu_1763_p2 - data_14_V_read15_reg_9987_pp0_iter5_reg);

assign sub_ln703_171_fu_1864_p2 = (add_ln703_260_reg_10817 - data_14_V_read15_reg_9987_pp0_iter5_reg);

assign sub_ln703_172_fu_1868_p2 = (sub_ln703_151_fu_1767_p2 - data_14_V_read15_reg_9987_pp0_iter5_reg);

assign sub_ln703_173_fu_1873_p2 = (sub_ln703_152_reg_10822 - data_14_V_read15_reg_9987_pp0_iter5_reg);

assign sub_ln703_174_fu_1877_p2 = (add_ln703_262_reg_10827 - data_14_V_read15_reg_9987_pp0_iter5_reg);

assign sub_ln703_175_fu_1881_p2 = (add_ln703_263_fu_1771_p2 - data_14_V_read15_reg_9987_pp0_iter5_reg);

assign sub_ln703_176_fu_1900_p2 = (sub_ln703_154_reg_10832 - data_14_V_read15_reg_9987_pp0_iter5_reg);

assign sub_ln703_177_fu_1904_p2 = (sub_ln703_156_fu_1785_p2 - data_14_V_read15_reg_9987_pp0_iter5_reg);

assign sub_ln703_178_fu_1909_p2 = (sub_ln703_157_fu_1790_p2 - data_14_V_read15_reg_9987_pp0_iter5_reg);

assign sub_ln703_179_fu_1919_p2 = (sub_ln703_160_fu_1804_p2 - data_14_V_read15_reg_9987_pp0_iter5_reg);

assign sub_ln703_17_fu_653_p2 = (sub_ln703_9_fu_611_p2 - data_4_V_read_10_reg_10273_pp0_iter2_reg);

assign sub_ln703_180_fu_1929_p2 = (sub_ln703_162_fu_1813_p2 - data_14_V_read15_reg_9987_pp0_iter5_reg);

assign sub_ln703_181_fu_1944_p2 = (add_ln703_264_fu_1821_p2 - data_14_V_read15_reg_9987_pp0_iter5_reg);

assign sub_ln703_182_fu_1949_p2 = (sub_ln703_164_fu_1826_p2 - data_14_V_read15_reg_9987_pp0_iter5_reg);

assign sub_ln703_183_fu_1959_p2 = (sub_ln703_168_fu_1844_p2 - data_15_V_read16_reg_9962_pp0_iter5_reg);

assign sub_ln703_184_fu_1984_p2 = (add_ln703_266_fu_1854_p2 - data_15_V_read16_reg_9962_pp0_iter5_reg);

assign sub_ln703_185_fu_1989_p2 = (sub_ln703_172_fu_1868_p2 - data_15_V_read16_reg_9962_pp0_iter5_reg);

assign sub_ln703_186_fu_1994_p2 = (sub_ln703_173_fu_1873_p2 - data_15_V_read16_reg_9962_pp0_iter5_reg);

assign sub_ln703_187_fu_1999_p2 = (sub_ln703_174_fu_1877_p2 - data_15_V_read16_reg_9962_pp0_iter5_reg);

assign sub_ln703_188_fu_2004_p2 = (add_ln703_268_fu_1886_p2 - data_15_V_read16_reg_9962_pp0_iter5_reg);

assign sub_ln703_189_fu_2014_p2 = (add_ln703_271_fu_1895_p2 - data_15_V_read16_reg_9962_pp0_iter5_reg);

assign sub_ln703_18_fu_658_p2 = (sub_ln703_8_reg_10392 - data_4_V_read_10_reg_10273_pp0_iter2_reg);

assign sub_ln703_190_fu_2024_p2 = (sub_ln703_178_fu_1909_p2 - data_15_V_read16_reg_9962_pp0_iter5_reg);

assign sub_ln703_191_fu_2029_p2 = (add_ln703_273_fu_1914_p2 - data_15_V_read16_reg_9962_pp0_iter5_reg);

assign sub_ln703_192_fu_2044_p2 = (add_ln703_274_fu_1924_p2 - data_15_V_read16_reg_9962_pp0_iter5_reg);

assign sub_ln703_193_fu_2049_p2 = (sub_ln703_180_fu_1929_p2 - data_15_V_read16_reg_9962_pp0_iter5_reg);

assign sub_ln703_194_fu_2054_p2 = (add_ln703_276_fu_1934_p2 - data_15_V_read16_reg_9962_pp0_iter5_reg);

assign sub_ln703_195_fu_2059_p2 = (add_ln703_277_fu_1939_p2 - data_15_V_read16_reg_9962_pp0_iter5_reg);

assign sub_ln703_196_fu_2074_p2 = (sub_ln703_181_fu_1944_p2 - data_15_V_read16_reg_9962_pp0_iter5_reg);

assign sub_ln703_197_fu_2079_p2 = (add_ln703_278_fu_1954_p2 - data_15_V_read16_reg_9962_pp0_iter5_reg);

assign sub_ln703_198_fu_2099_p2 = (add_ln703_282_fu_1973_p2 - data_16_V_read17_reg_9935_pp0_iter5_reg);

assign sub_ln703_199_fu_2246_p2 = (add_ln703_283_reg_10873 - data_16_V_read17_reg_9935_pp0_iter6_reg);

assign sub_ln703_19_fu_705_p2 = (sub_ln703_10_reg_10420 - data_4_V_read_10_reg_10273_pp0_iter3_reg);

assign sub_ln703_1_fu_540_p2 = (data_0_V_read_10_reg_10329 - data_1_V_read_10_reg_10323);

assign sub_ln703_200_fu_2115_p2 = (sub_ln703_188_fu_2004_p2 - data_16_V_read17_reg_9935_pp0_iter5_reg);

assign sub_ln703_201_fu_2258_p2 = (add_ln703_285_reg_10888 - data_16_V_read17_reg_9935_pp0_iter6_reg);

assign sub_ln703_202_fu_2120_p2 = (sub_ln703_189_fu_2014_p2 - data_16_V_read17_reg_9935_pp0_iter5_reg);

assign sub_ln703_203_fu_2131_p2 = (add_ln703_287_fu_2019_p2 - data_16_V_read17_reg_9935_pp0_iter5_reg);

assign sub_ln703_204_fu_2142_p2 = (sub_ln703_190_fu_2024_p2 - data_16_V_read17_reg_9935_pp0_iter5_reg);

assign sub_ln703_205_fu_2262_p2 = (sub_ln703_191_reg_10893 - data_16_V_read17_reg_9935_pp0_iter6_reg);

assign sub_ln703_206_fu_2266_p2 = (add_ln703_289_reg_10898 - data_16_V_read17_reg_9935_pp0_iter6_reg);

assign sub_ln703_207_fu_2274_p2 = (add_ln703_290_reg_10903 - data_16_V_read17_reg_9935_pp0_iter6_reg);

assign sub_ln703_208_fu_2152_p2 = (sub_ln703_192_fu_2044_p2 - data_16_V_read17_reg_9935_pp0_iter5_reg);

assign sub_ln703_209_fu_2157_p2 = (sub_ln703_195_fu_2059_p2 - data_16_V_read17_reg_9935_pp0_iter5_reg);

assign sub_ln703_20_fu_662_p2 = (add_ln703_134_reg_10385 - data_4_V_read_10_reg_10273_pp0_iter2_reg);

assign sub_ln703_210_fu_2162_p2 = (add_ln703_293_fu_2069_p2 - data_16_V_read17_reg_9935_pp0_iter5_reg);

assign sub_ln703_211_fu_2278_p2 = (sub_ln703_196_reg_10913 - data_16_V_read17_reg_9935_pp0_iter6_reg);

assign sub_ln703_212_fu_2173_p2 = (sub_ln703_197_fu_2079_p2 - data_16_V_read17_reg_9935_pp0_iter5_reg);

assign sub_ln703_213_fu_2282_p2 = (add_ln703_296_fu_2238_p2 - data_17_V_read18_reg_9904_pp0_iter6_reg);

assign sub_ln703_214_fu_2287_p2 = (add_ln703_298_fu_2242_p2 - data_17_V_read18_reg_9904_pp0_iter6_reg);

assign sub_ln703_215_fu_2292_p2 = (add_ln703_300_reg_10930 - data_17_V_read18_reg_9904_pp0_iter6_reg);

assign sub_ln703_216_fu_2296_p2 = (sub_ln703_198_reg_10935 - data_17_V_read18_reg_9904_pp0_iter6_reg);

assign sub_ln703_217_fu_2305_p2 = (add_ln703_301_fu_2250_p2 - data_17_V_read18_reg_9904_pp0_iter6_reg);

assign sub_ln703_218_fu_2310_p2 = (add_ln703_303_reg_10940 - data_17_V_read18_reg_9904_pp0_iter6_reg);

assign sub_ln703_219_fu_2314_p2 = (add_ln703_304_reg_10945 - data_17_V_read18_reg_9904_pp0_iter6_reg);

assign sub_ln703_21_fu_709_p2 = (sub_ln703_11_reg_10398_pp0_iter3_reg - data_4_V_read_10_reg_10273_pp0_iter3_reg);

assign sub_ln703_220_fu_2318_p2 = (add_ln703_305_fu_2254_p2 - data_17_V_read18_reg_9904_pp0_iter6_reg);

assign sub_ln703_221_fu_2332_p2 = (add_ln703_307_reg_10960 - data_17_V_read18_reg_9904_pp0_iter6_reg);

assign sub_ln703_222_fu_2340_p2 = (add_ln703_309_reg_10970 - data_17_V_read18_reg_9904_pp0_iter6_reg);

assign sub_ln703_223_fu_2344_p2 = (sub_ln703_204_reg_10975 - data_17_V_read18_reg_9904_pp0_iter6_reg);

assign sub_ln703_224_fu_2348_p2 = (sub_ln703_205_fu_2262_p2 - data_17_V_read18_reg_9904_pp0_iter6_reg);

assign sub_ln703_225_fu_2358_p2 = (add_ln703_312_fu_2270_p2 - data_17_V_read18_reg_9904_pp0_iter6_reg);

assign sub_ln703_226_fu_2363_p2 = (sub_ln703_207_fu_2274_p2 - data_17_V_read18_reg_9904_pp0_iter6_reg);

assign sub_ln703_227_fu_2368_p2 = (sub_ln703_209_reg_10990 - data_17_V_read18_reg_9904_pp0_iter6_reg);

assign sub_ln703_228_fu_2372_p2 = (sub_ln703_210_reg_10995 - data_17_V_read18_reg_9904_pp0_iter6_reg);

assign sub_ln703_229_fu_2376_p2 = (sub_ln703_211_fu_2278_p2 - data_17_V_read18_reg_9904_pp0_iter6_reg);

assign sub_ln703_22_fu_713_p2 = (add_ln703_135_reg_10425 - data_4_V_read_10_reg_10273_pp0_iter3_reg);

assign sub_ln703_230_fu_2194_p2 = (add_ln703_314_fu_2167_p2 - data_17_V_read18_reg_9904_pp0_iter5_reg);

assign sub_ln703_231_fu_2381_p2 = (sub_ln703_212_reg_11000 - data_17_V_read18_reg_9904_pp0_iter6_reg);

assign sub_ln703_232_fu_2385_p2 = (sub_ln703_213_fu_2282_p2 - data_18_V_read_8_reg_9874_pp0_iter6_reg);

assign sub_ln703_233_fu_2390_p2 = (sub_ln703_215_fu_2292_p2 - data_18_V_read_8_reg_9874_pp0_iter6_reg);

assign sub_ln703_234_fu_2395_p2 = (sub_ln703_216_fu_2296_p2 - data_18_V_read_8_reg_9874_pp0_iter6_reg);

assign sub_ln703_235_fu_2400_p2 = (add_ln703_315_fu_2300_p2 - data_18_V_read_8_reg_9874_pp0_iter6_reg);

assign sub_ln703_236_fu_2415_p2 = (sub_ln703_220_fu_2318_p2 - data_18_V_read_8_reg_9874_pp0_iter6_reg);

assign sub_ln703_237_fu_2214_p2 = (add_ln703_317_fu_2182_p2 - data_18_V_read_8_reg_9874_pp0_iter5_reg);

assign sub_ln703_238_fu_2424_p2 = (add_ln703_318_fu_2323_p2 - data_18_V_read_8_reg_9874_pp0_iter6_reg);

assign sub_ln703_239_fu_2429_p2 = (add_ln703_319_fu_2328_p2 - data_18_V_read_8_reg_9874_pp0_iter6_reg);

assign sub_ln703_23_fu_666_p2 = (add_ln703_136_fu_623_p2 - data_4_V_read_10_reg_10273_pp0_iter2_reg);

assign sub_ln703_240_fu_2434_p2 = (sub_ln703_221_fu_2332_p2 - data_18_V_read_8_reg_9874_pp0_iter6_reg);

assign sub_ln703_241_fu_2439_p2 = (add_ln703_320_fu_2336_p2 - data_18_V_read_8_reg_9874_pp0_iter6_reg);

assign sub_ln703_242_fu_2444_p2 = (sub_ln703_222_fu_2340_p2 - data_18_V_read_8_reg_9874_pp0_iter6_reg);

assign sub_ln703_243_fu_2454_p2 = (add_ln703_321_fu_2353_p2 - data_18_V_read_8_reg_9874_pp0_iter6_reg);

assign sub_ln703_244_fu_2468_p2 = (add_ln703_323_reg_11005 - data_18_V_read_8_reg_9874_pp0_iter6_reg);

assign sub_ln703_245_fu_2472_p2 = (sub_ln703_227_fu_2368_p2 - data_18_V_read_8_reg_9874_pp0_iter6_reg);

assign sub_ln703_246_fu_2477_p2 = (sub_ln703_228_fu_2372_p2 - data_18_V_read_8_reg_9874_pp0_iter6_reg);

assign sub_ln703_247_fu_2482_p2 = (sub_ln703_229_fu_2376_p2 - data_18_V_read_8_reg_9874_pp0_iter6_reg);

assign sub_ln703_248_fu_2487_p2 = (sub_ln703_230_reg_11010 - data_18_V_read_8_reg_9874_pp0_iter6_reg);

assign sub_ln703_249_fu_2496_p2 = (sub_ln703_232_fu_2385_p2 - data_19_V_read_8_reg_9845_pp0_iter6_reg);

assign sub_ln703_24_fu_717_p2 = (sub_ln703_13_fu_689_p2 - data_5_V_read_9_reg_10245_pp0_iter3_reg);

assign sub_ln703_250_fu_2501_p2 = (sub_ln703_235_fu_2400_p2 - data_19_V_read_8_reg_9845_pp0_iter6_reg);

assign sub_ln703_251_fu_2506_p2 = (add_ln703_324_fu_2405_p2 - data_19_V_read_8_reg_9845_pp0_iter6_reg);

assign sub_ln703_252_fu_2511_p2 = (add_ln703_328_reg_11015 - data_19_V_read_8_reg_9845_pp0_iter6_reg);

assign sub_ln703_253_fu_2515_p2 = (add_ln703_329_fu_2410_p2 - data_19_V_read_8_reg_9845_pp0_iter6_reg);

assign sub_ln703_254_fu_2525_p2 = (sub_ln703_236_fu_2415_p2 - data_19_V_read_8_reg_9845_pp0_iter6_reg);

assign sub_ln703_255_fu_2530_p2 = (add_ln703_333_reg_11025 - data_19_V_read_8_reg_9845_pp0_iter6_reg);

assign sub_ln703_256_fu_2534_p2 = (add_ln703_335_fu_2420_p2 - data_19_V_read_8_reg_9845_pp0_iter6_reg);

assign sub_ln703_257_fu_2539_p2 = (sub_ln703_238_fu_2424_p2 - data_19_V_read_8_reg_9845_pp0_iter6_reg);

assign sub_ln703_258_fu_2544_p2 = (sub_ln703_239_fu_2429_p2 - data_19_V_read_8_reg_9845_pp0_iter6_reg);

assign sub_ln703_259_fu_2549_p2 = (sub_ln703_240_fu_2434_p2 - data_19_V_read_8_reg_9845_pp0_iter6_reg);

assign sub_ln703_25_fu_722_p2 = (sub_ln703_14_fu_693_p2 - data_5_V_read_9_reg_10245_pp0_iter3_reg);

assign sub_ln703_260_fu_2559_p2 = (sub_ln703_242_fu_2444_p2 - data_19_V_read_8_reg_9845_pp0_iter6_reg);

assign sub_ln703_261_fu_2569_p2 = (add_ln703_336_fu_2449_p2 - data_19_V_read_8_reg_9845_pp0_iter6_reg);

assign sub_ln703_262_fu_2574_p2 = (sub_ln703_243_fu_2454_p2 - data_19_V_read_8_reg_9845_pp0_iter6_reg);

assign sub_ln703_263_fu_2579_p2 = (add_ln703_337_fu_2459_p2 - data_19_V_read_8_reg_9845_pp0_iter6_reg);

assign sub_ln703_264_fu_2584_p2 = (add_ln703_339_fu_2464_p2 - data_19_V_read_8_reg_9845_pp0_iter6_reg);

assign sub_ln703_265_fu_2613_p2 = (sub_ln703_247_fu_2482_p2 - data_19_V_read_8_reg_9845_pp0_iter6_reg);

assign sub_ln703_266_fu_2618_p2 = (sub_ln703_248_fu_2487_p2 - data_19_V_read_8_reg_9845_pp0_iter6_reg);

assign sub_ln703_267_fu_2623_p2 = (add_ln703_340_fu_2491_p2 - data_19_V_read_8_reg_9845_pp0_iter6_reg);

assign sub_ln703_268_fu_2783_p2 = (sub_ln703_249_reg_11056 - data_20_V_read21_reg_9814_pp0_iter7_reg);

assign sub_ln703_269_fu_2787_p2 = (sub_ln703_251_reg_11066 - data_20_V_read21_reg_9814_pp0_iter7_reg);

assign sub_ln703_26_fu_727_p2 = (add_ln703_137_fu_697_p2 - data_5_V_read_9_reg_10245_pp0_iter3_reg);

assign sub_ln703_270_fu_2628_p2 = (sub_ln703_252_fu_2511_p2 - data_20_V_read21_reg_9814_pp0_iter6_reg);

assign sub_ln703_271_fu_2791_p2 = (add_ln703_342_reg_11071 - data_20_V_read21_reg_9814_pp0_iter7_reg);

assign sub_ln703_272_fu_2647_p2 = (sub_ln703_255_fu_2530_p2 - data_20_V_read21_reg_9814_pp0_iter6_reg);

assign sub_ln703_273_fu_2799_p2 = (sub_ln703_256_reg_11081 - data_20_V_read21_reg_9814_pp0_iter7_reg);

assign sub_ln703_274_fu_2652_p2 = (sub_ln703_258_fu_2544_p2 - data_20_V_read21_reg_9814_pp0_iter6_reg);

assign sub_ln703_275_fu_2662_p2 = (add_ln703_343_fu_2554_p2 - data_20_V_read21_reg_9814_pp0_iter6_reg);

assign sub_ln703_276_fu_2667_p2 = (add_ln703_345_fu_2564_p2 - data_20_V_read21_reg_9814_pp0_iter6_reg);

assign sub_ln703_277_fu_2803_p2 = (sub_ln703_261_reg_11091 - data_20_V_read21_reg_9814_pp0_iter7_reg);

assign sub_ln703_278_fu_2807_p2 = (sub_ln703_262_reg_11096 - data_20_V_read21_reg_9814_pp0_iter7_reg);

assign sub_ln703_279_fu_2815_p2 = (add_ln703_346_reg_11106 - data_20_V_read21_reg_9814_pp0_iter7_reg);

assign sub_ln703_27_fu_732_p2 = (sub_ln703_15_reg_10430 - data_5_V_read_9_reg_10245_pp0_iter3_reg);

assign sub_ln703_280_fu_2819_p2 = (add_ln703_350_reg_11111 - data_20_V_read21_reg_9814_pp0_iter7_reg);

assign sub_ln703_281_fu_2688_p2 = (add_ln703_351_fu_2608_p2 - data_20_V_read21_reg_9814_pp0_iter6_reg);

assign sub_ln703_282_fu_2827_p2 = (sub_ln703_265_reg_11116 - data_20_V_read21_reg_9814_pp0_iter7_reg);

assign sub_ln703_283_fu_2693_p2 = (sub_ln703_266_fu_2618_p2 - data_20_V_read21_reg_9814_pp0_iter6_reg);

assign sub_ln703_284_fu_2698_p2 = (sub_ln703_267_fu_2623_p2 - data_20_V_read21_reg_9814_pp0_iter6_reg);

assign sub_ln703_285_fu_2836_p2 = (sub_ln703_269_fu_2787_p2 - data_21_V_read22_reg_9784_pp0_iter7_reg);

assign sub_ln703_286_fu_2845_p2 = (add_ln703_352_reg_11126 - data_21_V_read22_reg_9784_pp0_iter7_reg);

assign sub_ln703_287_fu_2849_p2 = (sub_ln703_271_fu_2791_p2 - data_21_V_read22_reg_9784_pp0_iter7_reg);

assign sub_ln703_288_fu_2854_p2 = (add_ln703_353_fu_2795_p2 - data_21_V_read22_reg_9784_pp0_iter7_reg);

assign sub_ln703_289_fu_2703_p2 = (add_ln703_355_fu_2642_p2 - data_21_V_read22_reg_9784_pp0_iter6_reg);

assign sub_ln703_28_fu_671_p2 = (data_5_V_read_9_reg_10245_pp0_iter2_reg - add_ln703_139_fu_636_p2);

assign sub_ln703_290_fu_2859_p2 = (sub_ln703_272_reg_11138 - data_21_V_read22_reg_9784_pp0_iter7_reg);

assign sub_ln703_291_fu_2863_p2 = (sub_ln703_274_reg_11143 - data_21_V_read22_reg_9784_pp0_iter7_reg);

assign sub_ln703_292_fu_2867_p2 = (add_ln703_356_reg_11148 - data_21_V_read22_reg_9784_pp0_iter7_reg);

assign sub_ln703_293_fu_2708_p2 = (sub_ln703_276_fu_2667_p2 - data_21_V_read22_reg_9784_pp0_iter6_reg);

assign sub_ln703_294_fu_2875_p2 = (add_ln703_357_fu_2811_p2 - data_21_V_read22_reg_9784_pp0_iter7_reg);

assign sub_ln703_295_fu_2880_p2 = (add_ln703_360_reg_11158 - data_21_V_read22_reg_9784_pp0_iter7_reg);

assign sub_ln703_296_fu_2713_p2 = (add_ln703_361_fu_2683_p2 - data_21_V_read22_reg_9784_pp0_iter6_reg);

assign sub_ln703_297_fu_2884_p2 = (sub_ln703_279_fu_2815_p2 - data_21_V_read22_reg_9784_pp0_iter7_reg);

assign sub_ln703_298_fu_2889_p2 = (sub_ln703_280_fu_2819_p2 - data_21_V_read22_reg_9784_pp0_iter7_reg);

assign sub_ln703_299_fu_2894_p2 = (sub_ln703_281_reg_11163 - data_21_V_read22_reg_9784_pp0_iter7_reg);

assign sub_ln703_29_fu_749_p2 = (sub_ln703_16_reg_10436 - data_5_V_read_9_reg_10245_pp0_iter3_reg);

assign sub_ln703_2_fu_552_p2 = (sub_ln703_reg_10342 - data_2_V_read_10_reg_10312_pp0_iter1_reg);

assign sub_ln703_300_fu_2898_p2 = (add_ln703_363_fu_2823_p2 - data_21_V_read22_reg_9784_pp0_iter7_reg);

assign sub_ln703_301_fu_2718_p2 = (sub_ln703_283_fu_2693_p2 - data_21_V_read22_reg_9784_pp0_iter6_reg);

assign sub_ln703_302_fu_2907_p2 = (add_ln703_364_fu_2831_p2 - data_22_V_read23_reg_9756_pp0_iter7_reg);

assign sub_ln703_303_fu_2912_p2 = (sub_ln703_285_fu_2836_p2 - data_22_V_read23_reg_9756_pp0_iter7_reg);

assign sub_ln703_304_fu_2917_p2 = (add_ln703_365_fu_2841_p2 - data_22_V_read23_reg_9756_pp0_iter7_reg);

assign sub_ln703_305_fu_2922_p2 = (sub_ln703_286_fu_2845_p2 - data_22_V_read23_reg_9756_pp0_iter7_reg);

assign sub_ln703_306_fu_2931_p2 = (sub_ln703_290_fu_2859_p2 - data_22_V_read23_reg_9756_pp0_iter7_reg);

assign sub_ln703_307_fu_2941_p2 = (sub_ln703_291_fu_2863_p2 - data_22_V_read23_reg_9756_pp0_iter7_reg);

assign sub_ln703_308_fu_2946_p2 = (sub_ln703_292_fu_2867_p2 - data_22_V_read23_reg_9756_pp0_iter7_reg);

assign sub_ln703_309_fu_2951_p2 = (add_ln703_366_fu_2871_p2 - data_22_V_read23_reg_9756_pp0_iter7_reg);

assign sub_ln703_30_fu_753_p2 = (add_ln703_140_reg_10442 - data_5_V_read_9_reg_10245_pp0_iter3_reg);

assign sub_ln703_310_fu_2978_p2 = (sub_ln703_298_fu_2889_p2 - data_22_V_read23_reg_9756_pp0_iter7_reg);

assign sub_ln703_311_fu_2988_p2 = (sub_ln703_300_fu_2898_p2 - data_22_V_read23_reg_9756_pp0_iter7_reg);

assign sub_ln703_312_fu_2993_p2 = (add_ln703_367_fu_2903_p2 - data_22_V_read23_reg_9756_pp0_iter7_reg);

assign sub_ln703_313_fu_2998_p2 = (sub_ln703_302_fu_2907_p2 - data_23_V_read24_reg_9730_pp0_iter7_reg);

assign sub_ln703_314_fu_3003_p2 = (add_ln703_371_reg_11193 - data_23_V_read24_reg_9730_pp0_iter7_reg);

assign sub_ln703_315_fu_3021_p2 = (sub_ln703_303_fu_2912_p2 - data_23_V_read24_reg_9730_pp0_iter7_reg);

assign sub_ln703_316_fu_3026_p2 = (sub_ln703_304_fu_2917_p2 - data_23_V_read24_reg_9730_pp0_iter7_reg);

assign sub_ln703_317_fu_3031_p2 = (add_ln703_372_fu_2927_p2 - data_23_V_read24_reg_9730_pp0_iter7_reg);

assign sub_ln703_318_fu_3036_p2 = (sub_ln703_306_fu_2931_p2 - data_23_V_read24_reg_9730_pp0_iter7_reg);

assign sub_ln703_319_fu_3041_p2 = (add_ln703_374_fu_2936_p2 - data_23_V_read24_reg_9730_pp0_iter7_reg);

assign sub_ln703_31_fu_761_p2 = (add_ln703_144_reg_10403_pp0_iter3_reg - data_5_V_read_9_reg_10245_pp0_iter3_reg);

assign sub_ln703_320_fu_3056_p2 = (sub_ln703_307_fu_2941_p2 - data_23_V_read24_reg_9730_pp0_iter7_reg);

assign sub_ln703_321_fu_3066_p2 = (sub_ln703_309_fu_2951_p2 - data_23_V_read24_reg_9730_pp0_iter7_reg);

assign sub_ln703_322_fu_3071_p2 = (add_ln703_377_fu_2956_p2 - data_23_V_read24_reg_9730_pp0_iter7_reg);

assign sub_ln703_323_fu_3076_p2 = (add_ln703_378_fu_2960_p2 - data_23_V_read24_reg_9730_pp0_iter7_reg);

assign sub_ln703_324_fu_3091_p2 = (add_ln703_379_fu_2964_p2 - data_23_V_read24_reg_9730_pp0_iter7_reg);

assign sub_ln703_325_fu_3096_p2 = (add_ln703_380_fu_2969_p2 - data_23_V_read24_reg_9730_pp0_iter7_reg);

assign sub_ln703_326_fu_3101_p2 = (add_ln703_381_fu_2973_p2 - data_23_V_read24_reg_9730_pp0_iter7_reg);

assign sub_ln703_327_fu_3106_p2 = (add_ln703_382_fu_2983_p2 - data_23_V_read24_reg_9730_pp0_iter7_reg);

assign sub_ln703_328_fu_3111_p2 = (sub_ln703_311_fu_2988_p2 - data_23_V_read24_reg_9730_pp0_iter7_reg);

assign sub_ln703_329_fu_3126_p2 = (sub_ln703_312_fu_2993_p2 - data_23_V_read24_reg_9730_pp0_iter7_reg);

assign sub_ln703_32_fu_765_p2 = (add_ln703_141_reg_10447 - data_5_V_read_9_reg_10245_pp0_iter3_reg);

assign sub_ln703_330_fu_3372_p2 = (sub_ln703_313_reg_11257 - data_24_V_read25_reg_9704_pp0_iter8_reg);

assign sub_ln703_331_fu_3140_p2 = (sub_ln703_314_fu_3003_p2 - data_24_V_read25_reg_9704_pp0_iter7_reg);

assign sub_ln703_332_fu_3376_p2 = (add_ln703_386_reg_11262 - data_24_V_read25_reg_9704_pp0_iter8_reg);

assign sub_ln703_333_fu_3155_p2 = (sub_ln703_316_fu_3026_p2 - data_24_V_read25_reg_9704_pp0_iter7_reg);

assign sub_ln703_334_fu_3175_p2 = (sub_ln703_318_fu_3036_p2 - data_24_V_read25_reg_9704_pp0_iter7_reg);

assign sub_ln703_335_fu_3384_p2 = (add_ln703_390_reg_11272 - data_24_V_read25_reg_9704_pp0_iter8_reg);

assign sub_ln703_336_fu_3180_p2 = (add_ln703_391_fu_3061_p2 - data_24_V_read25_reg_9704_pp0_iter7_reg);

assign sub_ln703_337_fu_3190_p2 = (sub_ln703_322_fu_3071_p2 - data_24_V_read25_reg_9704_pp0_iter7_reg);

assign sub_ln703_338_fu_3195_p2 = (sub_ln703_323_fu_3076_p2 - data_24_V_read25_reg_9704_pp0_iter7_reg);

assign sub_ln703_339_fu_3200_p2 = (add_ln703_394_fu_3086_p2 - data_24_V_read25_reg_9704_pp0_iter7_reg);

assign sub_ln703_33_fu_769_p2 = (sub_ln703_18_reg_10459 - data_5_V_read_9_reg_10245_pp0_iter3_reg);

assign sub_ln703_340_fu_3205_p2 = (sub_ln703_324_fu_3091_p2 - data_24_V_read25_reg_9704_pp0_iter7_reg);

assign sub_ln703_341_fu_3388_p2 = (sub_ln703_326_reg_11277 - data_24_V_read25_reg_9704_pp0_iter8_reg);

assign sub_ln703_342_fu_3215_p2 = (sub_ln703_327_fu_3106_p2 - data_24_V_read25_reg_9704_pp0_iter7_reg);

assign sub_ln703_343_fu_3392_p2 = (sub_ln703_328_reg_11282 - data_24_V_read25_reg_9704_pp0_iter8_reg);

assign sub_ln703_344_fu_3220_p2 = (add_ln703_397_fu_3121_p2 - data_24_V_read25_reg_9704_pp0_iter7_reg);

assign sub_ln703_345_fu_3234_p2 = (add_ln703_404_fu_3135_p2 - data_25_V_read26_reg_9677_pp0_iter7_reg);

assign sub_ln703_346_fu_3396_p2 = (add_ln703_410_reg_11287 - data_25_V_read26_reg_9677_pp0_iter8_reg);

assign sub_ln703_347_fu_3400_p2 = (sub_ln703_332_fu_3376_p2 - data_25_V_read26_reg_9677_pp0_iter8_reg);

assign sub_ln703_348_fu_3405_p2 = (add_ln703_411_fu_3380_p2 - data_25_V_read26_reg_9677_pp0_iter8_reg);

assign sub_ln703_349_fu_3410_p2 = (sub_ln703_333_reg_11292 - data_25_V_read26_reg_9677_pp0_iter8_reg);

assign sub_ln703_34_fu_778_p2 = (sub_ln703_20_reg_10465 - data_5_V_read_9_reg_10245_pp0_iter3_reg);

assign sub_ln703_350_fu_3244_p2 = (add_ln703_413_fu_3160_p2 - data_25_V_read26_reg_9677_pp0_iter7_reg);

assign sub_ln703_351_fu_3414_p2 = (add_ln703_416_reg_11297 - data_25_V_read26_reg_9677_pp0_iter8_reg);

assign sub_ln703_352_fu_3427_p2 = (add_ln703_417_reg_11312 - data_25_V_read26_reg_9677_pp0_iter8_reg);

assign sub_ln703_353_fu_3269_p2 = (sub_ln703_337_fu_3190_p2 - data_25_V_read26_reg_9677_pp0_iter7_reg);

assign sub_ln703_354_fu_3431_p2 = (sub_ln703_339_reg_11317 - data_25_V_read26_reg_9677_pp0_iter8_reg);

assign sub_ln703_355_fu_3435_p2 = (sub_ln703_340_reg_11322 - data_25_V_read26_reg_9677_pp0_iter8_reg);

assign sub_ln703_356_fu_3290_p2 = (add_ln703_418_fu_3210_p2 - data_25_V_read26_reg_9677_pp0_iter7_reg);

assign sub_ln703_357_fu_3295_p2 = (add_ln703_421_fu_3229_p2 - data_25_V_read26_reg_9677_pp0_iter7_reg);

assign sub_ln703_358_fu_3300_p2 = (add_ln703_422_fu_3239_p2 - data_26_V_read27_reg_9652_pp0_iter7_reg);

assign sub_ln703_359_fu_3448_p2 = (sub_ln703_349_fu_3410_p2 - data_26_V_read27_reg_9652_pp0_iter8_reg);

assign sub_ln703_35_fu_787_p2 = (sub_ln703_23_reg_10471 - data_5_V_read_9_reg_10245_pp0_iter3_reg);

assign sub_ln703_360_fu_3453_p2 = (sub_ln703_350_reg_11342 - data_26_V_read27_reg_9652_pp0_iter8_reg);

assign sub_ln703_361_fu_3457_p2 = (add_ln703_426_reg_11347 - data_26_V_read27_reg_9652_pp0_iter8_reg);

assign sub_ln703_362_fu_3305_p2 = (add_ln703_428_fu_3264_p2 - data_26_V_read27_reg_9652_pp0_iter7_reg);

assign sub_ln703_363_fu_3461_p2 = (add_ln703_429_fu_3418_p2 - data_26_V_read27_reg_9652_pp0_iter8_reg);

assign sub_ln703_364_fu_3470_p2 = (add_ln703_430_fu_3423_p2 - data_26_V_read27_reg_9652_pp0_iter8_reg);

assign sub_ln703_365_fu_3475_p2 = (sub_ln703_352_fu_3427_p2 - data_26_V_read27_reg_9652_pp0_iter8_reg);

assign sub_ln703_366_fu_3484_p2 = (add_ln703_431_reg_11357 - data_26_V_read27_reg_9652_pp0_iter8_reg);

assign sub_ln703_367_fu_3488_p2 = (sub_ln703_354_fu_3431_p2 - data_26_V_read27_reg_9652_pp0_iter8_reg);

assign sub_ln703_368_fu_3493_p2 = (add_ln703_435_reg_11362 - data_26_V_read27_reg_9652_pp0_iter8_reg);

assign sub_ln703_369_fu_3497_p2 = (sub_ln703_355_fu_3435_p2 - data_26_V_read27_reg_9652_pp0_iter8_reg);

assign sub_ln703_36_fu_795_p2 = (add_ln703_138_fu_701_p2 - data_5_V_read_9_reg_10245_pp0_iter3_reg);

assign sub_ln703_370_fu_3515_p2 = (add_ln703_436_fu_3439_p2 - data_26_V_read27_reg_9652_pp0_iter8_reg);

assign sub_ln703_371_fu_3324_p2 = (sub_ln703_357_fu_3295_p2 - data_26_V_read27_reg_9652_pp0_iter7_reg);

assign sub_ln703_372_fu_3532_p2 = (add_ln703_437_fu_3443_p2 - data_27_V_read28_reg_9625_pp0_iter8_reg);

assign sub_ln703_373_fu_3547_p2 = (sub_ln703_360_fu_3453_p2 - data_27_V_read28_reg_9625_pp0_iter8_reg);

assign sub_ln703_374_fu_3566_p2 = (add_ln703_440_fu_3466_p2 - data_27_V_read28_reg_9625_pp0_iter8_reg);

assign sub_ln703_375_fu_3576_p2 = (add_ln703_441_fu_3480_p2 - data_27_V_read28_reg_9625_pp0_iter8_reg);

assign sub_ln703_376_fu_3591_p2 = (sub_ln703_368_fu_3493_p2 - data_27_V_read28_reg_9625_pp0_iter8_reg);

assign sub_ln703_377_fu_3596_p2 = (sub_ln703_369_fu_3497_p2 - data_27_V_read28_reg_9625_pp0_iter8_reg);

assign sub_ln703_378_fu_3601_p2 = (add_ln703_442_fu_3502_p2 - data_27_V_read28_reg_9625_pp0_iter8_reg);

assign sub_ln703_379_fu_3606_p2 = (add_ln703_444_fu_3506_p2 - data_27_V_read28_reg_9625_pp0_iter8_reg);

assign sub_ln703_37_fu_800_p2 = (sub_ln703_17_reg_10453 - data_5_V_read_9_reg_10245_pp0_iter3_reg);

assign sub_ln703_380_fu_3611_p2 = (add_ln703_448_fu_3511_p2 - data_27_V_read28_reg_9625_pp0_iter8_reg);

assign sub_ln703_381_fu_3616_p2 = (sub_ln703_370_fu_3515_p2 - data_27_V_read28_reg_9625_pp0_iter8_reg);

assign sub_ln703_382_fu_3621_p2 = (add_ln703_450_fu_3520_p2 - data_27_V_read28_reg_9625_pp0_iter8_reg);

assign sub_ln703_383_fu_3626_p2 = (sub_ln703_371_reg_11397 - data_27_V_read28_reg_9625_pp0_iter8_reg);

assign sub_ln703_384_fu_3645_p2 = (add_ln703_452_fu_3524_p2 - data_28_V_read_8_reg_9598_pp0_iter8_reg);

assign sub_ln703_385_fu_3650_p2 = (add_ln703_453_fu_3528_p2 - data_28_V_read_8_reg_9598_pp0_iter8_reg);

assign sub_ln703_386_fu_3660_p2 = (add_ln703_455_fu_3537_p2 - data_28_V_read_8_reg_9598_pp0_iter8_reg);

assign sub_ln703_387_fu_3665_p2 = (add_ln703_456_fu_3542_p2 - data_28_V_read_8_reg_9598_pp0_iter8_reg);

assign sub_ln703_388_fu_3670_p2 = (add_ln703_458_fu_3552_p2 - data_28_V_read_8_reg_9598_pp0_iter8_reg);

assign sub_ln703_389_fu_3675_p2 = (add_ln703_461_fu_3561_p2 - data_28_V_read_8_reg_9598_pp0_iter8_reg);

assign sub_ln703_38_fu_814_p2 = (sub_ln703_27_fu_732_p2 - data_6_V_read_9_reg_10218_pp0_iter3_reg);

assign sub_ln703_390_fu_3690_p2 = (add_ln703_462_fu_3571_p2 - data_28_V_read_8_reg_9598_pp0_iter8_reg);

assign sub_ln703_391_fu_3695_p2 = (sub_ln703_375_fu_3576_p2 - data_28_V_read_8_reg_9598_pp0_iter8_reg);

assign sub_ln703_392_fu_3700_p2 = (add_ln703_463_fu_3581_p2 - data_28_V_read_8_reg_9598_pp0_iter8_reg);

assign sub_ln703_393_fu_3705_p2 = (add_ln703_464_fu_3586_p2 - data_28_V_read_8_reg_9598_pp0_iter8_reg);

assign sub_ln703_394_fu_3710_p2 = (sub_ln703_377_fu_3596_p2 - data_28_V_read_8_reg_9598_pp0_iter8_reg);

assign sub_ln703_395_fu_3720_p2 = (sub_ln703_379_fu_3606_p2 - data_28_V_read_8_reg_9598_pp0_iter8_reg);

assign sub_ln703_396_fu_3725_p2 = (sub_ln703_380_fu_3611_p2 - data_28_V_read_8_reg_9598_pp0_iter8_reg);

assign sub_ln703_397_fu_3746_p2 = (sub_ln703_382_fu_3621_p2 - data_28_V_read_8_reg_9598_pp0_iter8_reg);

assign sub_ln703_398_fu_3751_p2 = (sub_ln703_383_fu_3626_p2 - data_28_V_read_8_reg_9598_pp0_iter8_reg);

assign sub_ln703_399_fu_3761_p2 = (add_ln703_468_fu_3639_p2 - data_29_V_read_8_reg_9573_pp0_iter8_reg);

assign sub_ln703_39_fu_819_p2 = (add_ln703_145_fu_736_p2 - data_6_V_read_9_reg_10218_pp0_iter3_reg);

assign sub_ln703_3_fu_560_p2 = (sub_ln703_1_reg_10348 - data_2_V_read_10_reg_10312_pp0_iter1_reg);

assign sub_ln703_400_fu_3973_p2 = (add_ln703_469_reg_11479 - data_29_V_read_8_reg_9573_pp0_iter9_reg);

assign sub_ln703_401_fu_3781_p2 = (sub_ln703_388_fu_3670_p2 - data_29_V_read_8_reg_9573_pp0_iter8_reg);

assign sub_ln703_402_fu_3786_p2 = (sub_ln703_389_fu_3675_p2 - data_29_V_read_8_reg_9573_pp0_iter8_reg);

assign sub_ln703_403_fu_3791_p2 = (add_ln703_474_fu_3680_p2 - data_29_V_read_8_reg_9573_pp0_iter8_reg);

assign sub_ln703_404_fu_3977_p2 = (add_ln703_476_reg_11494 - data_29_V_read_8_reg_9573_pp0_iter9_reg);

assign sub_ln703_405_fu_3816_p2 = (sub_ln703_392_fu_3700_p2 - data_29_V_read_8_reg_9573_pp0_iter8_reg);

assign sub_ln703_406_fu_3981_p2 = (sub_ln703_393_reg_11504 - data_29_V_read_8_reg_9573_pp0_iter9_reg);

assign sub_ln703_407_fu_3985_p2 = (sub_ln703_394_reg_11509 - data_29_V_read_8_reg_9573_pp0_iter9_reg);

assign sub_ln703_408_fu_3845_p2 = (add_ln703_477_fu_3715_p2 - data_29_V_read_8_reg_9573_pp0_iter8_reg);

assign sub_ln703_409_fu_3989_p2 = (sub_ln703_395_reg_11514 - data_29_V_read_8_reg_9573_pp0_iter9_reg);

assign sub_ln703_40_fu_824_p2 = (add_ln703_146_fu_741_p2 - data_6_V_read_9_reg_10218_pp0_iter3_reg);

assign sub_ln703_410_fu_3993_p2 = (add_ln703_478_reg_11519 - data_29_V_read_8_reg_9573_pp0_iter9_reg);

assign sub_ln703_411_fu_3850_p2 = (add_ln703_482_fu_3740_p2 - data_29_V_read_8_reg_9573_pp0_iter8_reg);

assign sub_ln703_412_fu_3855_p2 = (add_ln703_487_fu_3756_p2 - data_29_V_read_8_reg_9573_pp0_iter8_reg);

assign sub_ln703_413_fu_3997_p2 = (sub_ln703_399_reg_11524 - data_30_V_read31_reg_9549_pp0_iter9_reg);

assign sub_ln703_414_fu_3860_p2 = (add_ln703_488_fu_3766_p2 - data_30_V_read31_reg_9549_pp0_iter8_reg);

assign sub_ln703_415_fu_4001_p2 = (sub_ln703_400_fu_3973_p2 - data_30_V_read31_reg_9549_pp0_iter9_reg);

assign sub_ln703_416_fu_3865_p2 = (add_ln703_491_fu_3776_p2 - data_30_V_read31_reg_9549_pp0_iter8_reg);

assign sub_ln703_417_fu_4010_p2 = (sub_ln703_402_reg_11534 - data_30_V_read31_reg_9549_pp0_iter9_reg);

assign sub_ln703_418_fu_4014_p2 = (sub_ln703_404_fu_3977_p2 - data_30_V_read31_reg_9549_pp0_iter9_reg);

assign sub_ln703_419_fu_3884_p2 = (add_ln703_493_fu_3796_p2 - data_30_V_read31_reg_9549_pp0_iter8_reg);

assign sub_ln703_41_fu_829_p2 = (sub_ln703_28_reg_10476 - data_6_V_read_9_reg_10218_pp0_iter3_reg);

assign sub_ln703_420_fu_4019_p2 = (add_ln703_496_reg_11544 - data_30_V_read31_reg_9549_pp0_iter9_reg);

assign sub_ln703_421_fu_4023_p2 = (add_ln703_497_reg_11549 - data_30_V_read31_reg_9549_pp0_iter9_reg);

assign sub_ln703_422_fu_4027_p2 = (sub_ln703_405_reg_11554 - data_30_V_read31_reg_9549_pp0_iter9_reg);

assign sub_ln703_423_fu_4031_p2 = (add_ln703_506_reg_11559 - data_30_V_read31_reg_9549_pp0_iter9_reg);

assign sub_ln703_424_fu_4040_p2 = (sub_ln703_408_reg_11564 - data_30_V_read31_reg_9549_pp0_iter9_reg);

assign sub_ln703_425_fu_4044_p2 = (sub_ln703_409_fu_3989_p2 - data_30_V_read31_reg_9549_pp0_iter9_reg);

assign sub_ln703_426_fu_4049_p2 = (sub_ln703_410_fu_3993_p2 - data_30_V_read31_reg_9549_pp0_iter9_reg);

assign sub_ln703_427_fu_4054_p2 = (sub_ln703_411_reg_11569 - data_30_V_read31_reg_9549_pp0_iter9_reg);

assign sub_ln703_428_fu_4080_p2 = (add_ln703_508_fu_4006_p2 - data_31_V_read32_reg_9521_pp0_iter9_reg);

assign sub_ln703_429_fu_4102_p2 = (add_ln703_512_reg_11589 - data_31_V_read32_reg_9521_pp0_iter9_reg);

assign sub_ln703_42_fu_833_p2 = (add_ln703_147_fu_745_p2 - data_6_V_read_9_reg_10218_pp0_iter3_reg);

assign sub_ln703_430_fu_4106_p2 = (sub_ln703_417_fu_4010_p2 - data_31_V_read32_reg_9521_pp0_iter9_reg);

assign sub_ln703_431_fu_4120_p2 = (sub_ln703_419_reg_11594 - data_31_V_read32_reg_9521_pp0_iter9_reg);

assign sub_ln703_432_fu_4124_p2 = (sub_ln703_420_fu_4019_p2 - data_31_V_read32_reg_9521_pp0_iter9_reg);

assign sub_ln703_433_fu_4129_p2 = (sub_ln703_421_fu_4023_p2 - data_31_V_read32_reg_9521_pp0_iter9_reg);

assign sub_ln703_434_fu_4134_p2 = (sub_ln703_422_fu_4027_p2 - data_31_V_read32_reg_9521_pp0_iter9_reg);

assign sub_ln703_435_fu_4144_p2 = (add_ln703_513_fu_4035_p2 - data_31_V_read32_reg_9521_pp0_iter9_reg);

assign sub_ln703_436_fu_4149_p2 = (sub_ln703_424_fu_4040_p2 - data_31_V_read32_reg_9521_pp0_iter9_reg);

assign sub_ln703_437_fu_4154_p2 = (add_ln703_515_reg_11599 - data_31_V_read32_reg_9521_pp0_iter9_reg);

assign sub_ln703_438_fu_4163_p2 = (sub_ln703_427_fu_4054_p2 - data_31_V_read32_reg_9521_pp0_iter9_reg);

assign sub_ln703_439_fu_4168_p2 = (add_ln703_517_reg_11604 - data_31_V_read32_reg_9521_pp0_iter9_reg);

assign sub_ln703_43_fu_838_p2 = (sub_ln703_29_fu_749_p2 - data_6_V_read_9_reg_10218_pp0_iter3_reg);

assign sub_ln703_440_fu_3938_p2 = (add_ln703_519_fu_3899_p2 - data_31_V_read32_reg_9521_pp0_iter8_reg);

assign sub_ln703_441_fu_4172_p2 = (add_ln703_520_fu_4058_p2 - data_31_V_read32_reg_9521_pp0_iter9_reg);

assign sub_ln703_442_fu_4177_p2 = (add_ln703_521_fu_4062_p2 - data_32_V_read_3_reg_9492_pp0_iter9_reg);

assign sub_ln703_443_fu_4182_p2 = (add_ln703_522_fu_4067_p2 - data_32_V_read_3_reg_9492_pp0_iter9_reg);

assign sub_ln703_444_fu_4187_p2 = (add_ln703_538_fu_4075_p2 - data_32_V_read_3_reg_9492_pp0_iter9_reg);

assign sub_ln703_445_fu_4192_p2 = (sub_ln703_428_fu_4080_p2 - data_32_V_read_3_reg_9492_pp0_iter9_reg);

assign sub_ln703_446_fu_4197_p2 = (add_ln703_541_fu_4089_p2 - data_32_V_read_3_reg_9492_pp0_iter9_reg);

assign sub_ln703_447_fu_4202_p2 = (add_ln703_545_reg_11614 - data_32_V_read_3_reg_9492_pp0_iter9_reg);

assign sub_ln703_448_fu_4206_p2 = (add_ln703_546_fu_4094_p2 - data_32_V_read_3_reg_9492_pp0_iter9_reg);

assign sub_ln703_449_fu_4211_p2 = (add_ln703_548_fu_4098_p2 - data_32_V_read_3_reg_9492_pp0_iter9_reg);

assign sub_ln703_44_fu_848_p2 = (add_ln703_148_fu_757_p2 - data_6_V_read_9_reg_10218_pp0_iter3_reg);

assign sub_ln703_450_fu_4221_p2 = (sub_ln703_430_fu_4106_p2 - data_32_V_read_3_reg_9492_pp0_iter9_reg);

assign sub_ln703_451_fu_4226_p2 = (add_ln703_550_fu_4111_p2 - data_32_V_read_3_reg_9492_pp0_iter9_reg);

assign sub_ln703_452_fu_4231_p2 = (add_ln703_551_fu_4115_p2 - data_32_V_read_3_reg_9492_pp0_iter9_reg);

assign sub_ln703_453_fu_4236_p2 = (sub_ln703_431_fu_4120_p2 - data_32_V_read_3_reg_9492_pp0_iter9_reg);

assign sub_ln703_454_fu_4246_p2 = (add_ln703_552_fu_4139_p2 - data_32_V_read_3_reg_9492_pp0_iter9_reg);

assign sub_ln703_455_fu_4251_p2 = (add_ln703_556_reg_11619 - data_32_V_read_3_reg_9492_pp0_iter9_reg);

assign sub_ln703_456_fu_4255_p2 = (sub_ln703_436_fu_4149_p2 - data_32_V_read_3_reg_9492_pp0_iter9_reg);

assign sub_ln703_457_fu_4265_p2 = (sub_ln703_437_fu_4154_p2 - data_32_V_read_3_reg_9492_pp0_iter9_reg);

assign sub_ln703_458_fu_4270_p2 = (add_ln703_557_fu_4158_p2 - data_32_V_read_3_reg_9492_pp0_iter9_reg);

assign sub_ln703_459_fu_4284_p2 = (sub_ln703_441_fu_4172_p2 - data_32_V_read_3_reg_9492_pp0_iter9_reg);

assign sub_ln703_45_fu_853_p2 = (sub_ln703_31_fu_761_p2 - data_6_V_read_9_reg_10218_pp0_iter3_reg);

assign sub_ln703_460_fu_4289_p2 = (sub_ln703_443_fu_4182_p2 - data_33_V_read_3_reg_9463_pp0_iter9_reg);

assign sub_ln703_461_fu_4303_p2 = (sub_ln703_445_fu_4192_p2 - data_33_V_read_3_reg_9463_pp0_iter9_reg);

assign sub_ln703_462_fu_4313_p2 = (sub_ln703_447_fu_4202_p2 - data_33_V_read_3_reg_9463_pp0_iter9_reg);

assign sub_ln703_463_fu_4558_p2 = (sub_ln703_448_reg_11673 - data_33_V_read_3_reg_9463_pp0_iter10_reg);

assign sub_ln703_464_fu_4318_p2 = (add_ln703_558_fu_4216_p2 - data_33_V_read_3_reg_9463_pp0_iter9_reg);

assign sub_ln703_465_fu_4328_p2 = (sub_ln703_451_fu_4226_p2 - data_33_V_read_3_reg_9463_pp0_iter9_reg);

assign sub_ln703_466_fu_4562_p2 = (sub_ln703_452_reg_11678 - data_33_V_read_3_reg_9463_pp0_iter10_reg);

assign sub_ln703_467_fu_4333_p2 = (add_ln703_559_fu_4241_p2 - data_33_V_read_3_reg_9463_pp0_iter9_reg);

assign sub_ln703_468_fu_4353_p2 = (sub_ln703_454_fu_4246_p2 - data_33_V_read_3_reg_9463_pp0_iter9_reg);

assign sub_ln703_469_fu_4368_p2 = (sub_ln703_456_fu_4255_p2 - data_33_V_read_3_reg_9463_pp0_iter9_reg);

assign sub_ln703_46_fu_858_p2 = (sub_ln703_32_fu_765_p2 - data_6_V_read_9_reg_10218_pp0_iter3_reg);

assign sub_ln703_470_fu_4373_p2 = (add_ln703_561_fu_4260_p2 - data_33_V_read_3_reg_9463_pp0_iter9_reg);

assign sub_ln703_471_fu_4378_p2 = (sub_ln703_457_fu_4265_p2 - data_33_V_read_3_reg_9463_pp0_iter9_reg);

assign sub_ln703_472_fu_4570_p2 = (sub_ln703_458_reg_11688 - data_33_V_read_3_reg_9463_pp0_iter10_reg);

assign sub_ln703_473_fu_4388_p2 = (add_ln703_562_fu_4275_p2 - data_33_V_read_3_reg_9463_pp0_iter9_reg);

assign sub_ln703_474_fu_4393_p2 = (add_ln703_563_fu_4280_p2 - data_33_V_read_3_reg_9463_pp0_iter9_reg);

assign sub_ln703_475_fu_4418_p2 = (add_ln703_571_fu_4298_p2 - data_34_V_read_3_reg_9434_pp0_iter9_reg);

assign sub_ln703_476_fu_4574_p2 = (sub_ln703_461_reg_11693 - data_34_V_read_3_reg_9434_pp0_iter10_reg);

assign sub_ln703_477_fu_4578_p2 = (add_ln703_572_reg_11698 - data_34_V_read_3_reg_9434_pp0_iter10_reg);

assign sub_ln703_478_fu_4582_p2 = (sub_ln703_462_reg_11703 - data_34_V_read_3_reg_9434_pp0_iter10_reg);

assign sub_ln703_479_fu_4586_p2 = (add_ln703_573_reg_11708 - data_34_V_read_3_reg_9434_pp0_iter10_reg);

assign sub_ln703_47_fu_863_p2 = (sub_ln703_33_fu_769_p2 - data_6_V_read_9_reg_10218_pp0_iter3_reg);

assign sub_ln703_480_fu_4590_p2 = (add_ln703_574_fu_4566_p2 - data_34_V_read_3_reg_9434_pp0_iter10_reg);

assign sub_ln703_481_fu_4595_p2 = (sub_ln703_467_reg_11713 - data_34_V_read_3_reg_9434_pp0_iter10_reg);

assign sub_ln703_482_fu_4447_p2 = (add_ln703_576_fu_4338_p2 - data_34_V_read_3_reg_9434_pp0_iter9_reg);

assign sub_ln703_483_fu_4452_p2 = (add_ln703_580_fu_4348_p2 - data_34_V_read_3_reg_9434_pp0_iter9_reg);

assign sub_ln703_484_fu_4599_p2 = (sub_ln703_468_reg_11718 - data_34_V_read_3_reg_9434_pp0_iter10_reg);

assign sub_ln703_485_fu_4603_p2 = (add_ln703_581_reg_11723 - data_34_V_read_3_reg_9434_pp0_iter10_reg);

assign sub_ln703_486_fu_4607_p2 = (add_ln703_583_reg_11728 - data_34_V_read_3_reg_9434_pp0_iter10_reg);

assign sub_ln703_487_fu_4611_p2 = (sub_ln703_470_reg_11738 - data_34_V_read_3_reg_9434_pp0_iter10_reg);

assign sub_ln703_488_fu_4457_p2 = (sub_ln703_471_fu_4378_p2 - data_34_V_read_3_reg_9434_pp0_iter9_reg);

assign sub_ln703_489_fu_4615_p2 = (sub_ln703_472_fu_4570_p2 - data_34_V_read_3_reg_9434_pp0_iter10_reg);

assign sub_ln703_48_fu_877_p2 = (add_ln703_149_fu_773_p2 - data_6_V_read_9_reg_10218_pp0_iter3_reg);

assign sub_ln703_490_fu_4462_p2 = (add_ln703_585_fu_4383_p2 - data_34_V_read_3_reg_9434_pp0_iter9_reg);

assign sub_ln703_491_fu_4467_p2 = (sub_ln703_473_fu_4388_p2 - data_34_V_read_3_reg_9434_pp0_iter9_reg);

assign sub_ln703_492_fu_4472_p2 = (sub_ln703_474_fu_4393_p2 - data_34_V_read_3_reg_9434_pp0_iter9_reg);

assign sub_ln703_493_fu_4624_p2 = (add_ln703_586_reg_11743 - data_35_V_read_3_reg_9410_pp0_iter10_reg);

assign sub_ln703_494_fu_4632_p2 = (add_ln703_590_reg_11748 - data_35_V_read_3_reg_9410_pp0_iter10_reg);

assign sub_ln703_495_fu_4636_p2 = (sub_ln703_475_reg_11753 - data_35_V_read_3_reg_9410_pp0_iter10_reg);

assign sub_ln703_496_fu_4650_p2 = (add_ln703_591_reg_11758 - data_35_V_read_3_reg_9410_pp0_iter10_reg);

assign sub_ln703_497_fu_4654_p2 = (sub_ln703_479_fu_4586_p2 - data_35_V_read_3_reg_9410_pp0_iter10_reg);

assign sub_ln703_498_fu_4659_p2 = (add_ln703_592_reg_11763 - data_35_V_read_3_reg_9410_pp0_iter10_reg);

assign sub_ln703_499_fu_4663_p2 = (sub_ln703_480_fu_4590_p2 - data_35_V_read_3_reg_9410_pp0_iter10_reg);

assign sub_ln703_49_fu_882_p2 = (sub_ln703_34_fu_778_p2 - data_6_V_read_9_reg_10218_pp0_iter3_reg);

assign sub_ln703_4_fu_548_p2 = (add_ln703_reg_10335 - data_2_V_read_10_reg_10312);

assign sub_ln703_500_fu_4668_p2 = (add_ln703_598_reg_11768 - data_35_V_read_3_reg_9410_pp0_iter10_reg);

assign sub_ln703_501_fu_4672_p2 = (sub_ln703_481_fu_4595_p2 - data_35_V_read_3_reg_9410_pp0_iter10_reg);

assign sub_ln703_502_fu_4682_p2 = (sub_ln703_485_fu_4603_p2 - data_35_V_read_3_reg_9410_pp0_iter10_reg);

assign sub_ln703_503_fu_4516_p2 = (sub_ln703_492_fu_4472_p2 - data_35_V_read_3_reg_9410_pp0_iter9_reg);

assign sub_ln703_504_fu_4700_p2 = (add_ln703_601_fu_4620_p2 - data_36_V_read_3_reg_9383_pp0_iter10_reg);

assign sub_ln703_505_fu_4521_p2 = (add_ln703_608_fu_4495_p2 - data_36_V_read_3_reg_9383_pp0_iter9_reg);

assign sub_ln703_506_fu_4705_p2 = (sub_ln703_493_fu_4624_p2 - data_36_V_read_3_reg_9383_pp0_iter10_reg);

assign sub_ln703_507_fu_4710_p2 = (add_ln703_611_fu_4628_p2 - data_36_V_read_3_reg_9383_pp0_iter10_reg);

assign sub_ln703_508_fu_4715_p2 = (sub_ln703_494_fu_4632_p2 - data_36_V_read_3_reg_9383_pp0_iter10_reg);

assign sub_ln703_509_fu_4725_p2 = (add_ln703_612_fu_4640_p2 - data_36_V_read_3_reg_9383_pp0_iter10_reg);

assign sub_ln703_50_fu_887_p2 = (add_ln703_150_fu_782_p2 - data_6_V_read_9_reg_10218_pp0_iter3_reg);

assign sub_ln703_510_fu_4730_p2 = (add_ln703_613_fu_4645_p2 - data_36_V_read_3_reg_9383_pp0_iter10_reg);

assign sub_ln703_511_fu_4735_p2 = (add_ln703_616_reg_11808 - data_36_V_read_3_reg_9383_pp0_iter10_reg);

assign sub_ln703_512_fu_4744_p2 = (sub_ln703_497_fu_4654_p2 - data_36_V_read_3_reg_9383_pp0_iter10_reg);

assign sub_ln703_513_fu_4749_p2 = (sub_ln703_498_fu_4659_p2 - data_36_V_read_3_reg_9383_pp0_iter10_reg);

assign sub_ln703_514_fu_4764_p2 = (sub_ln703_500_fu_4668_p2 - data_36_V_read_3_reg_9383_pp0_iter10_reg);

assign sub_ln703_515_fu_4778_p2 = (add_ln703_617_fu_4677_p2 - data_36_V_read_3_reg_9383_pp0_iter10_reg);

assign sub_ln703_516_fu_4783_p2 = (sub_ln703_502_fu_4682_p2 - data_36_V_read_3_reg_9383_pp0_iter10_reg);

assign sub_ln703_517_fu_4788_p2 = (add_ln703_618_fu_4687_p2 - data_36_V_read_3_reg_9383_pp0_iter10_reg);

assign sub_ln703_518_fu_4798_p2 = (add_ln703_619_fu_4692_p2 - data_36_V_read_3_reg_9383_pp0_iter10_reg);

assign sub_ln703_519_fu_4808_p2 = (add_ln703_620_fu_4696_p2 - data_36_V_read_3_reg_9383_pp0_iter10_reg);

assign sub_ln703_51_fu_897_p2 = (add_ln703_151_fu_791_p2 - data_6_V_read_9_reg_10218_pp0_iter3_reg);

assign sub_ln703_520_fu_4813_p2 = (sub_ln703_503_reg_11813 - data_36_V_read_3_reg_9383_pp0_iter10_reg);

assign sub_ln703_521_fu_4830_p2 = (sub_ln703_506_fu_4705_p2 - data_37_V_read_3_reg_9353_pp0_iter10_reg);

assign sub_ln703_522_fu_4840_p2 = (sub_ln703_508_fu_4715_p2 - data_37_V_read_3_reg_9353_pp0_iter10_reg);

assign sub_ln703_523_fu_4845_p2 = (add_ln703_622_fu_4720_p2 - data_37_V_read_3_reg_9353_pp0_iter10_reg);

assign sub_ln703_524_fu_4850_p2 = (sub_ln703_511_fu_4735_p2 - data_37_V_read_3_reg_9353_pp0_iter10_reg);

assign sub_ln703_525_fu_4855_p2 = (add_ln703_623_fu_4739_p2 - data_37_V_read_3_reg_9353_pp0_iter10_reg);

assign sub_ln703_526_fu_4860_p2 = (sub_ln703_512_fu_4744_p2 - data_37_V_read_3_reg_9353_pp0_iter10_reg);

assign sub_ln703_527_fu_4865_p2 = (add_ln703_626_fu_4759_p2 - data_37_V_read_3_reg_9353_pp0_iter10_reg);

assign sub_ln703_528_fu_4875_p2 = (sub_ln703_514_fu_4764_p2 - data_37_V_read_3_reg_9353_pp0_iter10_reg);

assign sub_ln703_529_fu_4880_p2 = (add_ln703_627_fu_4769_p2 - data_37_V_read_3_reg_9353_pp0_iter10_reg);

assign sub_ln703_52_fu_907_p2 = (sub_ln703_37_fu_800_p2 - data_6_V_read_9_reg_10218_pp0_iter3_reg);

assign sub_ln703_530_fu_4885_p2 = (add_ln703_629_fu_4774_p2 - data_37_V_read_3_reg_9353_pp0_iter10_reg);

assign sub_ln703_531_fu_4890_p2 = (add_ln703_634_reg_11828 - data_37_V_read_3_reg_9353_pp0_iter10_reg);

assign sub_ln703_532_fu_4894_p2 = (sub_ln703_515_fu_4778_p2 - data_37_V_read_3_reg_9353_pp0_iter10_reg);

assign sub_ln703_533_fu_4904_p2 = (sub_ln703_517_fu_4788_p2 - data_37_V_read_3_reg_9353_pp0_iter10_reg);

assign sub_ln703_534_fu_4909_p2 = (add_ln703_636_fu_4793_p2 - data_37_V_read_3_reg_9353_pp0_iter10_reg);

assign sub_ln703_535_fu_4919_p2 = (add_ln703_638_fu_4803_p2 - data_37_V_read_3_reg_9353_pp0_iter10_reg);

assign sub_ln703_536_fu_4924_p2 = (sub_ln703_520_fu_4813_p2 - data_37_V_read_3_reg_9353_pp0_iter10_reg);

assign sub_ln703_537_fu_4929_p2 = (add_ln703_642_fu_4817_p2 - data_37_V_read_3_reg_9353_pp0_iter10_reg);

assign sub_ln703_538_fu_4934_p2 = (add_ln703_643_fu_4821_p2 - data_38_V_read_3_reg_9328_pp0_iter10_reg);

assign sub_ln703_539_fu_4939_p2 = (add_ln703_644_fu_4826_p2 - data_38_V_read_3_reg_9328_pp0_iter10_reg);

assign sub_ln703_53_fu_912_p2 = (add_ln703_152_fu_804_p2 - data_7_V_read_9_reg_10191_pp0_iter3_reg);

assign sub_ln703_540_fu_4944_p2 = (add_ln703_645_fu_4835_p2 - data_38_V_read_3_reg_9328_pp0_iter10_reg);

assign sub_ln703_541_fu_4949_p2 = (sub_ln703_522_fu_4840_p2 - data_38_V_read_3_reg_9328_pp0_iter10_reg);

assign sub_ln703_542_fu_4954_p2 = (sub_ln703_523_fu_4845_p2 - data_38_V_read_3_reg_9328_pp0_iter10_reg);

assign sub_ln703_543_fu_4979_p2 = (sub_ln703_524_fu_4850_p2 - data_38_V_read_3_reg_9328_pp0_iter10_reg);

assign sub_ln703_544_fu_4984_p2 = (sub_ln703_525_fu_4855_p2 - data_38_V_read_3_reg_9328_pp0_iter10_reg);

assign sub_ln703_545_fu_5138_p2 = (sub_ln703_526_reg_11864 - data_38_V_read_3_reg_9328_pp0_iter11_reg);

assign sub_ln703_546_fu_5142_p2 = (sub_ln703_527_reg_11869 - data_38_V_read_3_reg_9328_pp0_iter11_reg);

assign sub_ln703_547_fu_5146_p2 = (add_ln703_647_reg_11874 - data_38_V_read_3_reg_9328_pp0_iter11_reg);

assign sub_ln703_548_fu_5154_p2 = (sub_ln703_532_reg_11884 - data_38_V_read_3_reg_9328_pp0_iter11_reg);

assign sub_ln703_549_fu_5158_p2 = (add_ln703_648_reg_11889 - data_38_V_read_3_reg_9328_pp0_iter11_reg);

assign sub_ln703_54_fu_1086_p2 = (add_ln703_153_reg_10503 - data_7_V_read_9_reg_10191_pp0_iter4_reg);

assign sub_ln703_550_fu_5162_p2 = (sub_ln703_533_reg_11894 - data_38_V_read_3_reg_9328_pp0_iter11_reg);

assign sub_ln703_551_fu_5004_p2 = (add_ln703_649_fu_4914_p2 - data_38_V_read_3_reg_9328_pp0_iter10_reg);

assign sub_ln703_552_fu_5170_p2 = (sub_ln703_539_reg_11909 - data_39_V_read_3_reg_9301_pp0_iter11_reg);

assign sub_ln703_553_fu_5174_p2 = (sub_ln703_540_reg_11914 - data_39_V_read_3_reg_9301_pp0_iter11_reg);

assign sub_ln703_554_fu_5178_p2 = (sub_ln703_542_reg_11924 - data_39_V_read_3_reg_9301_pp0_iter11_reg);

assign sub_ln703_555_fu_5182_p2 = (add_ln703_651_reg_11929 - data_39_V_read_3_reg_9301_pp0_iter11_reg);

assign sub_ln703_556_fu_5024_p2 = (add_ln703_656_fu_4973_p2 - data_39_V_read_3_reg_9301_pp0_iter10_reg);

assign sub_ln703_557_fu_5029_p2 = (sub_ln703_543_fu_4979_p2 - data_39_V_read_3_reg_9301_pp0_iter10_reg);

assign sub_ln703_558_fu_5034_p2 = (add_ln703_658_fu_4989_p2 - data_39_V_read_3_reg_9301_pp0_iter10_reg);

assign sub_ln703_559_fu_5190_p2 = (sub_ln703_546_fu_5142_p2 - data_39_V_read_3_reg_9301_pp0_iter11_reg);

assign sub_ln703_55_fu_1090_p2 = (sub_ln703_38_reg_10508 - data_7_V_read_9_reg_10191_pp0_iter4_reg);

assign sub_ln703_560_fu_5195_p2 = (sub_ln703_547_fu_5146_p2 - data_39_V_read_3_reg_9301_pp0_iter11_reg);

assign sub_ln703_561_fu_5200_p2 = (add_ln703_659_fu_5150_p2 - data_39_V_read_3_reg_9301_pp0_iter11_reg);

assign sub_ln703_562_fu_5205_p2 = (add_ln703_660_reg_11939 - data_39_V_read_3_reg_9301_pp0_iter11_reg);

assign sub_ln703_563_fu_5209_p2 = (sub_ln703_548_fu_5154_p2 - data_39_V_read_3_reg_9301_pp0_iter11_reg);

assign sub_ln703_564_fu_5214_p2 = (sub_ln703_550_fu_5162_p2 - data_39_V_read_3_reg_9301_pp0_iter11_reg);

assign sub_ln703_565_fu_5219_p2 = (add_ln703_661_reg_11944 - data_39_V_read_3_reg_9301_pp0_iter11_reg);

assign sub_ln703_566_fu_5223_p2 = (sub_ln703_551_reg_11949 - data_39_V_read_3_reg_9301_pp0_iter11_reg);

assign sub_ln703_567_fu_5227_p2 = (add_ln703_662_fu_5166_p2 - data_39_V_read_3_reg_9301_pp0_iter11_reg);

assign sub_ln703_568_fu_5232_p2 = (add_ln703_666_reg_11954 - data_39_V_read_3_reg_9301_pp0_iter11_reg);

assign sub_ln703_569_fu_5236_p2 = (add_ln703_668_reg_11959 - data_40_V_read41_reg_9272_pp0_iter11_reg);

assign sub_ln703_56_fu_1094_p2 = (sub_ln703_39_reg_10513 - data_7_V_read_9_reg_10191_pp0_iter4_reg);

assign sub_ln703_570_fu_5263_p2 = (sub_ln703_557_reg_11969 - data_40_V_read41_reg_9272_pp0_iter11_reg);

assign sub_ln703_571_fu_5267_p2 = (add_ln703_669_fu_5186_p2 - data_40_V_read41_reg_9272_pp0_iter11_reg);

assign sub_ln703_572_fu_5276_p2 = (sub_ln703_560_fu_5195_p2 - data_40_V_read41_reg_9272_pp0_iter11_reg);

assign sub_ln703_573_fu_5101_p2 = (add_ln703_671_fu_5039_p2 - data_40_V_read41_reg_9272_pp0_iter10_reg);

assign sub_ln703_574_fu_5290_p2 = (sub_ln703_562_fu_5205_p2 - data_40_V_read41_reg_9272_pp0_iter11_reg);

assign sub_ln703_575_fu_5295_p2 = (add_ln703_676_reg_11979 - data_40_V_read41_reg_9272_pp0_iter11_reg);

assign sub_ln703_576_fu_5299_p2 = (sub_ln703_564_fu_5214_p2 - data_40_V_read41_reg_9272_pp0_iter11_reg);

assign sub_ln703_577_fu_5304_p2 = (add_ln703_682_reg_11984 - data_40_V_read41_reg_9272_pp0_iter11_reg);

assign sub_ln703_578_fu_5308_p2 = (sub_ln703_565_fu_5219_p2 - data_40_V_read41_reg_9272_pp0_iter11_reg);

assign sub_ln703_579_fu_5318_p2 = (sub_ln703_567_fu_5227_p2 - data_40_V_read41_reg_9272_pp0_iter11_reg);

assign sub_ln703_57_fu_1102_p2 = (sub_ln703_40_reg_10519 - data_7_V_read_9_reg_10191_pp0_iter4_reg);

assign sub_ln703_580_fu_5323_p2 = (sub_ln703_568_fu_5232_p2 - data_40_V_read41_reg_9272_pp0_iter11_reg);

assign sub_ln703_581_fu_5328_p2 = (add_ln703_685_reg_11989 - data_40_V_read41_reg_9272_pp0_iter11_reg);

assign sub_ln703_582_fu_5106_p2 = (add_ln703_687_fu_5082_p2 - data_40_V_read41_reg_9272_pp0_iter10_reg);

assign sub_ln703_583_fu_5111_p2 = (add_ln703_689_fu_5087_p2 - data_40_V_read41_reg_9272_pp0_iter10_reg);

assign sub_ln703_584_fu_5341_p2 = (sub_ln703_569_fu_5236_p2 - data_41_V_read42_reg_9242_pp0_iter11_reg);

assign sub_ln703_585_fu_5346_p2 = (add_ln703_690_fu_5240_p2 - data_41_V_read42_reg_9242_pp0_iter11_reg);

assign sub_ln703_586_fu_5351_p2 = (add_ln703_692_fu_5245_p2 - data_41_V_read42_reg_9242_pp0_iter11_reg);

assign sub_ln703_587_fu_5356_p2 = (add_ln703_693_fu_5249_p2 - data_41_V_read42_reg_9242_pp0_iter11_reg);

assign sub_ln703_588_fu_5370_p2 = (add_ln703_694_fu_5254_p2 - data_41_V_read42_reg_9242_pp0_iter11_reg);

assign sub_ln703_589_fu_5375_p2 = (add_ln703_695_fu_5259_p2 - data_41_V_read42_reg_9242_pp0_iter11_reg);

assign sub_ln703_58_fu_922_p2 = (sub_ln703_41_fu_829_p2 - data_7_V_read_9_reg_10191_pp0_iter3_reg);

assign sub_ln703_590_fu_5380_p2 = (sub_ln703_570_fu_5263_p2 - data_41_V_read42_reg_9242_pp0_iter11_reg);

assign sub_ln703_591_fu_5385_p2 = (sub_ln703_571_fu_5267_p2 - data_41_V_read42_reg_9242_pp0_iter11_reg);

assign sub_ln703_592_fu_5400_p2 = (add_ln703_696_fu_5272_p2 - data_41_V_read42_reg_9242_pp0_iter11_reg);

assign sub_ln703_593_fu_5410_p2 = (sub_ln703_572_fu_5276_p2 - data_41_V_read42_reg_9242_pp0_iter11_reg);

assign sub_ln703_594_fu_5415_p2 = (add_ln703_699_fu_5281_p2 - data_41_V_read42_reg_9242_pp0_iter11_reg);

assign sub_ln703_595_fu_5420_p2 = (add_ln703_700_fu_5285_p2 - data_41_V_read42_reg_9242_pp0_iter11_reg);

assign sub_ln703_596_fu_5444_p2 = (sub_ln703_577_fu_5304_p2 - data_41_V_read42_reg_9242_pp0_iter11_reg);

assign sub_ln703_597_fu_5449_p2 = (add_ln703_701_fu_5313_p2 - data_41_V_read42_reg_9242_pp0_iter11_reg);

assign sub_ln703_598_fu_5454_p2 = (sub_ln703_579_fu_5318_p2 - data_41_V_read42_reg_9242_pp0_iter11_reg);

assign sub_ln703_599_fu_5459_p2 = (sub_ln703_580_fu_5323_p2 - data_41_V_read42_reg_9242_pp0_iter11_reg);

assign sub_ln703_59_fu_1106_p2 = (sub_ln703_43_reg_10524 - data_7_V_read_9_reg_10191_pp0_iter4_reg);

assign sub_ln703_5_fu_564_p2 = (data_2_V_read_10_reg_10312_pp0_iter1_reg - add_ln703_reg_10335_pp0_iter1_reg);

assign sub_ln703_600_fu_5464_p2 = (sub_ln703_581_fu_5328_p2 - data_41_V_read42_reg_9242_pp0_iter11_reg);

assign sub_ln703_601_fu_5473_p2 = (sub_ln703_583_reg_12017 - data_41_V_read42_reg_9242_pp0_iter11_reg);

assign sub_ln703_602_fu_5688_p2 = (add_ln703_704_reg_12056 - data_42_V_read_3_reg_9212_pp0_iter12_reg);

assign sub_ln703_603_fu_5491_p2 = (sub_ln703_587_fu_5356_p2 - data_42_V_read_3_reg_9212_pp0_iter11_reg);

assign sub_ln703_604_fu_5496_p2 = (add_ln703_709_fu_5365_p2 - data_42_V_read_3_reg_9212_pp0_iter11_reg);

assign sub_ln703_605_fu_5501_p2 = (sub_ln703_588_fu_5370_p2 - data_42_V_read_3_reg_9212_pp0_iter11_reg);

assign sub_ln703_606_fu_5696_p2 = (sub_ln703_589_reg_12066 - data_42_V_read_3_reg_9212_pp0_iter12_reg);

assign sub_ln703_607_fu_5506_p2 = (sub_ln703_590_fu_5380_p2 - data_42_V_read_3_reg_9212_pp0_iter11_reg);

assign sub_ln703_608_fu_5511_p2 = (sub_ln703_591_fu_5385_p2 - data_42_V_read_3_reg_9212_pp0_iter11_reg);

assign sub_ln703_609_fu_5516_p2 = (add_ln703_712_fu_5395_p2 - data_42_V_read_3_reg_9212_pp0_iter11_reg);

assign sub_ln703_60_fu_927_p2 = (add_ln703_154_fu_843_p2 - data_7_V_read_9_reg_10191_pp0_iter3_reg);

assign sub_ln703_610_fu_5521_p2 = (add_ln703_714_fu_5405_p2 - data_42_V_read_3_reg_9212_pp0_iter11_reg);

assign sub_ln703_611_fu_5704_p2 = (sub_ln703_594_reg_12076 - data_42_V_read_3_reg_9212_pp0_iter12_reg);

assign sub_ln703_612_fu_5526_p2 = (add_ln703_715_fu_5425_p2 - data_42_V_read_3_reg_9212_pp0_iter11_reg);

assign sub_ln703_613_fu_5531_p2 = (add_ln703_716_fu_5429_p2 - data_42_V_read_3_reg_9212_pp0_iter11_reg);

assign sub_ln703_614_fu_5536_p2 = (add_ln703_718_fu_5434_p2 - data_42_V_read_3_reg_9212_pp0_iter11_reg);

assign sub_ln703_615_fu_5708_p2 = (add_ln703_719_reg_12086 - data_42_V_read_3_reg_9212_pp0_iter12_reg);

assign sub_ln703_616_fu_5712_p2 = (sub_ln703_598_reg_12091 - data_42_V_read_3_reg_9212_pp0_iter12_reg);

assign sub_ln703_617_fu_5561_p2 = (sub_ln703_600_fu_5464_p2 - data_42_V_read_3_reg_9212_pp0_iter11_reg);

assign sub_ln703_618_fu_5566_p2 = (add_ln703_720_fu_5469_p2 - data_42_V_read_3_reg_9212_pp0_iter11_reg);

assign sub_ln703_619_fu_5716_p2 = (sub_ln703_602_fu_5688_p2 - data_43_V_read_3_reg_9184_pp0_iter12_reg);

assign sub_ln703_61_fu_932_p2 = (sub_ln703_44_fu_848_p2 - data_7_V_read_9_reg_10191_pp0_iter3_reg);

assign sub_ln703_620_fu_5721_p2 = (add_ln703_721_fu_5692_p2 - data_43_V_read_3_reg_9184_pp0_iter12_reg);

assign sub_ln703_621_fu_5726_p2 = (add_ln703_728_reg_12096 - data_43_V_read_3_reg_9184_pp0_iter12_reg);

assign sub_ln703_622_fu_5730_p2 = (sub_ln703_603_reg_12101 - data_43_V_read_3_reg_9184_pp0_iter12_reg);

assign sub_ln703_623_fu_5734_p2 = (sub_ln703_604_reg_12106 - data_43_V_read_3_reg_9184_pp0_iter12_reg);

assign sub_ln703_624_fu_5596_p2 = (sub_ln703_607_fu_5506_p2 - data_43_V_read_3_reg_9184_pp0_iter11_reg);

assign sub_ln703_625_fu_5742_p2 = (sub_ln703_609_reg_12121 - data_43_V_read_3_reg_9184_pp0_iter12_reg);

assign sub_ln703_626_fu_5746_p2 = (sub_ln703_610_reg_12126 - data_43_V_read_3_reg_9184_pp0_iter12_reg);

assign sub_ln703_627_fu_5750_p2 = (add_ln703_729_fu_5700_p2 - data_43_V_read_3_reg_9184_pp0_iter12_reg);

assign sub_ln703_628_fu_5755_p2 = (sub_ln703_613_reg_12136 - data_43_V_read_3_reg_9184_pp0_iter12_reg);

assign sub_ln703_629_fu_5763_p2 = (sub_ln703_615_fu_5708_p2 - data_43_V_read_3_reg_9184_pp0_iter12_reg);

assign sub_ln703_62_fu_942_p2 = (add_ln703_156_fu_872_p2 - data_7_V_read_9_reg_10191_pp0_iter3_reg);

assign sub_ln703_630_fu_5627_p2 = (add_ln703_730_fu_5541_p2 - data_43_V_read_3_reg_9184_pp0_iter11_reg);

assign sub_ln703_631_fu_5632_p2 = (add_ln703_732_fu_5546_p2 - data_43_V_read_3_reg_9184_pp0_iter11_reg);

assign sub_ln703_632_fu_5768_p2 = (add_ln703_733_reg_12146 - data_43_V_read_3_reg_9184_pp0_iter12_reg);

assign sub_ln703_633_fu_5772_p2 = (add_ln703_734_reg_12151 - data_43_V_read_3_reg_9184_pp0_iter12_reg);

assign sub_ln703_634_fu_5637_p2 = (sub_ln703_617_fu_5561_p2 - data_43_V_read_3_reg_9184_pp0_iter11_reg);

assign sub_ln703_635_fu_5780_p2 = (add_ln703_735_reg_12161 - data_43_V_read_3_reg_9184_pp0_iter12_reg);

assign sub_ln703_636_fu_5784_p2 = (sub_ln703_619_fu_5716_p2 - data_44_V_read_3_reg_9154_pp0_iter12_reg);

assign sub_ln703_637_fu_5642_p2 = (add_ln703_739_fu_5585_p2 - data_44_V_read_3_reg_9154_pp0_iter11_reg);

assign sub_ln703_638_fu_5647_p2 = (add_ln703_741_fu_5591_p2 - data_44_V_read_3_reg_9154_pp0_iter11_reg);

assign sub_ln703_639_fu_5789_p2 = (sub_ln703_620_fu_5721_p2 - data_44_V_read_3_reg_9154_pp0_iter12_reg);

assign sub_ln703_63_fu_947_p2 = (sub_ln703_48_fu_877_p2 - data_7_V_read_9_reg_10191_pp0_iter3_reg);

assign sub_ln703_640_fu_5794_p2 = (sub_ln703_622_fu_5730_p2 - data_44_V_read_3_reg_9154_pp0_iter12_reg);

assign sub_ln703_641_fu_5799_p2 = (sub_ln703_623_fu_5734_p2 - data_44_V_read_3_reg_9154_pp0_iter12_reg);

assign sub_ln703_642_fu_5804_p2 = (add_ln703_742_fu_5738_p2 - data_44_V_read_3_reg_9154_pp0_iter12_reg);

assign sub_ln703_643_fu_5822_p2 = (sub_ln703_625_fu_5742_p2 - data_44_V_read_3_reg_9154_pp0_iter12_reg);

assign sub_ln703_644_fu_5656_p2 = (add_ln703_744_fu_5601_p2 - data_44_V_read_3_reg_9154_pp0_iter11_reg);

assign sub_ln703_645_fu_5827_p2 = (sub_ln703_626_fu_5746_p2 - data_44_V_read_3_reg_9154_pp0_iter12_reg);

assign sub_ln703_646_fu_5832_p2 = (sub_ln703_627_fu_5750_p2 - data_44_V_read_3_reg_9154_pp0_iter12_reg);

assign sub_ln703_647_fu_5846_p2 = (sub_ln703_628_fu_5755_p2 - data_44_V_read_3_reg_9154_pp0_iter12_reg);

assign sub_ln703_648_fu_5661_p2 = (add_ln703_747_fu_5611_p2 - data_44_V_read_3_reg_9154_pp0_iter11_reg);

assign sub_ln703_649_fu_5851_p2 = (add_ln703_748_fu_5759_p2 - data_44_V_read_3_reg_9154_pp0_iter12_reg);

assign sub_ln703_64_fu_957_p2 = (sub_ln703_49_fu_882_p2 - data_7_V_read_9_reg_10191_pp0_iter3_reg);

assign sub_ln703_650_fu_5666_p2 = (add_ln703_753_fu_5621_p2 - data_44_V_read_3_reg_9154_pp0_iter11_reg);

assign sub_ln703_651_fu_5856_p2 = (sub_ln703_629_fu_5763_p2 - data_44_V_read_3_reg_9154_pp0_iter12_reg);

assign sub_ln703_652_fu_5865_p2 = (sub_ln703_632_fu_5768_p2 - data_44_V_read_3_reg_9154_pp0_iter12_reg);

assign sub_ln703_653_fu_5870_p2 = (sub_ln703_633_fu_5772_p2 - data_44_V_read_3_reg_9154_pp0_iter12_reg);

assign sub_ln703_654_fu_5875_p2 = (sub_ln703_634_reg_12181 - data_44_V_read_3_reg_9154_pp0_iter12_reg);

assign sub_ln703_655_fu_5879_p2 = (add_ln703_754_fu_5776_p2 - data_44_V_read_3_reg_9154_pp0_iter12_reg);

assign sub_ln703_656_fu_5884_p2 = (sub_ln703_635_fu_5780_p2 - data_44_V_read_3_reg_9154_pp0_iter12_reg);

assign sub_ln703_657_fu_5889_p2 = (sub_ln703_638_reg_12191 - data_45_V_read_3_reg_9125_pp0_iter12_reg);

assign sub_ln703_658_fu_5898_p2 = (sub_ln703_640_fu_5794_p2 - data_45_V_read_3_reg_9125_pp0_iter12_reg);

assign sub_ln703_659_fu_5903_p2 = (sub_ln703_642_fu_5804_p2 - data_45_V_read_3_reg_9125_pp0_iter12_reg);

assign sub_ln703_65_fu_1110_p2 = (add_ln703_157_reg_10529 - data_7_V_read_9_reg_10191_pp0_iter4_reg);

assign sub_ln703_660_fu_5908_p2 = (add_ln703_756_fu_5809_p2 - data_45_V_read_3_reg_9125_pp0_iter12_reg);

assign sub_ln703_661_fu_5913_p2 = (add_ln703_757_fu_5814_p2 - data_45_V_read_3_reg_9125_pp0_iter12_reg);

assign sub_ln703_662_fu_5918_p2 = (add_ln703_759_fu_5818_p2 - data_45_V_read_3_reg_9125_pp0_iter12_reg);

assign sub_ln703_663_fu_5923_p2 = (sub_ln703_643_fu_5822_p2 - data_45_V_read_3_reg_9125_pp0_iter12_reg);

assign sub_ln703_664_fu_5928_p2 = (sub_ln703_644_reg_12204 - data_45_V_read_3_reg_9125_pp0_iter12_reg);

assign sub_ln703_665_fu_5932_p2 = (sub_ln703_646_fu_5832_p2 - data_45_V_read_3_reg_9125_pp0_iter12_reg);

assign sub_ln703_666_fu_5937_p2 = (add_ln703_761_fu_5837_p2 - data_45_V_read_3_reg_9125_pp0_iter12_reg);

assign sub_ln703_667_fu_5956_p2 = (add_ln703_763_fu_5842_p2 - data_45_V_read_3_reg_9125_pp0_iter12_reg);

assign sub_ln703_668_fu_5971_p2 = (sub_ln703_650_reg_12214 - data_45_V_read_3_reg_9125_pp0_iter12_reg);

assign sub_ln703_669_fu_5975_p2 = (sub_ln703_651_fu_5856_p2 - data_45_V_read_3_reg_9125_pp0_iter12_reg);

assign sub_ln703_66_fu_987_p2 = (add_ln703_160_fu_902_p2 - data_7_V_read_9_reg_10191_pp0_iter3_reg);

assign sub_ln703_670_fu_5980_p2 = (add_ln703_764_fu_5861_p2 - data_45_V_read_3_reg_9125_pp0_iter12_reg);

assign sub_ln703_671_fu_5989_p2 = (sub_ln703_652_fu_5865_p2 - data_45_V_read_3_reg_9125_pp0_iter12_reg);

assign sub_ln703_672_fu_6004_p2 = (sub_ln703_653_fu_5870_p2 - data_45_V_read_3_reg_9125_pp0_iter12_reg);

assign sub_ln703_673_fu_6009_p2 = (sub_ln703_654_fu_5875_p2 - data_45_V_read_3_reg_9125_pp0_iter12_reg);

assign sub_ln703_674_fu_6014_p2 = (sub_ln703_655_fu_5879_p2 - data_45_V_read_3_reg_9125_pp0_iter12_reg);

assign sub_ln703_675_fu_6019_p2 = (sub_ln703_656_fu_5884_p2 - data_45_V_read_3_reg_9125_pp0_iter12_reg);

assign sub_ln703_676_fu_6033_p2 = (sub_ln703_657_fu_5889_p2 - data_46_V_read_3_reg_9094_pp0_iter12_reg);

assign sub_ln703_677_fu_6047_p2 = (add_ln703_766_fu_5893_p2 - data_46_V_read_3_reg_9094_pp0_iter12_reg);

assign sub_ln703_678_fu_6052_p2 = (sub_ln703_658_fu_5898_p2 - data_46_V_read_3_reg_9094_pp0_iter12_reg);

assign sub_ln703_679_fu_6057_p2 = (sub_ln703_659_fu_5903_p2 - data_46_V_read_3_reg_9094_pp0_iter12_reg);

assign sub_ln703_67_fu_1119_p2 = (add_ln703_162_reg_10539 - data_8_V_read_8_reg_10164_pp0_iter4_reg);

assign sub_ln703_680_fu_6062_p2 = (sub_ln703_660_fu_5908_p2 - data_46_V_read_3_reg_9094_pp0_iter12_reg);

assign sub_ln703_681_fu_6238_p2 = (sub_ln703_662_reg_12248 - data_46_V_read_3_reg_9094_pp0_iter13_reg);

assign sub_ln703_682_fu_6067_p2 = (sub_ln703_664_fu_5928_p2 - data_46_V_read_3_reg_9094_pp0_iter12_reg);

assign sub_ln703_683_fu_6242_p2 = (sub_ln703_665_reg_12253 - data_46_V_read_3_reg_9094_pp0_iter13_reg);

assign sub_ln703_684_fu_6072_p2 = (sub_ln703_666_fu_5937_p2 - data_46_V_read_3_reg_9094_pp0_iter12_reg);

assign sub_ln703_685_fu_6246_p2 = (add_ln703_770_reg_12258 - data_46_V_read_3_reg_9094_pp0_iter13_reg);

assign sub_ln703_686_fu_6077_p2 = (add_ln703_771_fu_5961_p2 - data_46_V_read_3_reg_9094_pp0_iter12_reg);

assign sub_ln703_687_fu_6086_p2 = (add_ln703_772_fu_5966_p2 - data_46_V_read_3_reg_9094_pp0_iter12_reg);

assign sub_ln703_688_fu_6091_p2 = (sub_ln703_668_fu_5971_p2 - data_46_V_read_3_reg_9094_pp0_iter12_reg);

assign sub_ln703_689_fu_6096_p2 = (sub_ln703_670_fu_5980_p2 - data_46_V_read_3_reg_9094_pp0_iter12_reg);

assign sub_ln703_68_fu_1133_p2 = (add_ln703_163_fu_1098_p2 - data_8_V_read_8_reg_10164_pp0_iter4_reg);

assign sub_ln703_690_fu_6101_p2 = (add_ln703_774_fu_5985_p2 - data_46_V_read_3_reg_9094_pp0_iter12_reg);

assign sub_ln703_691_fu_6106_p2 = (sub_ln703_671_fu_5989_p2 - data_46_V_read_3_reg_9094_pp0_iter12_reg);

assign sub_ln703_692_fu_6111_p2 = (add_ln703_777_fu_5999_p2 - data_46_V_read_3_reg_9094_pp0_iter12_reg);

assign sub_ln703_693_fu_6116_p2 = (sub_ln703_672_fu_6004_p2 - data_46_V_read_3_reg_9094_pp0_iter12_reg);

assign sub_ln703_694_fu_6126_p2 = (sub_ln703_674_fu_6014_p2 - data_46_V_read_3_reg_9094_pp0_iter12_reg);

assign sub_ln703_695_fu_6254_p2 = (add_ln703_779_reg_12273 - data_47_V_read_3_reg_9066_pp0_iter13_reg);

assign sub_ln703_696_fu_6136_p2 = (add_ln703_781_fu_6029_p2 - data_47_V_read_3_reg_9066_pp0_iter12_reg);

assign sub_ln703_697_fu_6141_p2 = (add_ln703_786_fu_6042_p2 - data_47_V_read_3_reg_9066_pp0_iter12_reg);

assign sub_ln703_698_fu_6267_p2 = (sub_ln703_682_reg_12298 - data_47_V_read_3_reg_9066_pp0_iter13_reg);

assign sub_ln703_699_fu_6271_p2 = (sub_ln703_683_fu_6242_p2 - data_47_V_read_3_reg_9066_pp0_iter13_reg);

assign sub_ln703_69_fu_1138_p2 = (sub_ln703_57_fu_1102_p2 - data_8_V_read_8_reg_10164_pp0_iter4_reg);

assign sub_ln703_6_fu_595_p2 = (sub_ln703_2_reg_10367 - data_3_V_read_10_reg_10295_pp0_iter2_reg);

assign sub_ln703_700_fu_6172_p2 = (add_ln703_788_fu_6082_p2 - data_47_V_read_3_reg_9066_pp0_iter12_reg);

assign sub_ln703_701_fu_6281_p2 = (sub_ln703_687_reg_12313 - data_47_V_read_3_reg_9066_pp0_iter13_reg);

assign sub_ln703_702_fu_6285_p2 = (sub_ln703_688_reg_12318 - data_47_V_read_3_reg_9066_pp0_iter13_reg);

assign sub_ln703_703_fu_6289_p2 = (add_ln703_789_fu_6250_p2 - data_47_V_read_3_reg_9066_pp0_iter13_reg);

assign sub_ln703_704_fu_6177_p2 = (sub_ln703_689_fu_6096_p2 - data_47_V_read_3_reg_9066_pp0_iter12_reg);

assign sub_ln703_705_fu_6294_p2 = (sub_ln703_691_reg_12328 - data_47_V_read_3_reg_9066_pp0_iter13_reg);

assign sub_ln703_706_fu_6298_p2 = (sub_ln703_693_reg_12338 - data_47_V_read_3_reg_9066_pp0_iter13_reg);

assign sub_ln703_707_fu_6182_p2 = (add_ln703_790_fu_6121_p2 - data_47_V_read_3_reg_9066_pp0_iter12_reg);

assign sub_ln703_708_fu_6302_p2 = (add_ln703_791_reg_12348 - data_47_V_read_3_reg_9066_pp0_iter13_reg);

assign sub_ln703_709_fu_6306_p2 = (sub_ln703_695_fu_6254_p2 - data_48_V_read_3_reg_9040_pp0_iter13_reg);

assign sub_ln703_70_fu_992_p2 = (sub_ln703_60_fu_927_p2 - data_8_V_read_8_reg_10164_pp0_iter3_reg);

assign sub_ln703_710_fu_6311_p2 = (sub_ln703_696_reg_12353 - data_48_V_read_3_reg_9040_pp0_iter13_reg);

assign sub_ln703_711_fu_6328_p2 = (add_ln703_792_reg_12363 - data_48_V_read_3_reg_9040_pp0_iter13_reg);

assign sub_ln703_712_fu_6332_p2 = (add_ln703_793_fu_6258_p2 - data_48_V_read_3_reg_9040_pp0_iter13_reg);

assign sub_ln703_713_fu_6337_p2 = (add_ln703_796_reg_12368 - data_48_V_read_3_reg_9040_pp0_iter13_reg);

assign sub_ln703_714_fu_6345_p2 = (add_ln703_797_fu_6262_p2 - data_48_V_read_3_reg_9040_pp0_iter13_reg);

assign sub_ln703_715_fu_6350_p2 = (add_ln703_798_reg_12373 - data_48_V_read_3_reg_9040_pp0_iter13_reg);

assign sub_ln703_716_fu_6354_p2 = (sub_ln703_698_fu_6267_p2 - data_48_V_read_3_reg_9040_pp0_iter13_reg);

assign sub_ln703_717_fu_6364_p2 = (add_ln703_799_fu_6276_p2 - data_48_V_read_3_reg_9040_pp0_iter13_reg);

assign sub_ln703_718_fu_6382_p2 = (sub_ln703_700_reg_12378 - data_48_V_read_3_reg_9040_pp0_iter13_reg);

assign sub_ln703_719_fu_6386_p2 = (sub_ln703_701_fu_6281_p2 - data_48_V_read_3_reg_9040_pp0_iter13_reg);

assign sub_ln703_71_fu_1002_p2 = (add_ln703_164_fu_937_p2 - data_8_V_read_8_reg_10164_pp0_iter3_reg);

assign sub_ln703_720_fu_6391_p2 = (sub_ln703_702_fu_6285_p2 - data_48_V_read_3_reg_9040_pp0_iter13_reg);

assign sub_ln703_721_fu_6413_p2 = (sub_ln703_707_reg_12388 - data_48_V_read_3_reg_9040_pp0_iter13_reg);

assign sub_ln703_722_fu_6422_p2 = (sub_ln703_709_fu_6306_p2 - data_49_V_read_3_reg_9012_pp0_iter13_reg);

assign sub_ln703_723_fu_6427_p2 = (add_ln703_800_fu_6315_p2 - data_49_V_read_3_reg_9012_pp0_iter13_reg);

assign sub_ln703_724_fu_6432_p2 = (add_ln703_804_fu_6323_p2 - data_49_V_read_3_reg_9012_pp0_iter13_reg);

assign sub_ln703_725_fu_6437_p2 = (sub_ln703_713_fu_6337_p2 - data_49_V_read_3_reg_9012_pp0_iter13_reg);

assign sub_ln703_726_fu_6442_p2 = (add_ln703_805_fu_6341_p2 - data_49_V_read_3_reg_9012_pp0_iter13_reg);

assign sub_ln703_727_fu_6452_p2 = (sub_ln703_715_fu_6350_p2 - data_49_V_read_3_reg_9012_pp0_iter13_reg);

assign sub_ln703_728_fu_6457_p2 = (add_ln703_806_fu_6359_p2 - data_49_V_read_3_reg_9012_pp0_iter13_reg);

assign sub_ln703_729_fu_6462_p2 = (add_ln703_808_fu_6373_p2 - data_49_V_read_3_reg_9012_pp0_iter13_reg);

assign sub_ln703_72_fu_1147_p2 = (sub_ln703_63_reg_10555 - data_8_V_read_8_reg_10164_pp0_iter4_reg);

assign sub_ln703_730_fu_6467_p2 = (add_ln703_809_fu_6378_p2 - data_49_V_read_3_reg_9012_pp0_iter13_reg);

assign sub_ln703_731_fu_6472_p2 = (sub_ln703_718_fu_6382_p2 - data_49_V_read_3_reg_9012_pp0_iter13_reg);

assign sub_ln703_732_fu_6477_p2 = (sub_ln703_719_fu_6386_p2 - data_49_V_read_3_reg_9012_pp0_iter13_reg);

assign sub_ln703_733_fu_6487_p2 = (add_ln703_810_fu_6396_p2 - data_49_V_read_3_reg_9012_pp0_iter13_reg);

assign sub_ln703_734_fu_6492_p2 = (add_ln703_811_fu_6401_p2 - data_49_V_read_3_reg_9012_pp0_iter13_reg);

assign sub_ln703_735_fu_6497_p2 = (add_ln703_812_fu_6405_p2 - data_49_V_read_3_reg_9012_pp0_iter13_reg);

assign sub_ln703_736_fu_6502_p2 = (add_ln703_813_fu_6409_p2 - data_49_V_read_3_reg_9012_pp0_iter13_reg);

assign sub_ln703_737_fu_6507_p2 = (sub_ln703_721_fu_6413_p2 - data_49_V_read_3_reg_9012_pp0_iter13_reg);

assign sub_ln703_738_fu_6521_p2 = (add_ln703_814_fu_6417_p2 - data_49_V_read_3_reg_9012_pp0_iter13_reg);

assign sub_ln703_739_fu_6541_p2 = (sub_ln703_725_fu_6437_p2 - data_50_V_read51_reg_8984_pp0_iter13_reg);

assign sub_ln703_73_fu_1026_p2 = (add_ln703_165_fu_952_p2 - data_8_V_read_8_reg_10164_pp0_iter3_reg);

assign sub_ln703_740_fu_6560_p2 = (sub_ln703_726_fu_6442_p2 - data_50_V_read51_reg_8984_pp0_iter13_reg);

assign sub_ln703_741_fu_6795_p2 = (add_ln703_818_reg_12409_pp0_iter14_reg - data_50_V_read51_reg_8984_pp0_iter14_reg);

assign sub_ln703_742_fu_6799_p2 = (add_ln703_819_reg_12455 - data_50_V_read51_reg_8984_pp0_iter14_reg);

assign sub_ln703_743_fu_6803_p2 = (sub_ln703_727_reg_12460 - data_50_V_read51_reg_8984_pp0_iter14_reg);

assign sub_ln703_744_fu_6565_p2 = (add_ln703_821_reg_12414 - data_50_V_read51_reg_8984_pp0_iter13_reg);

assign sub_ln703_745_fu_6807_p2 = (sub_ln703_728_reg_12465 - data_50_V_read51_reg_8984_pp0_iter14_reg);

assign sub_ln703_746_fu_6579_p2 = (sub_ln703_729_fu_6462_p2 - data_50_V_read51_reg_8984_pp0_iter13_reg);

assign sub_ln703_747_fu_6584_p2 = (sub_ln703_730_fu_6467_p2 - data_50_V_read51_reg_8984_pp0_iter13_reg);

assign sub_ln703_748_fu_6589_p2 = (sub_ln703_731_fu_6472_p2 - data_50_V_read51_reg_8984_pp0_iter13_reg);

assign sub_ln703_749_fu_6599_p2 = (add_ln703_822_fu_6482_p2 - data_50_V_read51_reg_8984_pp0_iter13_reg);

assign sub_ln703_74_fu_1151_p2 = (sub_ln703_64_reg_10560 - data_8_V_read_8_reg_10164_pp0_iter4_reg);

assign sub_ln703_750_fu_6811_p2 = (sub_ln703_733_reg_12470 - data_50_V_read51_reg_8984_pp0_iter14_reg);

assign sub_ln703_751_fu_6604_p2 = (sub_ln703_734_fu_6492_p2 - data_50_V_read51_reg_8984_pp0_iter13_reg);

assign sub_ln703_752_fu_6609_p2 = (sub_ln703_735_fu_6497_p2 - data_50_V_read51_reg_8984_pp0_iter13_reg);

assign sub_ln703_753_fu_6614_p2 = (sub_ln703_737_fu_6507_p2 - data_50_V_read51_reg_8984_pp0_iter13_reg);

assign sub_ln703_754_fu_6619_p2 = (add_ln703_824_fu_6516_p2 - data_50_V_read51_reg_8984_pp0_iter13_reg);

assign sub_ln703_755_fu_6819_p2 = (add_ln703_825_reg_12480 - data_51_V_read52_reg_8956_pp0_iter14_reg);

assign sub_ln703_756_fu_6823_p2 = (add_ln703_827_reg_12485 - data_51_V_read52_reg_8956_pp0_iter14_reg);

assign sub_ln703_757_fu_6629_p2 = (add_ln703_828_fu_6536_p2 - data_51_V_read52_reg_8956_pp0_iter13_reg);

assign sub_ln703_758_fu_6827_p2 = (add_ln703_831_reg_12490 - data_51_V_read52_reg_8956_pp0_iter14_reg);

assign sub_ln703_759_fu_6639_p2 = (sub_ln703_740_fu_6560_p2 - data_51_V_read52_reg_8956_pp0_iter13_reg);

assign sub_ln703_75_fu_1031_p2 = (add_ln703_168_fu_967_p2 - data_8_V_read_8_reg_10164_pp0_iter3_reg);

assign sub_ln703_760_fu_6831_p2 = (sub_ln703_741_fu_6795_p2 - data_51_V_read52_reg_8956_pp0_iter14_reg);

assign sub_ln703_761_fu_6644_p2 = (sub_ln703_744_fu_6565_p2 - data_51_V_read52_reg_8956_pp0_iter13_reg);

assign sub_ln703_762_fu_6841_p2 = (add_ln703_833_reg_12495 - data_51_V_read52_reg_8956_pp0_iter14_reg);

assign sub_ln703_763_fu_6654_p2 = (sub_ln703_748_fu_6589_p2 - data_51_V_read52_reg_8956_pp0_iter13_reg);

assign sub_ln703_764_fu_6845_p2 = (add_ln703_834_reg_12505 - data_51_V_read52_reg_8956_pp0_iter14_reg);

assign sub_ln703_765_fu_6849_p2 = (sub_ln703_749_reg_12510 - data_51_V_read52_reg_8956_pp0_iter14_reg);

assign sub_ln703_766_fu_6853_p2 = (sub_ln703_750_fu_6811_p2 - data_51_V_read52_reg_8956_pp0_iter14_reg);

assign sub_ln703_767_fu_6659_p2 = (sub_ln703_751_fu_6604_p2 - data_51_V_read52_reg_8956_pp0_iter13_reg);

assign sub_ln703_768_fu_6858_p2 = (add_ln703_835_fu_6815_p2 - data_51_V_read52_reg_8956_pp0_iter14_reg);

assign sub_ln703_769_fu_6684_p2 = (sub_ln703_753_fu_6614_p2 - data_51_V_read52_reg_8956_pp0_iter13_reg);

assign sub_ln703_76_fu_1155_p2 = (add_ln703_170_reg_10566 - data_8_V_read_8_reg_10164_pp0_iter4_reg);

assign sub_ln703_770_fu_6708_p2 = (add_ln703_837_fu_6624_p2 - data_52_V_read_3_reg_8928_pp0_iter13_reg);

assign sub_ln703_771_fu_6873_p2 = (add_ln703_838_reg_12520 - data_52_V_read_3_reg_8928_pp0_iter14_reg);

assign sub_ln703_772_fu_6877_p2 = (sub_ln703_758_fu_6827_p2 - data_52_V_read_3_reg_8928_pp0_iter14_reg);

assign sub_ln703_773_fu_6886_p2 = (sub_ln703_760_fu_6831_p2 - data_52_V_read_3_reg_8928_pp0_iter14_reg);

assign sub_ln703_774_fu_6896_p2 = (add_ln703_839_fu_6836_p2 - data_52_V_read_3_reg_8928_pp0_iter14_reg);

assign sub_ln703_775_fu_6910_p2 = (sub_ln703_762_fu_6841_p2 - data_52_V_read_3_reg_8928_pp0_iter14_reg);

assign sub_ln703_776_fu_6915_p2 = (add_ln703_840_reg_12535 - data_52_V_read_3_reg_8928_pp0_iter14_reg);

assign sub_ln703_777_fu_6928_p2 = (sub_ln703_765_fu_6849_p2 - data_52_V_read_3_reg_8928_pp0_iter14_reg);

assign sub_ln703_778_fu_6933_p2 = (sub_ln703_766_fu_6853_p2 - data_52_V_read_3_reg_8928_pp0_iter14_reg);

assign sub_ln703_779_fu_6938_p2 = (sub_ln703_767_reg_12545 - data_52_V_read_3_reg_8928_pp0_iter14_reg);

assign sub_ln703_77_fu_1159_p2 = (sub_ln703_65_fu_1110_p2 - data_8_V_read_8_reg_10164_pp0_iter4_reg);

assign sub_ln703_780_fu_6942_p2 = (add_ln703_841_reg_12550 - data_52_V_read_3_reg_8928_pp0_iter14_reg);

assign sub_ln703_781_fu_6739_p2 = (add_ln703_844_fu_6678_p2 - data_52_V_read_3_reg_8928_pp0_iter13_reg);

assign sub_ln703_782_fu_6946_p2 = (sub_ln703_769_reg_12555 - data_52_V_read_3_reg_8928_pp0_iter14_reg);

assign sub_ln703_783_fu_6950_p2 = (add_ln703_845_reg_12560 - data_52_V_read_3_reg_8928_pp0_iter14_reg);

assign sub_ln703_784_fu_6954_p2 = (add_ln703_846_fu_6863_p2 - data_53_V_read_3_reg_8899_pp0_iter14_reg);

assign sub_ln703_785_fu_6959_p2 = (add_ln703_847_fu_6868_p2 - data_53_V_read_3_reg_8899_pp0_iter14_reg);

assign sub_ln703_786_fu_6964_p2 = (add_ln703_851_reg_12565 - data_53_V_read_3_reg_8899_pp0_iter14_reg);

assign sub_ln703_787_fu_6759_p2 = (add_ln703_854_fu_6722_p2 - data_53_V_read_3_reg_8899_pp0_iter13_reg);

assign sub_ln703_788_fu_6981_p2 = (sub_ln703_772_fu_6877_p2 - data_53_V_read_3_reg_8899_pp0_iter14_reg);

assign sub_ln703_789_fu_6986_p2 = (add_ln703_855_fu_6882_p2 - data_53_V_read_3_reg_8899_pp0_iter14_reg);

assign sub_ln703_78_fu_1164_p2 = (add_ln703_171_reg_10571 - data_8_V_read_8_reg_10164_pp0_iter4_reg);

assign sub_ln703_790_fu_6991_p2 = (add_ln703_856_fu_6891_p2 - data_53_V_read_3_reg_8899_pp0_iter14_reg);

assign sub_ln703_791_fu_6996_p2 = (add_ln703_858_reg_12575 - data_53_V_read_3_reg_8899_pp0_iter14_reg);

assign sub_ln703_792_fu_7000_p2 = (add_ln703_859_fu_6901_p2 - data_53_V_read_3_reg_8899_pp0_iter14_reg);

assign sub_ln703_793_fu_7005_p2 = (add_ln703_860_fu_6905_p2 - data_53_V_read_3_reg_8899_pp0_iter14_reg);

assign sub_ln703_794_fu_7010_p2 = (sub_ln703_775_fu_6910_p2 - data_53_V_read_3_reg_8899_pp0_iter14_reg);

assign sub_ln703_795_fu_7015_p2 = (add_ln703_861_fu_6919_p2 - data_53_V_read_3_reg_8899_pp0_iter14_reg);

assign sub_ln703_796_fu_7020_p2 = (add_ln703_862_fu_6923_p2 - data_53_V_read_3_reg_8899_pp0_iter14_reg);

assign sub_ln703_797_fu_7030_p2 = (sub_ln703_778_fu_6933_p2 - data_53_V_read_3_reg_8899_pp0_iter14_reg);

assign sub_ln703_798_fu_7035_p2 = (sub_ln703_779_fu_6938_p2 - data_53_V_read_3_reg_8899_pp0_iter14_reg);

assign sub_ln703_799_fu_6764_p2 = (add_ln703_864_fu_6749_p2 - data_53_V_read_3_reg_8899_pp0_iter13_reg);

assign sub_ln703_79_fu_1168_p2 = (add_ln703_173_reg_10576 - data_8_V_read_8_reg_10164_pp0_iter4_reg);

assign sub_ln703_7_fu_607_p2 = (add_ln703_130_reg_10373 - data_3_V_read_10_reg_10295_pp0_iter2_reg);

assign sub_ln703_800_fu_7045_p2 = (sub_ln703_783_fu_6950_p2 - data_53_V_read_3_reg_8899_pp0_iter14_reg);

assign sub_ln703_801_fu_7060_p2 = (sub_ln703_786_fu_6964_p2 - data_54_V_read_3_reg_8873_pp0_iter14_reg);

assign sub_ln703_802_fu_7065_p2 = (add_ln703_865_fu_6968_p2 - data_54_V_read_3_reg_8873_pp0_iter14_reg);

assign sub_ln703_803_fu_7070_p2 = (add_ln703_869_fu_6976_p2 - data_54_V_read_3_reg_8873_pp0_iter14_reg);

assign sub_ln703_804_fu_7075_p2 = (sub_ln703_787_reg_12590 - data_54_V_read_3_reg_8873_pp0_iter14_reg);

assign sub_ln703_805_fu_7079_p2 = (sub_ln703_790_fu_6991_p2 - data_54_V_read_3_reg_8873_pp0_iter14_reg);

assign sub_ln703_806_fu_7089_p2 = (sub_ln703_792_fu_7000_p2 - data_54_V_read_3_reg_8873_pp0_iter14_reg);

assign sub_ln703_807_fu_7099_p2 = (sub_ln703_794_fu_7010_p2 - data_54_V_read_3_reg_8873_pp0_iter14_reg);

assign sub_ln703_808_fu_7137_p2 = (add_ln703_870_fu_7025_p2 - data_54_V_read_3_reg_8873_pp0_iter14_reg);

assign sub_ln703_809_fu_7165_p2 = (add_ln703_871_fu_7040_p2 - data_54_V_read_3_reg_8873_pp0_iter14_reg);

assign sub_ln703_80_fu_1184_p2 = (add_ln703_174_fu_1114_p2 - data_9_V_read_8_reg_10136_pp0_iter4_reg);

assign sub_ln703_810_fu_7170_p2 = (sub_ln703_800_fu_7045_p2 - data_54_V_read_3_reg_8873_pp0_iter14_reg);

assign sub_ln703_811_fu_7346_p2 = (add_ln703_872_reg_12650 - data_55_V_read_3_reg_8844_pp0_iter15_reg);

assign sub_ln703_812_fu_7350_p2 = (add_ln703_873_reg_12655 - data_55_V_read_3_reg_8844_pp0_iter15_reg);

assign sub_ln703_813_fu_7370_p2 = (add_ln703_874_reg_12675 - data_55_V_read_3_reg_8844_pp0_iter15_reg);

assign sub_ln703_814_fu_7200_p2 = (sub_ln703_806_fu_7089_p2 - data_55_V_read_3_reg_8844_pp0_iter14_reg);

assign sub_ln703_815_fu_7374_p2 = (add_ln703_875_reg_12680 - data_55_V_read_3_reg_8844_pp0_iter15_reg);

assign sub_ln703_816_fu_7205_p2 = (add_ln703_879_fu_7108_p2 - data_55_V_read_3_reg_8844_pp0_iter14_reg);

assign sub_ln703_817_fu_7382_p2 = (add_ln703_882_reg_12690 - data_55_V_read_3_reg_8844_pp0_iter15_reg);

assign sub_ln703_818_fu_7210_p2 = (add_ln703_883_fu_7127_p2 - data_55_V_read_3_reg_8844_pp0_iter14_reg);

assign sub_ln703_819_fu_7386_p2 = (add_ln703_884_reg_12695 - data_55_V_read_3_reg_8844_pp0_iter15_reg);

assign sub_ln703_81_fu_1194_p2 = (add_ln703_175_fu_1123_p2 - data_9_V_read_8_reg_10136_pp0_iter4_reg);

assign sub_ln703_820_fu_7215_p2 = (add_ln703_885_fu_7142_p2 - data_55_V_read_3_reg_8844_pp0_iter14_reg);

assign sub_ln703_821_fu_7220_p2 = (add_ln703_886_fu_7147_p2 - data_55_V_read_3_reg_8844_pp0_iter14_reg);

assign sub_ln703_822_fu_7398_p2 = (add_ln703_888_reg_12705 - data_55_V_read_3_reg_8844_pp0_iter15_reg);

assign sub_ln703_823_fu_7225_p2 = (add_ln703_889_fu_7161_p2 - data_55_V_read_3_reg_8844_pp0_iter14_reg);

assign sub_ln703_824_fu_7230_p2 = (sub_ln703_809_fu_7165_p2 - data_55_V_read_3_reg_8844_pp0_iter14_reg);

assign sub_ln703_825_fu_7235_p2 = (sub_ln703_810_fu_7170_p2 - data_55_V_read_3_reg_8844_pp0_iter14_reg);

assign sub_ln703_826_fu_7407_p2 = (sub_ln703_812_fu_7350_p2 - data_56_V_read_3_reg_8814_pp0_iter15_reg);

assign sub_ln703_827_fu_7412_p2 = (add_ln703_890_fu_7354_p2 - data_56_V_read_3_reg_8814_pp0_iter15_reg);

assign sub_ln703_828_fu_7417_p2 = (add_ln703_891_fu_7358_p2 - data_56_V_read_3_reg_8814_pp0_iter15_reg);

assign sub_ln703_829_fu_7422_p2 = (add_ln703_892_reg_12710 - data_56_V_read_3_reg_8814_pp0_iter15_reg);

assign sub_ln703_82_fu_1199_p2 = (add_ln703_176_fu_1128_p2 - data_9_V_read_8_reg_10136_pp0_iter4_reg);

assign sub_ln703_830_fu_7426_p2 = (add_ln703_893_reg_12715 - data_56_V_read_3_reg_8814_pp0_iter15_reg);

assign sub_ln703_831_fu_7430_p2 = (add_ln703_895_reg_12720 - data_56_V_read_3_reg_8814_pp0_iter15_reg);

assign sub_ln703_832_fu_7434_p2 = (add_ln703_897_fu_7362_p2 - data_56_V_read_3_reg_8814_pp0_iter15_reg);

assign sub_ln703_833_fu_7439_p2 = (add_ln703_899_fu_7366_p2 - data_56_V_read_3_reg_8814_pp0_iter15_reg);

assign sub_ln703_834_fu_7444_p2 = (sub_ln703_813_fu_7370_p2 - data_56_V_read_3_reg_8814_pp0_iter15_reg);

assign sub_ln703_835_fu_7449_p2 = (sub_ln703_814_reg_12735 - data_56_V_read_3_reg_8814_pp0_iter15_reg);

assign sub_ln703_836_fu_7453_p2 = (sub_ln703_815_fu_7374_p2 - data_56_V_read_3_reg_8814_pp0_iter15_reg);

assign sub_ln703_837_fu_7458_p2 = (add_ln703_900_fu_7378_p2 - data_56_V_read_3_reg_8814_pp0_iter15_reg);

assign sub_ln703_838_fu_7463_p2 = (sub_ln703_818_reg_12745 - data_56_V_read_3_reg_8814_pp0_iter15_reg);

assign sub_ln703_839_fu_7467_p2 = (add_ln703_901_fu_7390_p2 - data_56_V_read_3_reg_8814_pp0_iter15_reg);

assign sub_ln703_83_fu_1218_p2 = (sub_ln703_70_reg_10586 - data_9_V_read_8_reg_10136_pp0_iter4_reg);

assign sub_ln703_840_fu_7472_p2 = (add_ln703_902_fu_7394_p2 - data_56_V_read_3_reg_8814_pp0_iter15_reg);

assign sub_ln703_841_fu_7485_p2 = (sub_ln703_822_fu_7398_p2 - data_56_V_read_3_reg_8814_pp0_iter15_reg);

assign sub_ln703_842_fu_7498_p2 = (add_ln703_903_fu_7402_p2 - data_57_V_read_3_reg_8786_pp0_iter15_reg);

assign sub_ln703_843_fu_7503_p2 = (sub_ln703_826_fu_7407_p2 - data_57_V_read_3_reg_8786_pp0_iter15_reg);

assign sub_ln703_844_fu_7508_p2 = (sub_ln703_827_fu_7412_p2 - data_57_V_read_3_reg_8786_pp0_iter15_reg);

assign sub_ln703_845_fu_7518_p2 = (sub_ln703_829_fu_7422_p2 - data_57_V_read_3_reg_8786_pp0_iter15_reg);

assign sub_ln703_846_fu_7523_p2 = (sub_ln703_831_fu_7430_p2 - data_57_V_read_3_reg_8786_pp0_iter15_reg);

assign sub_ln703_847_fu_7528_p2 = (add_ln703_906_reg_12775 - data_57_V_read_3_reg_8786_pp0_iter15_reg);

assign sub_ln703_848_fu_7551_p2 = (sub_ln703_834_fu_7444_p2 - data_57_V_read_3_reg_8786_pp0_iter15_reg);

assign sub_ln703_849_fu_7556_p2 = (sub_ln703_836_fu_7453_p2 - data_57_V_read_3_reg_8786_pp0_iter15_reg);

assign sub_ln703_84_fu_1222_p2 = (add_ln703_177_reg_10591 - data_9_V_read_8_reg_10136_pp0_iter4_reg);

assign sub_ln703_850_fu_7566_p2 = (sub_ln703_839_fu_7467_p2 - data_57_V_read_3_reg_8786_pp0_iter15_reg);

assign sub_ln703_851_fu_7571_p2 = (add_ln703_907_fu_7477_p2 - data_57_V_read_3_reg_8786_pp0_iter15_reg);

assign sub_ln703_852_fu_7319_p2 = (add_ln703_910_fu_7259_p2 - data_57_V_read_3_reg_8786_pp0_iter14_reg);

assign sub_ln703_853_fu_7576_p2 = (add_ln703_911_fu_7481_p2 - data_57_V_read_3_reg_8786_pp0_iter15_reg);

assign sub_ln703_854_fu_7586_p2 = (add_ln703_912_fu_7490_p2 - data_57_V_read_3_reg_8786_pp0_iter15_reg);

assign sub_ln703_855_fu_7591_p2 = (add_ln703_913_fu_7494_p2 - data_57_V_read_3_reg_8786_pp0_iter15_reg);

assign sub_ln703_856_fu_7596_p2 = (add_ln703_917_reg_12780 - data_57_V_read_3_reg_8786_pp0_iter15_reg);

assign sub_ln703_857_fu_7600_p2 = (sub_ln703_842_fu_7498_p2 - data_58_V_read_3_reg_8756_pp0_iter15_reg);

assign sub_ln703_858_fu_7605_p2 = (sub_ln703_843_fu_7503_p2 - data_58_V_read_3_reg_8756_pp0_iter15_reg);

assign sub_ln703_859_fu_7615_p2 = (add_ln703_918_fu_7513_p2 - data_58_V_read_3_reg_8756_pp0_iter15_reg);

assign sub_ln703_85_fu_1230_p2 = (add_ln703_181_reg_10601 - data_9_V_read_8_reg_10136_pp0_iter4_reg);

assign sub_ln703_860_fu_7620_p2 = (sub_ln703_845_fu_7518_p2 - data_58_V_read_3_reg_8756_pp0_iter15_reg);

assign sub_ln703_861_fu_7625_p2 = (add_ln703_922_reg_12785 - data_58_V_read_3_reg_8756_pp0_iter15_reg);

assign sub_ln703_862_fu_7324_p2 = (add_ln703_925_fu_7302_p2 - data_58_V_read_3_reg_8756_pp0_iter14_reg);

assign sub_ln703_863_fu_7639_p2 = (add_ln703_926_fu_7532_p2 - data_58_V_read_3_reg_8756_pp0_iter15_reg);

assign sub_ln703_864_fu_7644_p2 = (add_ln703_928_fu_7541_p2 - data_58_V_read_3_reg_8756_pp0_iter15_reg);

assign sub_ln703_865_fu_7649_p2 = (add_ln703_929_fu_7546_p2 - data_58_V_read_3_reg_8756_pp0_iter15_reg);

assign sub_ln703_866_fu_7654_p2 = (sub_ln703_848_fu_7551_p2 - data_58_V_read_3_reg_8756_pp0_iter15_reg);

assign sub_ln703_867_fu_7669_p2 = (sub_ln703_849_fu_7556_p2 - data_58_V_read_3_reg_8756_pp0_iter15_reg);

assign sub_ln703_868_fu_7674_p2 = (add_ln703_930_fu_7561_p2 - data_58_V_read_3_reg_8756_pp0_iter15_reg);

assign sub_ln703_869_fu_7329_p2 = (add_ln703_932_fu_7313_p2 - data_58_V_read_3_reg_8756_pp0_iter14_reg);

assign sub_ln703_86_fu_1234_p2 = (add_ln703_183_reg_10606 - data_9_V_read_8_reg_10136_pp0_iter4_reg);

assign sub_ln703_870_fu_7685_p2 = (sub_ln703_850_fu_7566_p2 - data_58_V_read_3_reg_8756_pp0_iter15_reg);

assign sub_ln703_871_fu_7696_p2 = (sub_ln703_851_fu_7571_p2 - data_58_V_read_3_reg_8756_pp0_iter15_reg);

assign sub_ln703_872_fu_7705_p2 = (sub_ln703_853_fu_7576_p2 - data_58_V_read_3_reg_8756_pp0_iter15_reg);

assign sub_ln703_873_fu_7710_p2 = (add_ln703_933_fu_7581_p2 - data_58_V_read_3_reg_8756_pp0_iter15_reg);

assign sub_ln703_874_fu_7725_p2 = (sub_ln703_855_fu_7591_p2 - data_58_V_read_3_reg_8756_pp0_iter15_reg);

assign sub_ln703_875_fu_7730_p2 = (sub_ln703_856_fu_7596_p2 - data_58_V_read_3_reg_8756_pp0_iter15_reg);

assign sub_ln703_876_fu_7878_p2 = (sub_ln703_857_reg_12835 - data_59_V_read_3_reg_8724_pp0_iter16_reg);

assign sub_ln703_877_fu_7886_p2 = (add_ln703_934_reg_12845 - data_59_V_read_3_reg_8724_pp0_iter16_reg);

assign sub_ln703_878_fu_7890_p2 = (sub_ln703_859_reg_12850 - data_59_V_read_3_reg_8724_pp0_iter16_reg);

assign sub_ln703_879_fu_7735_p2 = (sub_ln703_860_fu_7620_p2 - data_59_V_read_3_reg_8724_pp0_iter15_reg);

assign sub_ln703_87_fu_1238_p2 = (add_ln703_184_fu_1143_p2 - data_9_V_read_8_reg_10136_pp0_iter4_reg);

assign sub_ln703_880_fu_7750_p2 = (sub_ln703_861_fu_7625_p2 - data_59_V_read_3_reg_8724_pp0_iter15_reg);

assign sub_ln703_881_fu_7755_p2 = (add_ln703_935_fu_7629_p2 - data_59_V_read_3_reg_8724_pp0_iter15_reg);

assign sub_ln703_882_fu_7894_p2 = (add_ln703_936_reg_12855 - data_59_V_read_3_reg_8724_pp0_iter16_reg);

assign sub_ln703_883_fu_7898_p2 = (sub_ln703_863_reg_12860 - data_59_V_read_3_reg_8724_pp0_iter16_reg);

assign sub_ln703_884_fu_7902_p2 = (sub_ln703_865_reg_12865 - data_59_V_read_3_reg_8724_pp0_iter16_reg);

assign sub_ln703_885_fu_7906_p2 = (sub_ln703_866_reg_12870 - data_59_V_read_3_reg_8724_pp0_iter16_reg);

assign sub_ln703_886_fu_7910_p2 = (add_ln703_938_reg_12875 - data_59_V_read_3_reg_8724_pp0_iter16_reg);

assign sub_ln703_887_fu_7914_p2 = (sub_ln703_867_reg_12880 - data_59_V_read_3_reg_8724_pp0_iter16_reg);

assign sub_ln703_888_fu_7918_p2 = (sub_ln703_868_reg_12885 - data_59_V_read_3_reg_8724_pp0_iter16_reg);

assign sub_ln703_889_fu_7922_p2 = (sub_ln703_869_reg_12800_pp0_iter16_reg - data_59_V_read_3_reg_8724_pp0_iter16_reg);

assign sub_ln703_88_fu_1248_p2 = (sub_ln703_73_reg_10611 - data_9_V_read_8_reg_10136_pp0_iter4_reg);

assign sub_ln703_890_fu_7926_p2 = (add_ln703_939_reg_12890 - data_59_V_read_3_reg_8724_pp0_iter16_reg);

assign sub_ln703_891_fu_7930_p2 = (sub_ln703_870_reg_12895 - data_59_V_read_3_reg_8724_pp0_iter16_reg);

assign sub_ln703_892_fu_7780_p2 = (add_ln703_940_fu_7690_p2 - data_59_V_read_3_reg_8724_pp0_iter15_reg);

assign sub_ln703_893_fu_7785_p2 = (sub_ln703_871_fu_7696_p2 - data_59_V_read_3_reg_8724_pp0_iter15_reg);

assign sub_ln703_894_fu_7790_p2 = (add_ln703_941_fu_7701_p2 - data_59_V_read_3_reg_8724_pp0_iter15_reg);

assign sub_ln703_895_fu_7795_p2 = (sub_ln703_872_fu_7705_p2 - data_59_V_read_3_reg_8724_pp0_iter15_reg);

assign sub_ln703_896_fu_7934_p2 = (sub_ln703_873_reg_12900 - data_59_V_read_3_reg_8724_pp0_iter16_reg);

assign sub_ln703_897_fu_7938_p2 = (add_ln703_943_reg_12905 - data_59_V_read_3_reg_8724_pp0_iter16_reg);

assign sub_ln703_898_fu_7805_p2 = (sub_ln703_874_fu_7725_p2 - data_59_V_read_3_reg_8724_pp0_iter15_reg);

assign sub_ln703_899_fu_7942_p2 = (sub_ln703_875_reg_12910 - data_59_V_read_3_reg_8724_pp0_iter16_reg);

assign sub_ln703_89_fu_1252_p2 = (sub_ln703_74_fu_1151_p2 - data_9_V_read_8_reg_10136_pp0_iter4_reg);

assign sub_ln703_8_fu_572_p2 = (sub_ln703_4_reg_10361 - data_3_V_read_10_reg_10295_pp0_iter1_reg);

assign sub_ln703_900_fu_7946_p2 = (sub_ln703_876_fu_7878_p2 - data_60_V_read61_reg_8691_pp0_iter16_reg);

assign sub_ln703_901_fu_7951_p2 = (add_ln703_944_fu_7882_p2 - data_60_V_read61_reg_8691_pp0_iter16_reg);

assign sub_ln703_902_fu_7961_p2 = (sub_ln703_878_fu_7890_p2 - data_60_V_read61_reg_8691_pp0_iter16_reg);

assign sub_ln703_903_fu_7966_p2 = (sub_ln703_879_reg_12915 - data_60_V_read61_reg_8691_pp0_iter16_reg);

assign sub_ln703_904_fu_7810_p2 = (add_ln703_947_fu_7745_p2 - data_60_V_read61_reg_8691_pp0_iter15_reg);

assign sub_ln703_905_fu_7970_p2 = (sub_ln703_880_reg_12920 - data_60_V_read61_reg_8691_pp0_iter16_reg);

assign sub_ln703_906_fu_7974_p2 = (sub_ln703_881_reg_12925 - data_60_V_read61_reg_8691_pp0_iter16_reg);

assign sub_ln703_907_fu_7978_p2 = (sub_ln703_883_fu_7898_p2 - data_60_V_read61_reg_8691_pp0_iter16_reg);

assign sub_ln703_908_fu_7983_p2 = (add_ln703_948_reg_12930 - data_60_V_read61_reg_8691_pp0_iter16_reg);

assign sub_ln703_909_fu_7987_p2 = (sub_ln703_885_fu_7906_p2 - data_60_V_read61_reg_8691_pp0_iter16_reg);

assign sub_ln703_90_fu_1257_p2 = (sub_ln703_75_reg_10616 - data_9_V_read_8_reg_10136_pp0_iter4_reg);

assign sub_ln703_910_fu_7992_p2 = (sub_ln703_888_fu_7918_p2 - data_60_V_read61_reg_8691_pp0_iter16_reg);

assign sub_ln703_911_fu_7833_p2 = (add_ln703_951_fu_7774_p2 - data_60_V_read61_reg_8691_pp0_iter15_reg);

assign sub_ln703_912_fu_8002_p2 = (sub_ln703_890_fu_7926_p2 - data_60_V_read61_reg_8691_pp0_iter16_reg);

assign sub_ln703_913_fu_8007_p2 = (sub_ln703_891_fu_7930_p2 - data_60_V_read61_reg_8691_pp0_iter16_reg);

assign sub_ln703_914_fu_8020_p2 = (sub_ln703_894_reg_12945 - data_60_V_read61_reg_8691_pp0_iter16_reg);

assign sub_ln703_915_fu_8024_p2 = (sub_ln703_895_reg_12950 - data_60_V_read61_reg_8691_pp0_iter16_reg);

assign sub_ln703_916_fu_8028_p2 = (sub_ln703_896_fu_7934_p2 - data_60_V_read61_reg_8691_pp0_iter16_reg);

assign sub_ln703_917_fu_7838_p2 = (add_ln703_952_fu_7800_p2 - data_60_V_read61_reg_8691_pp0_iter15_reg);

assign sub_ln703_918_fu_8033_p2 = (sub_ln703_898_reg_12955 - data_60_V_read61_reg_8691_pp0_iter16_reg);

assign sub_ln703_919_fu_8037_p2 = (add_ln703_953_fu_7956_p2 - data_61_V_read62_reg_8663_pp0_iter16_reg);

assign sub_ln703_91_fu_1261_p2 = (add_ln703_186_reg_10621 - data_9_V_read_8_reg_10136_pp0_iter4_reg);

assign sub_ln703_920_fu_8042_p2 = (sub_ln703_902_fu_7961_p2 - data_61_V_read62_reg_8663_pp0_iter16_reg);

assign sub_ln703_921_fu_8047_p2 = (sub_ln703_903_fu_7966_p2 - data_61_V_read62_reg_8663_pp0_iter16_reg);

assign sub_ln703_922_fu_7843_p2 = (add_ln703_955_fu_7815_p2 - data_61_V_read62_reg_8663_pp0_iter15_reg);

assign sub_ln703_923_fu_8057_p2 = (sub_ln703_906_fu_7974_p2 - data_61_V_read62_reg_8663_pp0_iter16_reg);

assign sub_ln703_924_fu_8072_p2 = (add_ln703_958_reg_12965 - data_61_V_read62_reg_8663_pp0_iter16_reg);

assign sub_ln703_925_fu_8076_p2 = (sub_ln703_911_reg_12970 - data_61_V_read62_reg_8663_pp0_iter16_reg);

assign sub_ln703_926_fu_8080_p2 = (add_ln703_959_fu_7997_p2 - data_61_V_read62_reg_8663_pp0_iter16_reg);

assign sub_ln703_927_fu_8085_p2 = (sub_ln703_913_fu_8007_p2 - data_61_V_read62_reg_8663_pp0_iter16_reg);

assign sub_ln703_928_fu_8090_p2 = (add_ln703_960_fu_8012_p2 - data_61_V_read62_reg_8663_pp0_iter16_reg);

assign sub_ln703_929_fu_8095_p2 = (add_ln703_961_fu_8016_p2 - data_61_V_read62_reg_8663_pp0_iter16_reg);

assign sub_ln703_92_fu_1054_p2 = (add_ln703_189_fu_1045_p2 - data_9_V_read_8_reg_10136_pp0_iter3_reg);

assign sub_ln703_930_fu_8120_p2 = (sub_ln703_921_fu_8047_p2 - data_62_V_read_3_reg_8645_pp0_iter16_reg);

assign sub_ln703_931_fu_8134_p2 = (add_ln703_962_fu_8052_p2 - data_62_V_read_3_reg_8645_pp0_iter16_reg);

assign sub_ln703_932_fu_8139_p2 = (sub_ln703_922_reg_12980 - data_62_V_read_3_reg_8645_pp0_iter16_reg);

assign sub_ln703_933_fu_8143_p2 = (sub_ln703_923_fu_8057_p2 - data_62_V_read_3_reg_8645_pp0_iter16_reg);

assign sub_ln703_934_fu_8165_p2 = (add_ln703_963_fu_8062_p2 - data_62_V_read_3_reg_8645_pp0_iter16_reg);

assign sub_ln703_935_fu_8181_p2 = (add_ln703_965_fu_8067_p2 - data_62_V_read_3_reg_8645_pp0_iter16_reg);

assign sub_ln703_936_fu_8209_p2 = (sub_ln703_928_fu_8090_p2 - data_62_V_read_3_reg_8645_pp0_iter16_reg);

assign sub_ln703_937_fu_8219_p2 = (add_ln703_966_fu_8100_p2 - data_62_V_read_3_reg_8645_pp0_iter16_reg);

assign sub_ln703_938_fu_8224_p2 = (add_ln703_967_fu_8105_p2 - data_62_V_read_3_reg_8645_pp0_iter16_reg);

assign sub_ln703_939_fu_8229_p2 = (add_ln703_968_fu_8110_p2 - data_62_V_read_3_reg_8645_pp0_iter16_reg);

assign sub_ln703_93_fu_1275_p2 = (sub_ln703_79_fu_1168_p2 - data_9_V_read_8_reg_10136_pp0_iter4_reg);

assign sub_ln703_940_fu_8234_p2 = (add_ln703_969_fu_8115_p2 - data_62_V_read_3_reg_8645_pp0_iter16_reg);

assign sub_ln703_94_fu_1280_p2 = (add_ln703_190_fu_1172_p2 - data_9_V_read_8_reg_10136_pp0_iter4_reg);

assign sub_ln703_95_fu_1285_p2 = (add_ln703_191_fu_1176_p2 - data_9_V_read_8_reg_10136_pp0_iter4_reg);

assign sub_ln703_96_fu_1294_p2 = (add_ln703_193_fu_1180_p2 - data_10_V_read11_reg_10105_pp0_iter4_reg);

assign sub_ln703_97_fu_1304_p2 = (add_ln703_194_fu_1189_p2 - data_10_V_read11_reg_10105_pp0_iter4_reg);

assign sub_ln703_98_fu_1319_p2 = (add_ln703_195_fu_1204_p2 - data_10_V_read11_reg_10105_pp0_iter4_reg);

assign sub_ln703_99_fu_1324_p2 = (add_ln703_197_fu_1209_p2 - data_10_V_read11_reg_10105_pp0_iter4_reg);

assign sub_ln703_9_fu_611_p2 = (sub_ln703_3_reg_10379 - data_3_V_read_10_reg_10295_pp0_iter2_reg);

assign sub_ln703_fu_536_p2 = (data_1_V_read_10_reg_10323 - data_0_V_read_10_reg_10329);

endmodule //dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_s
