
module normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1 (
        ap_clk,
        ap_rst,
        data_0_V_read,
        data_1_V_read,
        data_2_V_read,
        data_3_V_read,
        data_4_V_read,
        data_5_V_read,
        data_6_V_read,
        data_7_V_read,
        data_8_V_read,
        data_9_V_read,
        data_10_V_read,
        data_11_V_read,
        data_12_V_read,
        data_13_V_read,
        data_14_V_read,
        data_15_V_read,
        data_16_V_read,
        data_17_V_read,
        data_18_V_read,
        data_19_V_read,
        data_20_V_read,
        data_21_V_read,
        data_22_V_read,
        data_23_V_read,
        data_24_V_read,
        data_25_V_read,
        data_26_V_read,
        data_27_V_read,
        data_28_V_read,
        data_29_V_read,
        data_30_V_read,
        data_31_V_read,
        data_32_V_read,
        data_33_V_read,
        data_34_V_read,
        data_35_V_read,
        data_36_V_read,
        data_37_V_read,
        data_38_V_read,
        data_39_V_read,
        data_40_V_read,
        data_41_V_read,
        data_42_V_read,
        data_43_V_read,
        data_44_V_read,
        data_45_V_read,
        data_46_V_read,
        data_47_V_read,
        data_48_V_read,
        data_49_V_read,
        data_50_V_read,
        data_51_V_read,
        data_52_V_read,
        data_53_V_read,
        data_54_V_read,
        data_55_V_read,
        data_56_V_read,
        data_57_V_read,
        data_58_V_read,
        data_59_V_read,
        data_60_V_read,
        data_61_V_read,
        data_62_V_read,
        data_63_V_read,
        ap_return_0,
        ap_return_1,
        ap_return_2,
        ap_return_3,
        ap_return_4,
        ap_return_5,
        ap_return_6,
        ap_return_7,
        ap_return_8,
        ap_return_9,
        ap_return_10,
        ap_return_11,
        ap_return_12,
        ap_return_13,
        ap_return_14,
        ap_return_15,
        ap_return_16,
        ap_return_17,
        ap_return_18,
        ap_return_19,
        ap_return_20,
        ap_return_21,
        ap_return_22,
        ap_return_23,
        ap_return_24,
        ap_return_25,
        ap_return_26,
        ap_return_27,
        ap_return_28,
        ap_return_29,
        ap_return_30,
        ap_return_31,
        ap_return_32,
        ap_return_33,
        ap_return_34,
        ap_return_35,
        ap_return_36,
        ap_return_37,
        ap_return_38,
        ap_return_39,
        ap_return_40,
        ap_return_41,
        ap_return_42,
        ap_return_43,
        ap_return_44,
        ap_return_45,
        ap_return_46,
        ap_return_47,
        ap_return_48,
        ap_return_49,
        ap_return_50,
        ap_return_51,
        ap_return_52,
        ap_return_53,
        ap_return_54,
        ap_return_55,
        ap_return_56,
        ap_return_57,
        ap_return_58,
        ap_return_59,
        ap_return_60,
        ap_return_61,
        ap_return_62,
        ap_return_63,
        ap_ce
);


input   ap_clk;
input   ap_rst;
input  [15:0] data_0_V_read;
input  [15:0] data_1_V_read;
input  [15:0] data_2_V_read;
input  [15:0] data_3_V_read;
input  [15:0] data_4_V_read;
input  [15:0] data_5_V_read;
input  [15:0] data_6_V_read;
input  [15:0] data_7_V_read;
input  [15:0] data_8_V_read;
input  [15:0] data_9_V_read;
input  [15:0] data_10_V_read;
input  [15:0] data_11_V_read;
input  [15:0] data_12_V_read;
input  [15:0] data_13_V_read;
input  [15:0] data_14_V_read;
input  [15:0] data_15_V_read;
input  [15:0] data_16_V_read;
input  [15:0] data_17_V_read;
input  [15:0] data_18_V_read;
input  [15:0] data_19_V_read;
input  [15:0] data_20_V_read;
input  [15:0] data_21_V_read;
input  [15:0] data_22_V_read;
input  [15:0] data_23_V_read;
input  [15:0] data_24_V_read;
input  [15:0] data_25_V_read;
input  [15:0] data_26_V_read;
input  [15:0] data_27_V_read;
input  [15:0] data_28_V_read;
input  [15:0] data_29_V_read;
input  [15:0] data_30_V_read;
input  [15:0] data_31_V_read;
input  [15:0] data_32_V_read;
input  [15:0] data_33_V_read;
input  [15:0] data_34_V_read;
input  [15:0] data_35_V_read;
input  [15:0] data_36_V_read;
input  [15:0] data_37_V_read;
input  [15:0] data_38_V_read;
input  [15:0] data_39_V_read;
input  [15:0] data_40_V_read;
input  [15:0] data_41_V_read;
input  [15:0] data_42_V_read;
input  [15:0] data_43_V_read;
input  [15:0] data_44_V_read;
input  [15:0] data_45_V_read;
input  [15:0] data_46_V_read;
input  [15:0] data_47_V_read;
input  [15:0] data_48_V_read;
input  [15:0] data_49_V_read;
input  [15:0] data_50_V_read;
input  [15:0] data_51_V_read;
input  [15:0] data_52_V_read;
input  [15:0] data_53_V_read;
input  [15:0] data_54_V_read;
input  [15:0] data_55_V_read;
input  [15:0] data_56_V_read;
input  [15:0] data_57_V_read;
input  [15:0] data_58_V_read;
input  [15:0] data_59_V_read;
input  [15:0] data_60_V_read;
input  [15:0] data_61_V_read;
input  [15:0] data_62_V_read;
input  [15:0] data_63_V_read;
output  [15:0] ap_return_0;
output  [15:0] ap_return_1;
output  [15:0] ap_return_2;
output  [15:0] ap_return_3;
output  [15:0] ap_return_4;
output  [15:0] ap_return_5;
output  [15:0] ap_return_6;
output  [15:0] ap_return_7;
output  [15:0] ap_return_8;
output  [15:0] ap_return_9;
output  [15:0] ap_return_10;
output  [15:0] ap_return_11;
output  [15:0] ap_return_12;
output  [15:0] ap_return_13;
output  [15:0] ap_return_14;
output  [15:0] ap_return_15;
output  [15:0] ap_return_16;
output  [15:0] ap_return_17;
output  [15:0] ap_return_18;
output  [15:0] ap_return_19;
output  [15:0] ap_return_20;
output  [15:0] ap_return_21;
output  [15:0] ap_return_22;
output  [15:0] ap_return_23;
output  [15:0] ap_return_24;
output  [15:0] ap_return_25;
output  [15:0] ap_return_26;
output  [15:0] ap_return_27;
output  [15:0] ap_return_28;
output  [15:0] ap_return_29;
output  [15:0] ap_return_30;
output  [15:0] ap_return_31;
output  [15:0] ap_return_32;
output  [15:0] ap_return_33;
output  [15:0] ap_return_34;
output  [15:0] ap_return_35;
output  [15:0] ap_return_36;
output  [15:0] ap_return_37;
output  [15:0] ap_return_38;
output  [15:0] ap_return_39;
output  [15:0] ap_return_40;
output  [15:0] ap_return_41;
output  [15:0] ap_return_42;
output  [15:0] ap_return_43;
output  [15:0] ap_return_44;
output  [15:0] ap_return_45;
output  [15:0] ap_return_46;
output  [15:0] ap_return_47;
output  [15:0] ap_return_48;
output  [15:0] ap_return_49;
output  [15:0] ap_return_50;
output  [15:0] ap_return_51;
output  [15:0] ap_return_52;
output  [15:0] ap_return_53;
output  [15:0] ap_return_54;
output  [15:0] ap_return_55;
output  [15:0] ap_return_56;
output  [15:0] ap_return_57;
output  [15:0] ap_return_58;
output  [15:0] ap_return_59;
output  [15:0] ap_return_60;
output  [15:0] ap_return_61;
output  [15:0] ap_return_62;
output  [15:0] ap_return_63;
input   ap_ce;

reg[15:0] ap_return_0;
reg[15:0] ap_return_1;
reg[15:0] ap_return_2;
reg[15:0] ap_return_3;
reg[15:0] ap_return_4;
reg[15:0] ap_return_5;
reg[15:0] ap_return_6;
reg[15:0] ap_return_7;
reg[15:0] ap_return_8;
reg[15:0] ap_return_9;
reg[15:0] ap_return_10;
reg[15:0] ap_return_11;
reg[15:0] ap_return_12;
reg[15:0] ap_return_13;
reg[15:0] ap_return_14;
reg[15:0] ap_return_15;
reg[15:0] ap_return_16;
reg[15:0] ap_return_17;
reg[15:0] ap_return_18;
reg[15:0] ap_return_19;
reg[15:0] ap_return_20;
reg[15:0] ap_return_21;
reg[15:0] ap_return_22;
reg[15:0] ap_return_23;
reg[15:0] ap_return_24;
reg[15:0] ap_return_25;
reg[15:0] ap_return_26;
reg[15:0] ap_return_27;
reg[15:0] ap_return_28;
reg[15:0] ap_return_29;
reg[15:0] ap_return_30;
reg[15:0] ap_return_31;
reg[15:0] ap_return_32;
reg[15:0] ap_return_33;
reg[15:0] ap_return_34;
reg[15:0] ap_return_35;
reg[15:0] ap_return_36;
reg[15:0] ap_return_37;
reg[15:0] ap_return_38;
reg[15:0] ap_return_39;
reg[15:0] ap_return_40;
reg[15:0] ap_return_41;
reg[15:0] ap_return_42;
reg[15:0] ap_return_43;
reg[15:0] ap_return_44;
reg[15:0] ap_return_45;
reg[15:0] ap_return_46;
reg[15:0] ap_return_47;
reg[15:0] ap_return_48;
reg[15:0] ap_return_49;
reg[15:0] ap_return_50;
reg[15:0] ap_return_51;
reg[15:0] ap_return_52;
reg[15:0] ap_return_53;
reg[15:0] ap_return_54;
reg[15:0] ap_return_55;
reg[15:0] ap_return_56;
reg[15:0] ap_return_57;
reg[15:0] ap_return_58;
reg[15:0] ap_return_59;
reg[15:0] ap_return_60;
reg[15:0] ap_return_61;
reg[15:0] ap_return_62;
reg[15:0] ap_return_63;

reg   [15:0] data_46_V_read_2_reg_18625;
wire    ap_block_state1_pp0_stage0_iter0;
wire    ap_block_state2_pp0_stage0_iter1;
wire    ap_block_state3_pp0_stage0_iter2;
wire    ap_block_pp0_stage0_11001;
reg   [15:0] data_42_V_read_2_reg_18631;
reg   [15:0] data_39_V_read_2_reg_18637;
reg   [15:0] trunc_ln_reg_18948;
reg   [15:0] trunc_ln708_31_reg_18953;
reg   [15:0] trunc_ln708_32_reg_18958;
reg   [15:0] trunc_ln708_s_reg_18963;
reg   [15:0] trunc_ln708_33_reg_18968;
reg   [15:0] trunc_ln708_34_reg_18973;
reg   [15:0] trunc_ln708_35_reg_18978;
reg   [15:0] trunc_ln708_36_reg_18983;
reg   [15:0] trunc_ln708_37_reg_18988;
reg   [15:0] trunc_ln708_38_reg_18993;
reg   [15:0] trunc_ln708_39_reg_18998;
reg   [15:0] trunc_ln708_40_reg_19003;
reg   [15:0] trunc_ln708_41_reg_19008;
reg   [15:0] trunc_ln708_42_reg_19013;
reg   [15:0] trunc_ln708_43_reg_19018;
reg   [15:0] trunc_ln708_44_reg_19023;
reg   [15:0] trunc_ln708_45_reg_19028;
reg   [15:0] trunc_ln708_46_reg_19033;
reg   [15:0] trunc_ln708_47_reg_19038;
reg   [15:0] trunc_ln708_48_reg_19043;
reg   [15:0] trunc_ln708_49_reg_19048;
reg   [15:0] trunc_ln708_50_reg_19053;
reg   [15:0] trunc_ln708_51_reg_19058;
reg   [15:0] trunc_ln708_52_reg_19063;
reg   [15:0] trunc_ln708_53_reg_19068;
reg   [15:0] trunc_ln708_54_reg_19073;
reg   [15:0] trunc_ln708_55_reg_19078;
reg   [15:0] trunc_ln708_56_reg_19083;
reg   [15:0] trunc_ln708_57_reg_19088;
reg   [15:0] trunc_ln708_58_reg_19093;
reg   [15:0] trunc_ln708_59_reg_19098;
reg   [15:0] trunc_ln708_60_reg_19103;
reg   [15:0] trunc_ln708_61_reg_19108;
reg   [15:0] trunc_ln708_62_reg_19113;
reg   [15:0] trunc_ln708_63_reg_19118;
reg   [15:0] trunc_ln708_64_reg_19123;
reg   [15:0] trunc_ln708_65_reg_19128;
reg   [15:0] trunc_ln708_66_reg_19133;
reg   [15:0] trunc_ln708_67_reg_19138;
reg   [15:0] trunc_ln708_68_reg_19143;
reg   [15:0] trunc_ln708_69_reg_19148;
reg   [15:0] trunc_ln708_70_reg_19153;
reg   [15:0] trunc_ln708_71_reg_19158;
reg   [15:0] trunc_ln708_72_reg_19163;
reg   [15:0] trunc_ln708_73_reg_19168;
reg   [15:0] trunc_ln708_74_reg_19173;
reg   [15:0] trunc_ln708_75_reg_19178;
reg   [15:0] trunc_ln708_76_reg_19183;
reg   [15:0] trunc_ln708_77_reg_19188;
reg   [15:0] trunc_ln708_78_reg_19193;
reg   [15:0] trunc_ln708_79_reg_19198;
reg   [15:0] trunc_ln708_80_reg_19203;
reg   [15:0] trunc_ln708_81_reg_19208;
reg   [15:0] trunc_ln708_82_reg_19213;
reg   [15:0] trunc_ln708_83_reg_19218;
reg   [15:0] trunc_ln708_84_reg_19223;
reg   [15:0] trunc_ln708_85_reg_19228;
reg   [15:0] trunc_ln708_86_reg_19233;
reg   [15:0] trunc_ln708_87_reg_19238;
reg   [15:0] trunc_ln708_88_reg_19243;
reg   [15:0] trunc_ln708_89_reg_19248;
reg   [15:0] trunc_ln708_90_reg_19253;
reg   [15:0] trunc_ln708_91_reg_19258;
reg   [15:0] trunc_ln708_92_reg_19263;
wire   [11:0] grp_fu_804_p1;
wire    ap_block_pp0_stage0;
wire   [11:0] grp_fu_805_p1;
wire   [11:0] grp_fu_806_p1;
wire   [11:0] grp_fu_807_p1;
wire   [10:0] grp_fu_808_p1;
wire   [10:0] grp_fu_809_p1;
wire   [11:0] grp_fu_810_p1;
wire   [10:0] grp_fu_811_p1;
wire   [11:0] grp_fu_812_p1;
wire   [12:0] grp_fu_813_p1;
wire   [11:0] grp_fu_814_p1;
wire   [11:0] grp_fu_815_p1;
wire   [11:0] grp_fu_816_p1;
wire   [11:0] grp_fu_818_p1;
wire   [10:0] grp_fu_819_p1;
wire   [11:0] grp_fu_820_p1;
wire   [11:0] grp_fu_821_p1;
wire   [11:0] grp_fu_822_p1;
wire   [11:0] grp_fu_823_p1;
wire   [11:0] grp_fu_824_p1;
wire   [10:0] grp_fu_825_p1;
wire   [11:0] grp_fu_826_p1;
wire   [11:0] grp_fu_827_p1;
wire   [10:0] grp_fu_828_p1;
wire   [10:0] grp_fu_829_p1;
wire   [11:0] grp_fu_830_p1;
wire   [10:0] grp_fu_831_p1;
wire   [10:0] grp_fu_832_p1;
wire   [11:0] grp_fu_833_p1;
wire   [10:0] grp_fu_834_p1;
wire   [11:0] grp_fu_835_p1;
wire   [11:0] grp_fu_837_p1;
wire   [12:0] grp_fu_838_p1;
wire   [10:0] grp_fu_839_p1;
wire   [11:0] grp_fu_840_p1;
wire   [10:0] grp_fu_841_p1;
wire   [11:0] grp_fu_842_p1;
wire   [10:0] grp_fu_843_p1;
wire   [10:0] grp_fu_844_p1;
wire   [10:0] grp_fu_845_p1;
wire   [11:0] grp_fu_846_p1;
wire   [11:0] grp_fu_847_p1;
wire   [10:0] grp_fu_848_p1;
wire   [11:0] grp_fu_849_p1;
wire   [10:0] grp_fu_850_p1;
wire   [11:0] grp_fu_851_p1;
wire   [11:0] grp_fu_852_p1;
wire   [10:0] grp_fu_853_p1;
wire   [12:0] grp_fu_854_p1;
wire   [11:0] grp_fu_855_p1;
wire   [10:0] grp_fu_856_p1;
wire   [11:0] grp_fu_857_p1;
wire   [10:0] grp_fu_858_p1;
wire   [11:0] grp_fu_859_p1;
wire   [11:0] grp_fu_860_p1;
wire   [11:0] grp_fu_861_p1;
wire   [11:0] grp_fu_862_p1;
wire   [11:0] grp_fu_863_p1;
wire   [10:0] grp_fu_864_p1;
wire   [11:0] grp_fu_866_p1;
wire   [12:0] grp_fu_867_p1;
wire   [25:0] grp_fu_852_p2;
wire   [25:0] grp_fu_832_p2;
wire   [25:0] grp_fu_860_p2;
wire   [25:0] grp_fu_828_p2;
wire   [25:0] grp_fu_857_p2;
wire   [25:0] grp_fu_846_p2;
wire   [25:0] grp_fu_829_p2;
wire   [25:0] grp_fu_866_p2;
wire   [25:0] grp_fu_819_p2;
wire   [25:0] grp_fu_844_p2;
wire   [25:0] grp_fu_859_p2;
wire   [25:0] grp_fu_856_p2;
wire   [25:0] grp_fu_834_p2;
wire   [25:0] grp_fu_813_p2;
wire   [25:0] grp_fu_816_p2;
wire   [25:0] grp_fu_812_p2;
wire   [25:0] grp_fu_837_p2;
wire   [25:0] grp_fu_849_p2;
wire   [25:0] grp_fu_818_p2;
wire   [25:0] grp_fu_810_p2;
wire   [25:0] grp_fu_815_p2;
wire   [25:0] grp_fu_811_p2;
wire   [25:0] grp_fu_824_p2;
wire   [25:0] grp_fu_830_p2;
wire   [25:0] grp_fu_839_p2;
wire   [25:0] grp_fu_850_p2;
wire   [25:0] grp_fu_827_p2;
wire   [25:0] grp_fu_847_p2;
wire   [25:0] grp_fu_845_p2;
wire   [25:0] grp_fu_853_p2;
wire   [25:0] grp_fu_814_p2;
wire   [25:0] grp_fu_840_p2;
wire   [25:0] grp_fu_808_p2;
wire   [25:0] grp_fu_858_p2;
wire   [25:0] grp_fu_835_p2;
wire   [25:0] grp_fu_804_p2;
wire   [25:0] grp_fu_841_p2;
wire   [25:0] grp_fu_807_p2;
wire   [25:0] grp_fu_825_p2;
wire   [22:0] shl_ln1118_5_fu_17614_p3;
wire   [25:0] shl_ln_fu_17607_p3;
wire   [25:0] sext_ln1118_73_fu_17621_p1;
wire   [25:0] add_ln1118_fu_17625_p2;
wire   [25:0] grp_fu_867_p2;
wire   [25:0] grp_fu_822_p2;
wire   [25:0] sext_ln1118_76_fu_17661_p1;
wire   [25:0] shl_ln1118_6_fu_17664_p3;
wire   [25:0] add_ln1118_1_fu_17671_p2;
wire   [25:0] grp_fu_851_p2;
wire   [25:0] grp_fu_826_p2;
wire   [25:0] grp_fu_855_p2;
wire   [21:0] shl_ln1118_8_fu_17724_p3;
wire   [25:0] shl_ln1118_7_fu_17717_p3;
wire   [25:0] sext_ln1118_80_fu_17731_p1;
wire   [25:0] add_ln1118_2_fu_17735_p2;
wire   [25:0] grp_fu_838_p2;
wire   [25:0] grp_fu_861_p2;
wire   [25:0] grp_fu_843_p2;
wire   [25:0] grp_fu_862_p2;
wire   [25:0] grp_fu_863_p2;
wire   [25:0] grp_fu_823_p2;
wire   [25:0] grp_fu_848_p2;
wire   [25:0] grp_fu_854_p2;
wire   [25:0] grp_fu_821_p2;
wire   [25:0] grp_fu_831_p2;
wire   [25:0] grp_fu_864_p2;
wire   [25:0] grp_fu_809_p2;
wire   [25:0] grp_fu_842_p2;
wire   [25:0] grp_fu_805_p2;
wire   [25:0] grp_fu_833_p2;
wire   [25:0] grp_fu_806_p2;
wire   [25:0] grp_fu_820_p2;
wire   [15:0] add_ln703_fu_17921_p2;
wire   [15:0] add_ln703_36_fu_17926_p2;
wire   [15:0] add_ln703_37_fu_17931_p2;
wire   [15:0] add_ln703_38_fu_17936_p2;
wire   [15:0] add_ln703_39_fu_17941_p2;
wire   [15:0] add_ln703_40_fu_17946_p2;
wire   [15:0] add_ln703_41_fu_17951_p2;
wire   [15:0] add_ln703_42_fu_17956_p2;
wire   [15:0] add_ln703_43_fu_17961_p2;
wire   [15:0] add_ln703_44_fu_17966_p2;
wire   [15:0] add_ln703_45_fu_17971_p2;
wire   [15:0] add_ln703_46_fu_17976_p2;
wire   [15:0] add_ln703_47_fu_17981_p2;
wire   [15:0] add_ln703_48_fu_17986_p2;
wire   [15:0] add_ln703_49_fu_17991_p2;
wire   [15:0] add_ln703_50_fu_17996_p2;
wire   [15:0] add_ln703_51_fu_18001_p2;
wire   [15:0] add_ln703_52_fu_18006_p2;
wire   [15:0] add_ln703_53_fu_18011_p2;
wire   [15:0] add_ln703_54_fu_18016_p2;
wire   [15:0] add_ln703_55_fu_18021_p2;
wire   [15:0] add_ln703_56_fu_18026_p2;
wire   [15:0] add_ln703_57_fu_18031_p2;
wire   [15:0] add_ln703_58_fu_18036_p2;
wire   [15:0] add_ln703_59_fu_18041_p2;
wire   [15:0] add_ln703_60_fu_18046_p2;
wire   [15:0] add_ln703_61_fu_18051_p2;
wire   [15:0] add_ln703_62_fu_18056_p2;
wire   [15:0] add_ln703_63_fu_18061_p2;
wire   [15:0] add_ln703_64_fu_18066_p2;
wire   [15:0] add_ln703_65_fu_18071_p2;
wire   [15:0] add_ln703_66_fu_18076_p2;
wire   [15:0] add_ln703_67_fu_18081_p2;
wire   [15:0] add_ln703_68_fu_18086_p2;
wire   [15:0] add_ln703_69_fu_18091_p2;
wire   [15:0] add_ln703_70_fu_18096_p2;
wire   [15:0] add_ln703_71_fu_18101_p2;
wire   [15:0] add_ln703_72_fu_18106_p2;
wire   [15:0] add_ln703_73_fu_18111_p2;
wire   [15:0] add_ln703_74_fu_18116_p2;
wire   [15:0] add_ln703_75_fu_18121_p2;
wire   [15:0] add_ln703_76_fu_18126_p2;
wire   [15:0] add_ln703_77_fu_18131_p2;
wire   [15:0] add_ln703_78_fu_18136_p2;
wire   [15:0] add_ln703_79_fu_18141_p2;
wire   [15:0] add_ln703_80_fu_18146_p2;
wire   [15:0] add_ln703_81_fu_18151_p2;
wire   [15:0] add_ln703_82_fu_18156_p2;
wire   [15:0] add_ln703_83_fu_18161_p2;
wire   [15:0] add_ln703_84_fu_18166_p2;
wire   [15:0] add_ln703_85_fu_18171_p2;
wire   [15:0] add_ln703_86_fu_18176_p2;
wire   [15:0] add_ln703_87_fu_18181_p2;
wire   [15:0] add_ln703_88_fu_18186_p2;
wire   [15:0] add_ln703_89_fu_18191_p2;
wire   [15:0] add_ln703_90_fu_18196_p2;
wire   [15:0] add_ln703_91_fu_18201_p2;
wire   [15:0] add_ln703_92_fu_18206_p2;
wire   [15:0] add_ln703_93_fu_18211_p2;
wire   [15:0] add_ln703_94_fu_18216_p2;
wire   [15:0] add_ln703_95_fu_18221_p2;
wire   [15:0] add_ln703_96_fu_18226_p2;
wire   [15:0] add_ln703_97_fu_18231_p2;
wire   [15:0] add_ln703_98_fu_18236_p2;
reg    grp_fu_804_ce;
reg    grp_fu_805_ce;
reg    grp_fu_806_ce;
reg    grp_fu_807_ce;
reg    grp_fu_808_ce;
reg    grp_fu_809_ce;
reg    grp_fu_810_ce;
reg    grp_fu_811_ce;
reg    grp_fu_812_ce;
reg    grp_fu_813_ce;
reg    grp_fu_814_ce;
reg    grp_fu_815_ce;
reg    grp_fu_816_ce;
reg    grp_fu_818_ce;
reg    grp_fu_819_ce;
reg    grp_fu_820_ce;
reg    grp_fu_821_ce;
reg    grp_fu_822_ce;
reg    grp_fu_823_ce;
reg    grp_fu_824_ce;
reg    grp_fu_825_ce;
reg    grp_fu_826_ce;
reg    grp_fu_827_ce;
reg    grp_fu_828_ce;
reg    grp_fu_829_ce;
reg    grp_fu_830_ce;
reg    grp_fu_831_ce;
reg    grp_fu_832_ce;
reg    grp_fu_833_ce;
reg    grp_fu_834_ce;
reg    grp_fu_835_ce;
reg    grp_fu_837_ce;
reg    grp_fu_838_ce;
reg    grp_fu_839_ce;
reg    grp_fu_840_ce;
reg    grp_fu_841_ce;
reg    grp_fu_842_ce;
reg    grp_fu_843_ce;
reg    grp_fu_844_ce;
reg    grp_fu_845_ce;
reg    grp_fu_846_ce;
reg    grp_fu_847_ce;
reg    grp_fu_848_ce;
reg    grp_fu_849_ce;
reg    grp_fu_850_ce;
reg    grp_fu_851_ce;
reg    grp_fu_852_ce;
reg    grp_fu_853_ce;
reg    grp_fu_854_ce;
reg    grp_fu_855_ce;
reg    grp_fu_856_ce;
reg    grp_fu_857_ce;
reg    grp_fu_858_ce;
reg    grp_fu_859_ce;
reg    grp_fu_860_ce;
reg    grp_fu_861_ce;
reg    grp_fu_862_ce;
reg    grp_fu_863_ce;
reg    grp_fu_864_ce;
reg    grp_fu_866_ce;
reg    grp_fu_867_ce;
reg    ap_ce_reg;
reg   [15:0] data_0_V_read_int_reg;
reg   [15:0] data_1_V_read_int_reg;
reg   [15:0] data_2_V_read_int_reg;
reg   [15:0] data_3_V_read_int_reg;
reg   [15:0] data_4_V_read_int_reg;
reg   [15:0] data_5_V_read_int_reg;
reg   [15:0] data_6_V_read_int_reg;
reg   [15:0] data_7_V_read_int_reg;
reg   [15:0] data_8_V_read_int_reg;
reg   [15:0] data_9_V_read_int_reg;
reg   [15:0] data_10_V_read_int_reg;
reg   [15:0] data_11_V_read_int_reg;
reg   [15:0] data_12_V_read_int_reg;
reg   [15:0] data_13_V_read_int_reg;
reg   [15:0] data_14_V_read_int_reg;
reg   [15:0] data_15_V_read_int_reg;
reg   [15:0] data_16_V_read_int_reg;
reg   [15:0] data_17_V_read_int_reg;
reg   [15:0] data_18_V_read_int_reg;
reg   [15:0] data_19_V_read_int_reg;
reg   [15:0] data_20_V_read_int_reg;
reg   [15:0] data_21_V_read_int_reg;
reg   [15:0] data_22_V_read_int_reg;
reg   [15:0] data_23_V_read_int_reg;
reg   [15:0] data_24_V_read_int_reg;
reg   [15:0] data_25_V_read_int_reg;
reg   [15:0] data_26_V_read_int_reg;
reg   [15:0] data_27_V_read_int_reg;
reg   [15:0] data_28_V_read_int_reg;
reg   [15:0] data_29_V_read_int_reg;
reg   [15:0] data_30_V_read_int_reg;
reg   [15:0] data_31_V_read_int_reg;
reg   [15:0] data_32_V_read_int_reg;
reg   [15:0] data_33_V_read_int_reg;
reg   [15:0] data_34_V_read_int_reg;
reg   [15:0] data_35_V_read_int_reg;
reg   [15:0] data_36_V_read_int_reg;
reg   [15:0] data_37_V_read_int_reg;
reg   [15:0] data_38_V_read_int_reg;
reg   [15:0] data_39_V_read_int_reg;
reg   [15:0] data_40_V_read_int_reg;
reg   [15:0] data_41_V_read_int_reg;
reg   [15:0] data_42_V_read_int_reg;
reg   [15:0] data_43_V_read_int_reg;
reg   [15:0] data_44_V_read_int_reg;
reg   [15:0] data_45_V_read_int_reg;
reg   [15:0] data_46_V_read_int_reg;
reg   [15:0] data_47_V_read_int_reg;
reg   [15:0] data_48_V_read_int_reg;
reg   [15:0] data_49_V_read_int_reg;
reg   [15:0] data_50_V_read_int_reg;
reg   [15:0] data_51_V_read_int_reg;
reg   [15:0] data_52_V_read_int_reg;
reg   [15:0] data_53_V_read_int_reg;
reg   [15:0] data_54_V_read_int_reg;
reg   [15:0] data_55_V_read_int_reg;
reg   [15:0] data_56_V_read_int_reg;
reg   [15:0] data_57_V_read_int_reg;
reg   [15:0] data_58_V_read_int_reg;
reg   [15:0] data_59_V_read_int_reg;
reg   [15:0] data_60_V_read_int_reg;
reg   [15:0] data_61_V_read_int_reg;
reg   [15:0] data_62_V_read_int_reg;
reg   [15:0] data_63_V_read_int_reg;
reg   [15:0] ap_return_0_int_reg;
reg   [15:0] ap_return_1_int_reg;
reg   [15:0] ap_return_2_int_reg;
reg   [15:0] ap_return_3_int_reg;
reg   [15:0] ap_return_4_int_reg;
reg   [15:0] ap_return_5_int_reg;
reg   [15:0] ap_return_6_int_reg;
reg   [15:0] ap_return_7_int_reg;
reg   [15:0] ap_return_8_int_reg;
reg   [15:0] ap_return_9_int_reg;
reg   [15:0] ap_return_10_int_reg;
reg   [15:0] ap_return_11_int_reg;
reg   [15:0] ap_return_12_int_reg;
reg   [15:0] ap_return_13_int_reg;
reg   [15:0] ap_return_14_int_reg;
reg   [15:0] ap_return_15_int_reg;
reg   [15:0] ap_return_16_int_reg;
reg   [15:0] ap_return_17_int_reg;
reg   [15:0] ap_return_18_int_reg;
reg   [15:0] ap_return_19_int_reg;
reg   [15:0] ap_return_20_int_reg;
reg   [15:0] ap_return_21_int_reg;
reg   [15:0] ap_return_22_int_reg;
reg   [15:0] ap_return_23_int_reg;
reg   [15:0] ap_return_24_int_reg;
reg   [15:0] ap_return_25_int_reg;
reg   [15:0] ap_return_26_int_reg;
reg   [15:0] ap_return_27_int_reg;
reg   [15:0] ap_return_28_int_reg;
reg   [15:0] ap_return_29_int_reg;
reg   [15:0] ap_return_30_int_reg;
reg   [15:0] ap_return_31_int_reg;
reg   [15:0] ap_return_32_int_reg;
reg   [15:0] ap_return_33_int_reg;
reg   [15:0] ap_return_34_int_reg;
reg   [15:0] ap_return_35_int_reg;
reg   [15:0] ap_return_36_int_reg;
reg   [15:0] ap_return_37_int_reg;
reg   [15:0] ap_return_38_int_reg;
reg   [15:0] ap_return_39_int_reg;
reg   [15:0] ap_return_40_int_reg;
reg   [15:0] ap_return_41_int_reg;
reg   [15:0] ap_return_42_int_reg;
reg   [15:0] ap_return_43_int_reg;
reg   [15:0] ap_return_44_int_reg;
reg   [15:0] ap_return_45_int_reg;
reg   [15:0] ap_return_46_int_reg;
reg   [15:0] ap_return_47_int_reg;
reg   [15:0] ap_return_48_int_reg;
reg   [15:0] ap_return_49_int_reg;
reg   [15:0] ap_return_50_int_reg;
reg   [15:0] ap_return_51_int_reg;
reg   [15:0] ap_return_52_int_reg;
reg   [15:0] ap_return_53_int_reg;
reg   [15:0] ap_return_54_int_reg;
reg   [15:0] ap_return_55_int_reg;
reg   [15:0] ap_return_56_int_reg;
reg   [15:0] ap_return_57_int_reg;
reg   [15:0] ap_return_58_int_reg;
reg   [15:0] ap_return_59_int_reg;
reg   [15:0] ap_return_60_int_reg;
reg   [15:0] ap_return_61_int_reg;
reg   [15:0] ap_return_62_int_reg;
reg   [15:0] ap_return_63_int_reg;

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U2(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_35_V_read_int_reg),
    .din1(grp_fu_804_p1),
    .ce(grp_fu_804_ce),
    .dout(grp_fu_804_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U3(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_60_V_read_int_reg),
    .din1(grp_fu_805_p1),
    .ce(grp_fu_805_ce),
    .dout(grp_fu_805_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U4(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_62_V_read_int_reg),
    .din1(grp_fu_806_p1),
    .ce(grp_fu_806_ce),
    .dout(grp_fu_806_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U5(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_37_V_read_int_reg),
    .din1(grp_fu_807_p1),
    .ce(grp_fu_807_ce),
    .dout(grp_fu_807_p2)
);

myproject_mul_16s_11ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_11ns_26_2_0_U6(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_32_V_read_int_reg),
    .din1(grp_fu_808_p1),
    .ce(grp_fu_808_ce),
    .dout(grp_fu_808_p2)
);

myproject_mul_16s_11ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_11ns_26_2_0_U7(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_58_V_read_int_reg),
    .din1(grp_fu_809_p1),
    .ce(grp_fu_809_ce),
    .dout(grp_fu_809_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U8(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_19_V_read_int_reg),
    .din1(grp_fu_810_p1),
    .ce(grp_fu_810_ce),
    .dout(grp_fu_810_p2)
);

myproject_mul_16s_11ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_11ns_26_2_0_U9(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_21_V_read_int_reg),
    .din1(grp_fu_811_p1),
    .ce(grp_fu_811_ce),
    .dout(grp_fu_811_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U10(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_15_V_read_int_reg),
    .din1(grp_fu_812_p1),
    .ce(grp_fu_812_ce),
    .dout(grp_fu_812_p2)
);

myproject_mul_16s_13ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 13 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_13ns_26_2_0_U11(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_13_V_read_int_reg),
    .din1(grp_fu_813_p1),
    .ce(grp_fu_813_ce),
    .dout(grp_fu_813_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U12(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_30_V_read_int_reg),
    .din1(grp_fu_814_p1),
    .ce(grp_fu_814_ce),
    .dout(grp_fu_814_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U13(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_20_V_read_int_reg),
    .din1(grp_fu_815_p1),
    .ce(grp_fu_815_ce),
    .dout(grp_fu_815_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U14(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_14_V_read_int_reg),
    .din1(grp_fu_816_p1),
    .ce(grp_fu_816_ce),
    .dout(grp_fu_816_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U15(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_18_V_read_int_reg),
    .din1(grp_fu_818_p1),
    .ce(grp_fu_818_ce),
    .dout(grp_fu_818_p2)
);

myproject_mul_16s_11ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_11ns_26_2_0_U16(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_8_V_read_int_reg),
    .din1(grp_fu_819_p1),
    .ce(grp_fu_819_ce),
    .dout(grp_fu_819_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U17(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_63_V_read_int_reg),
    .din1(grp_fu_820_p1),
    .ce(grp_fu_820_ce),
    .dout(grp_fu_820_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U18(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_55_V_read_int_reg),
    .din1(grp_fu_821_p1),
    .ce(grp_fu_821_ce),
    .dout(grp_fu_821_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U19(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_41_V_read_int_reg),
    .din1(grp_fu_822_p1),
    .ce(grp_fu_822_ce),
    .dout(grp_fu_822_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U20(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_52_V_read_int_reg),
    .din1(grp_fu_823_p1),
    .ce(grp_fu_823_ce),
    .dout(grp_fu_823_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U21(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_22_V_read_int_reg),
    .din1(grp_fu_824_p1),
    .ce(grp_fu_824_ce),
    .dout(grp_fu_824_p2)
);

myproject_mul_16s_11ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_11ns_26_2_0_U22(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_38_V_read_int_reg),
    .din1(grp_fu_825_p1),
    .ce(grp_fu_825_ce),
    .dout(grp_fu_825_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U23(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_44_V_read_int_reg),
    .din1(grp_fu_826_p1),
    .ce(grp_fu_826_ce),
    .dout(grp_fu_826_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U24(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_26_V_read_int_reg),
    .din1(grp_fu_827_p1),
    .ce(grp_fu_827_ce),
    .dout(grp_fu_827_p2)
);

myproject_mul_16s_11ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_11ns_26_2_0_U25(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_3_V_read_int_reg),
    .din1(grp_fu_828_p1),
    .ce(grp_fu_828_ce),
    .dout(grp_fu_828_p2)
);

myproject_mul_16s_11ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_11ns_26_2_0_U26(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_6_V_read_int_reg),
    .din1(grp_fu_829_p1),
    .ce(grp_fu_829_ce),
    .dout(grp_fu_829_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U27(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_23_V_read_int_reg),
    .din1(grp_fu_830_p1),
    .ce(grp_fu_830_ce),
    .dout(grp_fu_830_p2)
);

myproject_mul_16s_11ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_11ns_26_2_0_U28(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_56_V_read_int_reg),
    .din1(grp_fu_831_p1),
    .ce(grp_fu_831_ce),
    .dout(grp_fu_831_p2)
);

myproject_mul_16s_11ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_11ns_26_2_0_U29(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_1_V_read_int_reg),
    .din1(grp_fu_832_p1),
    .ce(grp_fu_832_ce),
    .dout(grp_fu_832_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U30(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_61_V_read_int_reg),
    .din1(grp_fu_833_p1),
    .ce(grp_fu_833_ce),
    .dout(grp_fu_833_p2)
);

myproject_mul_16s_11ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_11ns_26_2_0_U31(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_12_V_read_int_reg),
    .din1(grp_fu_834_p1),
    .ce(grp_fu_834_ce),
    .dout(grp_fu_834_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U32(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_34_V_read_int_reg),
    .din1(grp_fu_835_p1),
    .ce(grp_fu_835_ce),
    .dout(grp_fu_835_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U33(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_16_V_read_int_reg),
    .din1(grp_fu_837_p1),
    .ce(grp_fu_837_ce),
    .dout(grp_fu_837_p2)
);

myproject_mul_16s_13ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 13 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_13ns_26_2_0_U34(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_47_V_read_int_reg),
    .din1(grp_fu_838_p1),
    .ce(grp_fu_838_ce),
    .dout(grp_fu_838_p2)
);

myproject_mul_16s_11ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_11ns_26_2_0_U35(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_24_V_read_int_reg),
    .din1(grp_fu_839_p1),
    .ce(grp_fu_839_ce),
    .dout(grp_fu_839_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U36(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_31_V_read_int_reg),
    .din1(grp_fu_840_p1),
    .ce(grp_fu_840_ce),
    .dout(grp_fu_840_p2)
);

myproject_mul_16s_11ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_11ns_26_2_0_U37(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_36_V_read_int_reg),
    .din1(grp_fu_841_p1),
    .ce(grp_fu_841_ce),
    .dout(grp_fu_841_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U38(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_59_V_read_int_reg),
    .din1(grp_fu_842_p1),
    .ce(grp_fu_842_ce),
    .dout(grp_fu_842_p2)
);

myproject_mul_16s_11ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_11ns_26_2_0_U39(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_49_V_read_int_reg),
    .din1(grp_fu_843_p1),
    .ce(grp_fu_843_ce),
    .dout(grp_fu_843_p2)
);

myproject_mul_16s_11ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_11ns_26_2_0_U40(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_9_V_read_int_reg),
    .din1(grp_fu_844_p1),
    .ce(grp_fu_844_ce),
    .dout(grp_fu_844_p2)
);

myproject_mul_16s_11ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_11ns_26_2_0_U41(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_28_V_read_int_reg),
    .din1(grp_fu_845_p1),
    .ce(grp_fu_845_ce),
    .dout(grp_fu_845_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U42(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_5_V_read_int_reg),
    .din1(grp_fu_846_p1),
    .ce(grp_fu_846_ce),
    .dout(grp_fu_846_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U43(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_27_V_read_int_reg),
    .din1(grp_fu_847_p1),
    .ce(grp_fu_847_ce),
    .dout(grp_fu_847_p2)
);

myproject_mul_16s_11ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_11ns_26_2_0_U44(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_53_V_read_int_reg),
    .din1(grp_fu_848_p1),
    .ce(grp_fu_848_ce),
    .dout(grp_fu_848_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U45(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_17_V_read_int_reg),
    .din1(grp_fu_849_p1),
    .ce(grp_fu_849_ce),
    .dout(grp_fu_849_p2)
);

myproject_mul_16s_11ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_11ns_26_2_0_U46(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_25_V_read_int_reg),
    .din1(grp_fu_850_p1),
    .ce(grp_fu_850_ce),
    .dout(grp_fu_850_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U47(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_43_V_read_int_reg),
    .din1(grp_fu_851_p1),
    .ce(grp_fu_851_ce),
    .dout(grp_fu_851_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U48(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_0_V_read_int_reg),
    .din1(grp_fu_852_p1),
    .ce(grp_fu_852_ce),
    .dout(grp_fu_852_p2)
);

myproject_mul_16s_11ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_11ns_26_2_0_U49(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_29_V_read_int_reg),
    .din1(grp_fu_853_p1),
    .ce(grp_fu_853_ce),
    .dout(grp_fu_853_p2)
);

myproject_mul_16s_13ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 13 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_13ns_26_2_0_U50(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_54_V_read_int_reg),
    .din1(grp_fu_854_p1),
    .ce(grp_fu_854_ce),
    .dout(grp_fu_854_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U51(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_45_V_read_int_reg),
    .din1(grp_fu_855_p1),
    .ce(grp_fu_855_ce),
    .dout(grp_fu_855_p2)
);

myproject_mul_16s_11ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_11ns_26_2_0_U52(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_11_V_read_int_reg),
    .din1(grp_fu_856_p1),
    .ce(grp_fu_856_ce),
    .dout(grp_fu_856_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U53(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_4_V_read_int_reg),
    .din1(grp_fu_857_p1),
    .ce(grp_fu_857_ce),
    .dout(grp_fu_857_p2)
);

myproject_mul_16s_11ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_11ns_26_2_0_U54(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_33_V_read_int_reg),
    .din1(grp_fu_858_p1),
    .ce(grp_fu_858_ce),
    .dout(grp_fu_858_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U55(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_10_V_read_int_reg),
    .din1(grp_fu_859_p1),
    .ce(grp_fu_859_ce),
    .dout(grp_fu_859_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U56(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_2_V_read_int_reg),
    .din1(grp_fu_860_p1),
    .ce(grp_fu_860_ce),
    .dout(grp_fu_860_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U57(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_48_V_read_int_reg),
    .din1(grp_fu_861_p1),
    .ce(grp_fu_861_ce),
    .dout(grp_fu_861_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U58(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_50_V_read_int_reg),
    .din1(grp_fu_862_p1),
    .ce(grp_fu_862_ce),
    .dout(grp_fu_862_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U59(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_51_V_read_int_reg),
    .din1(grp_fu_863_p1),
    .ce(grp_fu_863_ce),
    .dout(grp_fu_863_p2)
);

myproject_mul_16s_11ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 11 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_11ns_26_2_0_U60(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_57_V_read_int_reg),
    .din1(grp_fu_864_p1),
    .ce(grp_fu_864_ce),
    .dout(grp_fu_864_p2)
);

myproject_mul_16s_12ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 12 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_12ns_26_2_0_U61(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_7_V_read_int_reg),
    .din1(grp_fu_866_p1),
    .ce(grp_fu_866_ce),
    .dout(grp_fu_866_p2)
);

myproject_mul_16s_13ns_26_2_0 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 13 ),
    .dout_WIDTH( 26 ))
myproject_mul_16s_13ns_26_2_0_U62(
    .clk(ap_clk),
    .reset(ap_rst),
    .din0(data_40_V_read_int_reg),
    .din1(grp_fu_867_p1),
    .ce(grp_fu_867_ce),
    .dout(grp_fu_867_p2)
);

always @ (posedge ap_clk) begin
    ap_ce_reg <= ap_ce;
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_ce_reg)) begin
        ap_return_0_int_reg <= add_ln703_fu_17921_p2;
        ap_return_10_int_reg <= add_ln703_45_fu_17971_p2;
        ap_return_11_int_reg <= add_ln703_46_fu_17976_p2;
        ap_return_12_int_reg <= add_ln703_47_fu_17981_p2;
        ap_return_13_int_reg <= add_ln703_48_fu_17986_p2;
        ap_return_14_int_reg <= add_ln703_49_fu_17991_p2;
        ap_return_15_int_reg <= add_ln703_50_fu_17996_p2;
        ap_return_16_int_reg <= add_ln703_51_fu_18001_p2;
        ap_return_17_int_reg <= add_ln703_52_fu_18006_p2;
        ap_return_18_int_reg <= add_ln703_53_fu_18011_p2;
        ap_return_19_int_reg <= add_ln703_54_fu_18016_p2;
        ap_return_1_int_reg <= add_ln703_36_fu_17926_p2;
        ap_return_20_int_reg <= add_ln703_55_fu_18021_p2;
        ap_return_21_int_reg <= add_ln703_56_fu_18026_p2;
        ap_return_22_int_reg <= add_ln703_57_fu_18031_p2;
        ap_return_23_int_reg <= add_ln703_58_fu_18036_p2;
        ap_return_24_int_reg <= add_ln703_59_fu_18041_p2;
        ap_return_25_int_reg <= add_ln703_60_fu_18046_p2;
        ap_return_26_int_reg <= add_ln703_61_fu_18051_p2;
        ap_return_27_int_reg <= add_ln703_62_fu_18056_p2;
        ap_return_28_int_reg <= add_ln703_63_fu_18061_p2;
        ap_return_29_int_reg <= add_ln703_64_fu_18066_p2;
        ap_return_2_int_reg <= add_ln703_37_fu_17931_p2;
        ap_return_30_int_reg <= add_ln703_65_fu_18071_p2;
        ap_return_31_int_reg <= add_ln703_66_fu_18076_p2;
        ap_return_32_int_reg <= add_ln703_67_fu_18081_p2;
        ap_return_33_int_reg <= add_ln703_68_fu_18086_p2;
        ap_return_34_int_reg <= add_ln703_69_fu_18091_p2;
        ap_return_35_int_reg <= add_ln703_70_fu_18096_p2;
        ap_return_36_int_reg <= add_ln703_71_fu_18101_p2;
        ap_return_37_int_reg <= add_ln703_72_fu_18106_p2;
        ap_return_38_int_reg <= add_ln703_73_fu_18111_p2;
        ap_return_39_int_reg <= add_ln703_74_fu_18116_p2;
        ap_return_3_int_reg <= add_ln703_38_fu_17936_p2;
        ap_return_40_int_reg <= add_ln703_75_fu_18121_p2;
        ap_return_41_int_reg <= add_ln703_76_fu_18126_p2;
        ap_return_42_int_reg <= add_ln703_77_fu_18131_p2;
        ap_return_43_int_reg <= add_ln703_78_fu_18136_p2;
        ap_return_44_int_reg <= add_ln703_79_fu_18141_p2;
        ap_return_45_int_reg <= add_ln703_80_fu_18146_p2;
        ap_return_46_int_reg <= add_ln703_81_fu_18151_p2;
        ap_return_47_int_reg <= add_ln703_82_fu_18156_p2;
        ap_return_48_int_reg <= add_ln703_83_fu_18161_p2;
        ap_return_49_int_reg <= add_ln703_84_fu_18166_p2;
        ap_return_4_int_reg <= add_ln703_39_fu_17941_p2;
        ap_return_50_int_reg <= add_ln703_85_fu_18171_p2;
        ap_return_51_int_reg <= add_ln703_86_fu_18176_p2;
        ap_return_52_int_reg <= add_ln703_87_fu_18181_p2;
        ap_return_53_int_reg <= add_ln703_88_fu_18186_p2;
        ap_return_54_int_reg <= add_ln703_89_fu_18191_p2;
        ap_return_55_int_reg <= add_ln703_90_fu_18196_p2;
        ap_return_56_int_reg <= add_ln703_91_fu_18201_p2;
        ap_return_57_int_reg <= add_ln703_92_fu_18206_p2;
        ap_return_58_int_reg <= add_ln703_93_fu_18211_p2;
        ap_return_59_int_reg <= add_ln703_94_fu_18216_p2;
        ap_return_5_int_reg <= add_ln703_40_fu_17946_p2;
        ap_return_60_int_reg <= add_ln703_95_fu_18221_p2;
        ap_return_61_int_reg <= add_ln703_96_fu_18226_p2;
        ap_return_62_int_reg <= add_ln703_97_fu_18231_p2;
        ap_return_63_int_reg <= add_ln703_98_fu_18236_p2;
        ap_return_6_int_reg <= add_ln703_41_fu_17951_p2;
        ap_return_7_int_reg <= add_ln703_42_fu_17956_p2;
        ap_return_8_int_reg <= add_ln703_43_fu_17961_p2;
        ap_return_9_int_reg <= add_ln703_44_fu_17966_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_ce)) begin
        data_0_V_read_int_reg <= data_0_V_read;
        data_10_V_read_int_reg <= data_10_V_read;
        data_11_V_read_int_reg <= data_11_V_read;
        data_12_V_read_int_reg <= data_12_V_read;
        data_13_V_read_int_reg <= data_13_V_read;
        data_14_V_read_int_reg <= data_14_V_read;
        data_15_V_read_int_reg <= data_15_V_read;
        data_16_V_read_int_reg <= data_16_V_read;
        data_17_V_read_int_reg <= data_17_V_read;
        data_18_V_read_int_reg <= data_18_V_read;
        data_19_V_read_int_reg <= data_19_V_read;
        data_1_V_read_int_reg <= data_1_V_read;
        data_20_V_read_int_reg <= data_20_V_read;
        data_21_V_read_int_reg <= data_21_V_read;
        data_22_V_read_int_reg <= data_22_V_read;
        data_23_V_read_int_reg <= data_23_V_read;
        data_24_V_read_int_reg <= data_24_V_read;
        data_25_V_read_int_reg <= data_25_V_read;
        data_26_V_read_int_reg <= data_26_V_read;
        data_27_V_read_int_reg <= data_27_V_read;
        data_28_V_read_int_reg <= data_28_V_read;
        data_29_V_read_int_reg <= data_29_V_read;
        data_2_V_read_int_reg <= data_2_V_read;
        data_30_V_read_int_reg <= data_30_V_read;
        data_31_V_read_int_reg <= data_31_V_read;
        data_32_V_read_int_reg <= data_32_V_read;
        data_33_V_read_int_reg <= data_33_V_read;
        data_34_V_read_int_reg <= data_34_V_read;
        data_35_V_read_int_reg <= data_35_V_read;
        data_36_V_read_int_reg <= data_36_V_read;
        data_37_V_read_int_reg <= data_37_V_read;
        data_38_V_read_int_reg <= data_38_V_read;
        data_39_V_read_int_reg <= data_39_V_read;
        data_3_V_read_int_reg <= data_3_V_read;
        data_40_V_read_int_reg <= data_40_V_read;
        data_41_V_read_int_reg <= data_41_V_read;
        data_42_V_read_int_reg <= data_42_V_read;
        data_43_V_read_int_reg <= data_43_V_read;
        data_44_V_read_int_reg <= data_44_V_read;
        data_45_V_read_int_reg <= data_45_V_read;
        data_46_V_read_int_reg <= data_46_V_read;
        data_47_V_read_int_reg <= data_47_V_read;
        data_48_V_read_int_reg <= data_48_V_read;
        data_49_V_read_int_reg <= data_49_V_read;
        data_4_V_read_int_reg <= data_4_V_read;
        data_50_V_read_int_reg <= data_50_V_read;
        data_51_V_read_int_reg <= data_51_V_read;
        data_52_V_read_int_reg <= data_52_V_read;
        data_53_V_read_int_reg <= data_53_V_read;
        data_54_V_read_int_reg <= data_54_V_read;
        data_55_V_read_int_reg <= data_55_V_read;
        data_56_V_read_int_reg <= data_56_V_read;
        data_57_V_read_int_reg <= data_57_V_read;
        data_58_V_read_int_reg <= data_58_V_read;
        data_59_V_read_int_reg <= data_59_V_read;
        data_5_V_read_int_reg <= data_5_V_read;
        data_60_V_read_int_reg <= data_60_V_read;
        data_61_V_read_int_reg <= data_61_V_read;
        data_62_V_read_int_reg <= data_62_V_read;
        data_63_V_read_int_reg <= data_63_V_read;
        data_6_V_read_int_reg <= data_6_V_read;
        data_7_V_read_int_reg <= data_7_V_read;
        data_8_V_read_int_reg <= data_8_V_read;
        data_9_V_read_int_reg <= data_9_V_read;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        data_39_V_read_2_reg_18637 <= data_39_V_read_int_reg;
        data_42_V_read_2_reg_18631 <= data_42_V_read_int_reg;
        data_46_V_read_2_reg_18625 <= data_46_V_read_int_reg;
        trunc_ln708_31_reg_18953 <= {{grp_fu_832_p2[25:10]}};
        trunc_ln708_32_reg_18958 <= {{grp_fu_860_p2[25:10]}};
        trunc_ln708_33_reg_18968 <= {{grp_fu_857_p2[25:10]}};
        trunc_ln708_34_reg_18973 <= {{grp_fu_846_p2[25:10]}};
        trunc_ln708_35_reg_18978 <= {{grp_fu_829_p2[25:10]}};
        trunc_ln708_36_reg_18983 <= {{grp_fu_866_p2[25:10]}};
        trunc_ln708_37_reg_18988 <= {{grp_fu_819_p2[25:10]}};
        trunc_ln708_38_reg_18993 <= {{grp_fu_844_p2[25:10]}};
        trunc_ln708_39_reg_18998 <= {{grp_fu_859_p2[25:10]}};
        trunc_ln708_40_reg_19003 <= {{grp_fu_856_p2[25:10]}};
        trunc_ln708_41_reg_19008 <= {{grp_fu_834_p2[25:10]}};
        trunc_ln708_42_reg_19013 <= {{grp_fu_813_p2[25:10]}};
        trunc_ln708_43_reg_19018 <= {{grp_fu_816_p2[25:10]}};
        trunc_ln708_44_reg_19023 <= {{grp_fu_812_p2[25:10]}};
        trunc_ln708_45_reg_19028 <= {{grp_fu_837_p2[25:10]}};
        trunc_ln708_46_reg_19033 <= {{grp_fu_849_p2[25:10]}};
        trunc_ln708_47_reg_19038 <= {{grp_fu_818_p2[25:10]}};
        trunc_ln708_48_reg_19043 <= {{grp_fu_810_p2[25:10]}};
        trunc_ln708_49_reg_19048 <= {{grp_fu_815_p2[25:10]}};
        trunc_ln708_50_reg_19053 <= {{grp_fu_811_p2[25:10]}};
        trunc_ln708_51_reg_19058 <= {{grp_fu_824_p2[25:10]}};
        trunc_ln708_52_reg_19063 <= {{grp_fu_830_p2[25:10]}};
        trunc_ln708_53_reg_19068 <= {{grp_fu_839_p2[25:10]}};
        trunc_ln708_54_reg_19073 <= {{grp_fu_850_p2[25:10]}};
        trunc_ln708_55_reg_19078 <= {{grp_fu_827_p2[25:10]}};
        trunc_ln708_56_reg_19083 <= {{grp_fu_847_p2[25:10]}};
        trunc_ln708_57_reg_19088 <= {{grp_fu_845_p2[25:10]}};
        trunc_ln708_58_reg_19093 <= {{grp_fu_853_p2[25:10]}};
        trunc_ln708_59_reg_19098 <= {{grp_fu_814_p2[25:10]}};
        trunc_ln708_60_reg_19103 <= {{grp_fu_840_p2[25:10]}};
        trunc_ln708_61_reg_19108 <= {{grp_fu_808_p2[25:10]}};
        trunc_ln708_62_reg_19113 <= {{grp_fu_858_p2[25:10]}};
        trunc_ln708_63_reg_19118 <= {{grp_fu_835_p2[25:10]}};
        trunc_ln708_64_reg_19123 <= {{grp_fu_804_p2[25:10]}};
        trunc_ln708_65_reg_19128 <= {{grp_fu_841_p2[25:10]}};
        trunc_ln708_66_reg_19133 <= {{grp_fu_807_p2[25:10]}};
        trunc_ln708_67_reg_19138 <= {{grp_fu_825_p2[25:10]}};
        trunc_ln708_68_reg_19143 <= {{add_ln1118_fu_17625_p2[25:10]}};
        trunc_ln708_69_reg_19148 <= {{grp_fu_867_p2[25:10]}};
        trunc_ln708_70_reg_19153 <= {{grp_fu_822_p2[25:10]}};
        trunc_ln708_71_reg_19158 <= {{add_ln1118_1_fu_17671_p2[25:10]}};
        trunc_ln708_72_reg_19163 <= {{grp_fu_851_p2[25:10]}};
        trunc_ln708_73_reg_19168 <= {{grp_fu_826_p2[25:10]}};
        trunc_ln708_74_reg_19173 <= {{grp_fu_855_p2[25:10]}};
        trunc_ln708_75_reg_19178 <= {{add_ln1118_2_fu_17735_p2[25:10]}};
        trunc_ln708_76_reg_19183 <= {{grp_fu_838_p2[25:10]}};
        trunc_ln708_77_reg_19188 <= {{grp_fu_861_p2[25:10]}};
        trunc_ln708_78_reg_19193 <= {{grp_fu_843_p2[25:10]}};
        trunc_ln708_79_reg_19198 <= {{grp_fu_862_p2[25:10]}};
        trunc_ln708_80_reg_19203 <= {{grp_fu_863_p2[25:10]}};
        trunc_ln708_81_reg_19208 <= {{grp_fu_823_p2[25:10]}};
        trunc_ln708_82_reg_19213 <= {{grp_fu_848_p2[25:10]}};
        trunc_ln708_83_reg_19218 <= {{grp_fu_854_p2[25:10]}};
        trunc_ln708_84_reg_19223 <= {{grp_fu_821_p2[25:10]}};
        trunc_ln708_85_reg_19228 <= {{grp_fu_831_p2[25:10]}};
        trunc_ln708_86_reg_19233 <= {{grp_fu_864_p2[25:10]}};
        trunc_ln708_87_reg_19238 <= {{grp_fu_809_p2[25:10]}};
        trunc_ln708_88_reg_19243 <= {{grp_fu_842_p2[25:10]}};
        trunc_ln708_89_reg_19248 <= {{grp_fu_805_p2[25:10]}};
        trunc_ln708_90_reg_19253 <= {{grp_fu_833_p2[25:10]}};
        trunc_ln708_91_reg_19258 <= {{grp_fu_806_p2[25:10]}};
        trunc_ln708_92_reg_19263 <= {{grp_fu_820_p2[25:10]}};
        trunc_ln708_s_reg_18963 <= {{grp_fu_828_p2[25:10]}};
        trunc_ln_reg_18948 <= {{grp_fu_852_p2[25:10]}};
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_0 = ap_return_0_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_0 = add_ln703_fu_17921_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_1 = ap_return_1_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_1 = add_ln703_36_fu_17926_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_10 = ap_return_10_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_10 = add_ln703_45_fu_17971_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_11 = ap_return_11_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_11 = add_ln703_46_fu_17976_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_12 = ap_return_12_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_12 = add_ln703_47_fu_17981_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_13 = ap_return_13_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_13 = add_ln703_48_fu_17986_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_14 = ap_return_14_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_14 = add_ln703_49_fu_17991_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_15 = ap_return_15_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_15 = add_ln703_50_fu_17996_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_16 = ap_return_16_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_16 = add_ln703_51_fu_18001_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_17 = ap_return_17_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_17 = add_ln703_52_fu_18006_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_18 = ap_return_18_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_18 = add_ln703_53_fu_18011_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_19 = ap_return_19_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_19 = add_ln703_54_fu_18016_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_2 = ap_return_2_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_2 = add_ln703_37_fu_17931_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_20 = ap_return_20_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_20 = add_ln703_55_fu_18021_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_21 = ap_return_21_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_21 = add_ln703_56_fu_18026_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_22 = ap_return_22_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_22 = add_ln703_57_fu_18031_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_23 = ap_return_23_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_23 = add_ln703_58_fu_18036_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_24 = ap_return_24_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_24 = add_ln703_59_fu_18041_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_25 = ap_return_25_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_25 = add_ln703_60_fu_18046_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_26 = ap_return_26_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_26 = add_ln703_61_fu_18051_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_27 = ap_return_27_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_27 = add_ln703_62_fu_18056_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_28 = ap_return_28_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_28 = add_ln703_63_fu_18061_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_29 = ap_return_29_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_29 = add_ln703_64_fu_18066_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_3 = ap_return_3_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_3 = add_ln703_38_fu_17936_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_30 = ap_return_30_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_30 = add_ln703_65_fu_18071_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_31 = ap_return_31_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_31 = add_ln703_66_fu_18076_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_32 = ap_return_32_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_32 = add_ln703_67_fu_18081_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_33 = ap_return_33_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_33 = add_ln703_68_fu_18086_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_34 = ap_return_34_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_34 = add_ln703_69_fu_18091_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_35 = ap_return_35_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_35 = add_ln703_70_fu_18096_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_36 = ap_return_36_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_36 = add_ln703_71_fu_18101_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_37 = ap_return_37_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_37 = add_ln703_72_fu_18106_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_38 = ap_return_38_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_38 = add_ln703_73_fu_18111_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_39 = ap_return_39_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_39 = add_ln703_74_fu_18116_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_4 = ap_return_4_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_4 = add_ln703_39_fu_17941_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_40 = ap_return_40_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_40 = add_ln703_75_fu_18121_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_41 = ap_return_41_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_41 = add_ln703_76_fu_18126_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_42 = ap_return_42_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_42 = add_ln703_77_fu_18131_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_43 = ap_return_43_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_43 = add_ln703_78_fu_18136_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_44 = ap_return_44_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_44 = add_ln703_79_fu_18141_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_45 = ap_return_45_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_45 = add_ln703_80_fu_18146_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_46 = ap_return_46_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_46 = add_ln703_81_fu_18151_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_47 = ap_return_47_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_47 = add_ln703_82_fu_18156_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_48 = ap_return_48_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_48 = add_ln703_83_fu_18161_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_49 = ap_return_49_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_49 = add_ln703_84_fu_18166_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_5 = ap_return_5_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_5 = add_ln703_40_fu_17946_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_50 = ap_return_50_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_50 = add_ln703_85_fu_18171_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_51 = ap_return_51_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_51 = add_ln703_86_fu_18176_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_52 = ap_return_52_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_52 = add_ln703_87_fu_18181_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_53 = ap_return_53_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_53 = add_ln703_88_fu_18186_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_54 = ap_return_54_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_54 = add_ln703_89_fu_18191_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_55 = ap_return_55_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_55 = add_ln703_90_fu_18196_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_56 = ap_return_56_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_56 = add_ln703_91_fu_18201_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_57 = ap_return_57_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_57 = add_ln703_92_fu_18206_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_58 = ap_return_58_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_58 = add_ln703_93_fu_18211_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_59 = ap_return_59_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_59 = add_ln703_94_fu_18216_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_6 = ap_return_6_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_6 = add_ln703_41_fu_17951_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_60 = ap_return_60_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_60 = add_ln703_95_fu_18221_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_61 = ap_return_61_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_61 = add_ln703_96_fu_18226_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_62 = ap_return_62_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_62 = add_ln703_97_fu_18231_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_63 = ap_return_63_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_63 = add_ln703_98_fu_18236_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_7 = ap_return_7_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_7 = add_ln703_42_fu_17956_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_8 = ap_return_8_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_8 = add_ln703_43_fu_17961_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_9 = ap_return_9_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_9 = add_ln703_44_fu_17966_p2;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_804_ce = 1'b1;
    end else begin
        grp_fu_804_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_805_ce = 1'b1;
    end else begin
        grp_fu_805_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_806_ce = 1'b1;
    end else begin
        grp_fu_806_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_807_ce = 1'b1;
    end else begin
        grp_fu_807_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_808_ce = 1'b1;
    end else begin
        grp_fu_808_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_809_ce = 1'b1;
    end else begin
        grp_fu_809_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_810_ce = 1'b1;
    end else begin
        grp_fu_810_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_811_ce = 1'b1;
    end else begin
        grp_fu_811_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_812_ce = 1'b1;
    end else begin
        grp_fu_812_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_813_ce = 1'b1;
    end else begin
        grp_fu_813_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_814_ce = 1'b1;
    end else begin
        grp_fu_814_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_815_ce = 1'b1;
    end else begin
        grp_fu_815_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_816_ce = 1'b1;
    end else begin
        grp_fu_816_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_818_ce = 1'b1;
    end else begin
        grp_fu_818_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_819_ce = 1'b1;
    end else begin
        grp_fu_819_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_820_ce = 1'b1;
    end else begin
        grp_fu_820_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_821_ce = 1'b1;
    end else begin
        grp_fu_821_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_822_ce = 1'b1;
    end else begin
        grp_fu_822_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_823_ce = 1'b1;
    end else begin
        grp_fu_823_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_824_ce = 1'b1;
    end else begin
        grp_fu_824_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_825_ce = 1'b1;
    end else begin
        grp_fu_825_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_826_ce = 1'b1;
    end else begin
        grp_fu_826_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_827_ce = 1'b1;
    end else begin
        grp_fu_827_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_828_ce = 1'b1;
    end else begin
        grp_fu_828_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_829_ce = 1'b1;
    end else begin
        grp_fu_829_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_830_ce = 1'b1;
    end else begin
        grp_fu_830_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_831_ce = 1'b1;
    end else begin
        grp_fu_831_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_832_ce = 1'b1;
    end else begin
        grp_fu_832_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_833_ce = 1'b1;
    end else begin
        grp_fu_833_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_834_ce = 1'b1;
    end else begin
        grp_fu_834_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_835_ce = 1'b1;
    end else begin
        grp_fu_835_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_837_ce = 1'b1;
    end else begin
        grp_fu_837_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_838_ce = 1'b1;
    end else begin
        grp_fu_838_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_839_ce = 1'b1;
    end else begin
        grp_fu_839_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_840_ce = 1'b1;
    end else begin
        grp_fu_840_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_841_ce = 1'b1;
    end else begin
        grp_fu_841_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_842_ce = 1'b1;
    end else begin
        grp_fu_842_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_843_ce = 1'b1;
    end else begin
        grp_fu_843_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_844_ce = 1'b1;
    end else begin
        grp_fu_844_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_845_ce = 1'b1;
    end else begin
        grp_fu_845_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_846_ce = 1'b1;
    end else begin
        grp_fu_846_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_847_ce = 1'b1;
    end else begin
        grp_fu_847_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_848_ce = 1'b1;
    end else begin
        grp_fu_848_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_849_ce = 1'b1;
    end else begin
        grp_fu_849_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_850_ce = 1'b1;
    end else begin
        grp_fu_850_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_851_ce = 1'b1;
    end else begin
        grp_fu_851_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_852_ce = 1'b1;
    end else begin
        grp_fu_852_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_853_ce = 1'b1;
    end else begin
        grp_fu_853_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_854_ce = 1'b1;
    end else begin
        grp_fu_854_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_855_ce = 1'b1;
    end else begin
        grp_fu_855_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_856_ce = 1'b1;
    end else begin
        grp_fu_856_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_857_ce = 1'b1;
    end else begin
        grp_fu_857_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_858_ce = 1'b1;
    end else begin
        grp_fu_858_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_859_ce = 1'b1;
    end else begin
        grp_fu_859_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_860_ce = 1'b1;
    end else begin
        grp_fu_860_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_861_ce = 1'b1;
    end else begin
        grp_fu_861_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_862_ce = 1'b1;
    end else begin
        grp_fu_862_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_863_ce = 1'b1;
    end else begin
        grp_fu_863_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_864_ce = 1'b1;
    end else begin
        grp_fu_864_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_866_ce = 1'b1;
    end else begin
        grp_fu_866_ce = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        grp_fu_867_ce = 1'b1;
    end else begin
        grp_fu_867_ce = 1'b0;
    end
end

assign add_ln1118_1_fu_17671_p2 = ((sext_ln1118_76_fu_17661_p1) + (shl_ln1118_6_fu_17664_p3));

assign add_ln1118_2_fu_17735_p2 = ((shl_ln1118_7_fu_17717_p3) + (sext_ln1118_80_fu_17731_p1));

assign add_ln1118_fu_17625_p2 = ((shl_ln_fu_17607_p3) + (sext_ln1118_73_fu_17621_p1));

assign add_ln703_36_fu_17926_p2 = (trunc_ln708_31_reg_18953 + 16'd2428);

assign add_ln703_37_fu_17931_p2 = ((trunc_ln708_32_reg_18958) + (16'd63557));

assign add_ln703_38_fu_17936_p2 = (trunc_ln708_s_reg_18963 + 16'd2668);

assign add_ln703_39_fu_17941_p2 = (trunc_ln708_33_reg_18968 + 16'd770);

assign add_ln703_40_fu_17946_p2 = ((trunc_ln708_34_reg_18973) + (16'd65261));

assign add_ln703_41_fu_17951_p2 = (trunc_ln708_35_reg_18978 + 16'd1774);

assign add_ln703_42_fu_17956_p2 = ((trunc_ln708_36_reg_18983) + (16'd61620));

assign add_ln703_43_fu_17961_p2 = (trunc_ln708_37_reg_18988 + 16'd1134);

assign add_ln703_44_fu_17966_p2 = (trunc_ln708_38_reg_18993 + 16'd3344);

assign add_ln703_45_fu_17971_p2 = (trunc_ln708_39_reg_18998 + 16'd476);

assign add_ln703_46_fu_17976_p2 = ((trunc_ln708_40_reg_19003) + (16'd65055));

assign add_ln703_47_fu_17981_p2 = ((trunc_ln708_41_reg_19008) + (16'd63350));

assign add_ln703_48_fu_17986_p2 = (trunc_ln708_42_reg_19013 + 16'd6336);

assign add_ln703_49_fu_17991_p2 = (trunc_ln708_43_reg_19018 + 16'd779);

assign add_ln703_50_fu_17996_p2 = ((trunc_ln708_44_reg_19023) + (16'd65093));

assign add_ln703_51_fu_18001_p2 = ((trunc_ln708_45_reg_19028) + (16'd64452));

assign add_ln703_52_fu_18006_p2 = (trunc_ln708_46_reg_19033 + 16'd150);

assign add_ln703_53_fu_18011_p2 = ((trunc_ln708_47_reg_19038) + (16'd64356));

assign add_ln703_54_fu_18016_p2 = ((trunc_ln708_48_reg_19043) + (16'd61833));

assign add_ln703_55_fu_18021_p2 = ((trunc_ln708_49_reg_19048) + (16'd62693));

assign add_ln703_56_fu_18026_p2 = ((trunc_ln708_50_reg_19053) + (16'd65182));

assign add_ln703_57_fu_18031_p2 = ((trunc_ln708_51_reg_19058) + (16'd65467));

assign add_ln703_58_fu_18036_p2 = ((trunc_ln708_52_reg_19063) + (16'd65273));

assign add_ln703_59_fu_18041_p2 = ((trunc_ln708_53_reg_19068) + (16'd64093));

assign add_ln703_60_fu_18046_p2 = (trunc_ln708_54_reg_19073 + 16'd639);

assign add_ln703_61_fu_18051_p2 = ((trunc_ln708_55_reg_19078) + (16'd61811));

assign add_ln703_62_fu_18056_p2 = (trunc_ln708_56_reg_19083 + 16'd2997);

assign add_ln703_63_fu_18061_p2 = ((trunc_ln708_57_reg_19088) + (16'd65397));

assign add_ln703_64_fu_18066_p2 = ((trunc_ln708_58_reg_19093) + (16'd62604));

assign add_ln703_65_fu_18071_p2 = ((trunc_ln708_59_reg_19098) + (16'd60961));

assign add_ln703_66_fu_18076_p2 = (trunc_ln708_60_reg_19103 + 16'd3539);

assign add_ln703_67_fu_18081_p2 = ((trunc_ln708_61_reg_19108) + (16'd64305));

assign add_ln703_68_fu_18086_p2 = ((trunc_ln708_62_reg_19113) + (16'd64971));

assign add_ln703_69_fu_18091_p2 = (trunc_ln708_63_reg_19118 + 16'd427);

assign add_ln703_70_fu_18096_p2 = (trunc_ln708_64_reg_19123 + 16'd942);

assign add_ln703_71_fu_18101_p2 = ((trunc_ln708_65_reg_19128) + (16'd64448));

assign add_ln703_72_fu_18106_p2 = ((trunc_ln708_66_reg_19133) + (16'd61149));

assign add_ln703_73_fu_18111_p2 = ((trunc_ln708_67_reg_19138) + (16'd63555));

assign add_ln703_74_fu_18116_p2 = ((trunc_ln708_68_reg_19143) + (16'd64965));

assign add_ln703_75_fu_18121_p2 = ((trunc_ln708_69_reg_19148) + (16'd65184));

assign add_ln703_76_fu_18126_p2 = ((trunc_ln708_70_reg_19153) + (16'd65085));

assign add_ln703_77_fu_18131_p2 = ((trunc_ln708_71_reg_19158) + (16'd63019));

assign add_ln703_78_fu_18136_p2 = (trunc_ln708_72_reg_19163 + 16'd436);

assign add_ln703_79_fu_18141_p2 = ((trunc_ln708_73_reg_19168) + (16'd62012));

assign add_ln703_80_fu_18146_p2 = (trunc_ln708_74_reg_19173 + 16'd946);

assign add_ln703_81_fu_18151_p2 = ((trunc_ln708_75_reg_19178) + (16'd65281));

assign add_ln703_82_fu_18156_p2 = (trunc_ln708_76_reg_19183 + 16'd473);

assign add_ln703_83_fu_18161_p2 = ((trunc_ln708_77_reg_19188) + (16'd64458));

assign add_ln703_84_fu_18166_p2 = ((trunc_ln708_78_reg_19193) + (16'd65219));

assign add_ln703_85_fu_18171_p2 = (trunc_ln708_79_reg_19198 + 16'd1658);

assign add_ln703_86_fu_18176_p2 = (trunc_ln708_80_reg_19203 + 16'd2181);

assign add_ln703_87_fu_18181_p2 = (trunc_ln708_81_reg_19208 + 16'd1895);

assign add_ln703_88_fu_18186_p2 = (trunc_ln708_82_reg_19213 + 16'd792);

assign add_ln703_89_fu_18191_p2 = ((trunc_ln708_83_reg_19218) + (16'd62636));

assign add_ln703_90_fu_18196_p2 = (trunc_ln708_84_reg_19223 + 16'd1428);

assign add_ln703_91_fu_18201_p2 = ((trunc_ln708_85_reg_19228) + (16'd64938));

assign add_ln703_92_fu_18206_p2 = (trunc_ln708_86_reg_19233 + 16'd931);

assign add_ln703_93_fu_18211_p2 = ((trunc_ln708_87_reg_19238) + (16'd63398));

assign add_ln703_94_fu_18216_p2 = (trunc_ln708_88_reg_19243 + 16'd1118);

assign add_ln703_95_fu_18221_p2 = (trunc_ln708_89_reg_19248 + 16'd139);

assign add_ln703_96_fu_18226_p2 = (trunc_ln708_90_reg_19253 + 16'd1493);

assign add_ln703_97_fu_18231_p2 = (trunc_ln708_91_reg_19258 + 16'd396);

assign add_ln703_98_fu_18236_p2 = ((trunc_ln708_92_reg_19263) + (16'd61920));

assign add_ln703_fu_17921_p2 = ((trunc_ln_reg_18948) + (16'd64219));

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_state1_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign grp_fu_804_p1 = 26'd1206;

assign grp_fu_805_p1 = 26'd1155;

assign grp_fu_806_p1 = 26'd1317;

assign grp_fu_807_p1 = 26'd1776;

assign grp_fu_808_p1 = 26'd753;

assign grp_fu_809_p1 = 26'd689;

assign grp_fu_810_p1 = 26'd1209;

assign grp_fu_811_p1 = 26'd880;

assign grp_fu_812_p1 = 26'd1483;

assign grp_fu_813_p1 = 26'd2953;

assign grp_fu_814_p1 = 26'd1379;

assign grp_fu_815_p1 = 26'd1208;

assign grp_fu_816_p1 = 26'd1089;

assign grp_fu_818_p1 = 26'd1827;

assign grp_fu_819_p1 = 26'd811;

assign grp_fu_820_p1 = 26'd1718;

assign grp_fu_821_p1 = 26'd1103;

assign grp_fu_822_p1 = 26'd1465;

assign grp_fu_823_p1 = 26'd1094;

assign grp_fu_824_p1 = 26'd1816;

assign grp_fu_825_p1 = 26'd850;

assign grp_fu_826_p1 = 26'd1241;

assign grp_fu_827_p1 = 26'd1315;

assign grp_fu_828_p1 = 26'd929;

assign grp_fu_829_p1 = 26'd931;

assign grp_fu_830_p1 = 26'd1361;

assign grp_fu_831_p1 = 26'd793;

assign grp_fu_832_p1 = 26'd999;

assign grp_fu_833_p1 = 26'd1589;

assign grp_fu_834_p1 = 26'd667;

assign grp_fu_835_p1 = 26'd1731;

assign grp_fu_837_p1 = 26'd1192;

assign grp_fu_838_p1 = 26'd2114;

assign grp_fu_839_p1 = 26'd832;

assign grp_fu_840_p1 = 26'd1254;

assign grp_fu_841_p1 = 26'd998;

assign grp_fu_842_p1 = 26'd1583;

assign grp_fu_843_p1 = 26'd947;

assign grp_fu_844_p1 = 26'd882;

assign grp_fu_845_p1 = 26'd936;

assign grp_fu_846_p1 = 26'd1168;

assign grp_fu_847_p1 = 26'd1604;

assign grp_fu_848_p1 = 26'd991;

assign grp_fu_849_p1 = 26'd1117;

assign grp_fu_850_p1 = 26'd817;

assign grp_fu_851_p1 = 26'd1116;

assign grp_fu_852_p1 = 26'd1611;

assign grp_fu_853_p1 = 26'd773;

assign grp_fu_854_p1 = 26'd2327;

assign grp_fu_855_p1 = 26'd1031;

assign grp_fu_856_p1 = 26'd868;

assign grp_fu_857_p1 = 26'd1751;

assign grp_fu_858_p1 = 26'd669;

assign grp_fu_859_p1 = 26'd1054;

assign grp_fu_860_p1 = 26'd1055;

assign grp_fu_861_p1 = 26'd1256;

assign grp_fu_862_p1 = 26'd1713;

assign grp_fu_863_p1 = 26'd1267;

assign grp_fu_864_p1 = 26'd901;

assign grp_fu_866_p1 = 26'd1881;

assign grp_fu_867_p1 = 26'd2145;

assign sext_ln1118_73_fu_17621_p1 = (shl_ln1118_5_fu_17614_p3);

assign sext_ln1118_76_fu_17661_p1 = data_42_V_read_2_reg_18631;

assign sext_ln1118_80_fu_17731_p1 = (shl_ln1118_8_fu_17724_p3);

assign shl_ln1118_5_fu_17614_p3 = {{data_39_V_read_2_reg_18637}, {7'd0}};

assign shl_ln1118_6_fu_17664_p3 = {{data_42_V_read_2_reg_18631}, {10'd0}};

assign shl_ln1118_7_fu_17717_p3 = {{data_46_V_read_2_reg_18625}, {10'd0}};

assign shl_ln1118_8_fu_17724_p3 = {{data_46_V_read_2_reg_18625}, {6'd0}};

assign shl_ln_fu_17607_p3 = {{data_39_V_read_2_reg_18637}, {10'd0}};

endmodule //normalize_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1
module myproject_mul_16s_13ns_26_2_0(
    clk,
    reset,
    ce,
    din0,
    din1,
    dout);

parameter ID = 32'd1;
parameter NUM_STAGE = 32'd1;
parameter din0_WIDTH = 32'd1;
parameter din1_WIDTH = 32'd1;
parameter dout_WIDTH = 32'd1;
input clk;
input reset;
input ce;
input[din0_WIDTH - 1:0] din0;
input[din1_WIDTH - 1:0] din1;
output[dout_WIDTH - 1:0] dout;



myproject_mul_16s_13ns_26_2_0_MulnS_2 myproject_mul_16s_13ns_26_2_0_MulnS_2_U(
    .clk( clk ),
    .ce( ce ),
    .a( din0 ),
    .b( din1 ),
    .p( dout ));

endmodule
module myproject_mul_16s_13ns_26_2_0_MulnS_2(clk, ce, a, b, p);
input clk;
input ce;
input  [16 - 1 : 0] a;
input [13 - 1 : 0] b;
output[26 - 1 : 0] p;
reg  [26 - 1 : 0] p;
wire  [26 - 1 : 0] tmp_product;

assign tmp_product = (a) * ({1'b0, b});
always @ (posedge clk) begin
    if (ce) begin
        p <= tmp_product;
    end
end
endmodule
module myproject_mul_16s_12ns_26_2_0(
    clk,
    reset,
    ce,
    din0,
    din1,
    dout);

parameter ID = 32'd1;
parameter NUM_STAGE = 32'd1;
parameter din0_WIDTH = 32'd1;
parameter din1_WIDTH = 32'd1;
parameter dout_WIDTH = 32'd1;
input clk;
input reset;
input ce;
input[din0_WIDTH - 1:0] din0;
input[din1_WIDTH - 1:0] din1;
output[dout_WIDTH - 1:0] dout;



myproject_mul_16s_12ns_26_2_0_MulnS_0 myproject_mul_16s_12ns_26_2_0_MulnS_0_U(
    .clk( clk ),
    .ce( ce ),
    .a( din0 ),
    .b( din1 ),
    .p( dout ));

endmodule
module myproject_mul_16s_12ns_26_2_0_MulnS_0(clk, ce, a, b, p);
input clk;
input ce;
input  [16 - 1 : 0] a;
input [12 - 1 : 0] b;
output[26 - 1 : 0] p;
reg  [26 - 1 : 0] p;
wire  [26 - 1 : 0] tmp_product;

assign tmp_product = (a) * ({1'b0, b});
always @ (posedge clk) begin
    if (ce) begin
        p <= tmp_product;
    end
end
endmodule

module myproject_mul_16s_11ns_26_2_0(
    clk,
    reset,
    ce,
    din0,
    din1,
    dout);

parameter ID = 32'd1;
parameter NUM_STAGE = 32'd1;
parameter din0_WIDTH = 32'd1;
parameter din1_WIDTH = 32'd1;
parameter dout_WIDTH = 32'd1;
input clk;
input reset;
input ce;
input[din0_WIDTH - 1:0] din0;
input[din1_WIDTH - 1:0] din1;
output[dout_WIDTH - 1:0] dout;



myproject_mul_16s_11ns_26_2_0_MulnS_1 myproject_mul_16s_11ns_26_2_0_MulnS_1_U(
    .clk( clk ),
    .ce( ce ),
    .a( din0 ),
    .b( din1 ),
    .p( dout ));

endmodule
module myproject_mul_16s_11ns_26_2_0_MulnS_1(clk, ce, a, b, p);
input clk;
input ce;
input  [16 - 1 : 0] a;
input [11 - 1 : 0] b;
output[26 - 1 : 0] p;
reg  [26 - 1 : 0] p;
wire  [26 - 1 : 0] tmp_product;

assign tmp_product = (a) * ({1'b0, b});
always @ (posedge clk) begin
    if (ce) begin
        p <= tmp_product;
    end
end
endmodule



