
module relu_max_ap_fixed_ap_fixed_1_relu1_config5_s (
        ap_ready,
        data_0_V_read,
        data_1_V_read,
        data_2_V_read,
        data_3_V_read,
        data_4_V_read,
        data_5_V_read,
        data_6_V_read,
        data_7_V_read,
        data_8_V_read,
        data_9_V_read,
        data_10_V_read,
        data_11_V_read,
        data_12_V_read,
        data_13_V_read,
        data_14_V_read,
        data_15_V_read,
        data_16_V_read,
        data_17_V_read,
        data_18_V_read,
        data_19_V_read,
        data_20_V_read,
        data_21_V_read,
        data_22_V_read,
        data_23_V_read,
        data_24_V_read,
        data_25_V_read,
        data_26_V_read,
        data_27_V_read,
        data_28_V_read,
        data_29_V_read,
        data_30_V_read,
        data_31_V_read,
        data_32_V_read,
        data_33_V_read,
        data_34_V_read,
        data_35_V_read,
        data_36_V_read,
        data_37_V_read,
        data_38_V_read,
        data_39_V_read,
        data_40_V_read,
        data_41_V_read,
        data_42_V_read,
        data_43_V_read,
        data_44_V_read,
        data_45_V_read,
        data_46_V_read,
        data_47_V_read,
        data_48_V_read,
        data_49_V_read,
        data_50_V_read,
        data_51_V_read,
        data_52_V_read,
        data_53_V_read,
        data_54_V_read,
        data_55_V_read,
        data_56_V_read,
        data_57_V_read,
        data_58_V_read,
        data_59_V_read,
        data_60_V_read,
        data_61_V_read,
        data_62_V_read,
        data_63_V_read,
        ap_return_0,
        ap_return_1,
        ap_return_2,
        ap_return_3,
        ap_return_4,
        ap_return_5,
        ap_return_6,
        ap_return_7,
        ap_return_8,
        ap_return_9,
        ap_return_10,
        ap_return_11,
        ap_return_12,
        ap_return_13,
        ap_return_14,
        ap_return_15,
        ap_return_16,
        ap_return_17,
        ap_return_18,
        ap_return_19,
        ap_return_20,
        ap_return_21,
        ap_return_22,
        ap_return_23,
        ap_return_24,
        ap_return_25,
        ap_return_26,
        ap_return_27,
        ap_return_28,
        ap_return_29,
        ap_return_30,
        ap_return_31,
        ap_return_32,
        ap_return_33,
        ap_return_34,
        ap_return_35,
        ap_return_36,
        ap_return_37,
        ap_return_38,
        ap_return_39,
        ap_return_40,
        ap_return_41,
        ap_return_42,
        ap_return_43,
        ap_return_44,
        ap_return_45,
        ap_return_46,
        ap_return_47,
        ap_return_48,
        ap_return_49,
        ap_return_50,
        ap_return_51,
        ap_return_52,
        ap_return_53,
        ap_return_54,
        ap_return_55,
        ap_return_56,
        ap_return_57,
        ap_return_58,
        ap_return_59,
        ap_return_60,
        ap_return_61,
        ap_return_62,
        ap_return_63
);


output   ap_ready;
input  [15:0] data_0_V_read;
input  [15:0] data_1_V_read;
input  [15:0] data_2_V_read;
input  [15:0] data_3_V_read;
input  [15:0] data_4_V_read;
input  [15:0] data_5_V_read;
input  [15:0] data_6_V_read;
input  [15:0] data_7_V_read;
input  [15:0] data_8_V_read;
input  [15:0] data_9_V_read;
input  [15:0] data_10_V_read;
input  [15:0] data_11_V_read;
input  [15:0] data_12_V_read;
input  [15:0] data_13_V_read;
input  [15:0] data_14_V_read;
input  [15:0] data_15_V_read;
input  [15:0] data_16_V_read;
input  [15:0] data_17_V_read;
input  [15:0] data_18_V_read;
input  [15:0] data_19_V_read;
input  [15:0] data_20_V_read;
input  [15:0] data_21_V_read;
input  [15:0] data_22_V_read;
input  [15:0] data_23_V_read;
input  [15:0] data_24_V_read;
input  [15:0] data_25_V_read;
input  [15:0] data_26_V_read;
input  [15:0] data_27_V_read;
input  [15:0] data_28_V_read;
input  [15:0] data_29_V_read;
input  [15:0] data_30_V_read;
input  [15:0] data_31_V_read;
input  [15:0] data_32_V_read;
input  [15:0] data_33_V_read;
input  [15:0] data_34_V_read;
input  [15:0] data_35_V_read;
input  [15:0] data_36_V_read;
input  [15:0] data_37_V_read;
input  [15:0] data_38_V_read;
input  [15:0] data_39_V_read;
input  [15:0] data_40_V_read;
input  [15:0] data_41_V_read;
input  [15:0] data_42_V_read;
input  [15:0] data_43_V_read;
input  [15:0] data_44_V_read;
input  [15:0] data_45_V_read;
input  [15:0] data_46_V_read;
input  [15:0] data_47_V_read;
input  [15:0] data_48_V_read;
input  [15:0] data_49_V_read;
input  [15:0] data_50_V_read;
input  [15:0] data_51_V_read;
input  [15:0] data_52_V_read;
input  [15:0] data_53_V_read;
input  [15:0] data_54_V_read;
input  [15:0] data_55_V_read;
input  [15:0] data_56_V_read;
input  [15:0] data_57_V_read;
input  [15:0] data_58_V_read;
input  [15:0] data_59_V_read;
input  [15:0] data_60_V_read;
input  [15:0] data_61_V_read;
input  [15:0] data_62_V_read;
input  [15:0] data_63_V_read;
output  [15:0] ap_return_0;
output  [15:0] ap_return_1;
output  [15:0] ap_return_2;
output  [15:0] ap_return_3;
output  [15:0] ap_return_4;
output  [15:0] ap_return_5;
output  [15:0] ap_return_6;
output  [15:0] ap_return_7;
output  [15:0] ap_return_8;
output  [15:0] ap_return_9;
output  [15:0] ap_return_10;
output  [15:0] ap_return_11;
output  [15:0] ap_return_12;
output  [15:0] ap_return_13;
output  [15:0] ap_return_14;
output  [15:0] ap_return_15;
output  [15:0] ap_return_16;
output  [15:0] ap_return_17;
output  [15:0] ap_return_18;
output  [15:0] ap_return_19;
output  [15:0] ap_return_20;
output  [15:0] ap_return_21;
output  [15:0] ap_return_22;
output  [15:0] ap_return_23;
output  [15:0] ap_return_24;
output  [15:0] ap_return_25;
output  [15:0] ap_return_26;
output  [15:0] ap_return_27;
output  [15:0] ap_return_28;
output  [15:0] ap_return_29;
output  [15:0] ap_return_30;
output  [15:0] ap_return_31;
output  [15:0] ap_return_32;
output  [15:0] ap_return_33;
output  [15:0] ap_return_34;
output  [15:0] ap_return_35;
output  [15:0] ap_return_36;
output  [15:0] ap_return_37;
output  [15:0] ap_return_38;
output  [15:0] ap_return_39;
output  [15:0] ap_return_40;
output  [15:0] ap_return_41;
output  [15:0] ap_return_42;
output  [15:0] ap_return_43;
output  [15:0] ap_return_44;
output  [15:0] ap_return_45;
output  [15:0] ap_return_46;
output  [15:0] ap_return_47;
output  [15:0] ap_return_48;
output  [15:0] ap_return_49;
output  [15:0] ap_return_50;
output  [15:0] ap_return_51;
output  [15:0] ap_return_52;
output  [15:0] ap_return_53;
output  [15:0] ap_return_54;
output  [15:0] ap_return_55;
output  [15:0] ap_return_56;
output  [15:0] ap_return_57;
output  [15:0] ap_return_58;
output  [15:0] ap_return_59;
output  [15:0] ap_return_60;
output  [15:0] ap_return_61;
output  [15:0] ap_return_62;
output  [15:0] ap_return_63;

wire   [0:0] tmp_98_fu_558_p3;
wire   [0:0] xor_ln1495_fu_566_p2;
wire   [10:0] tmp_99_fu_572_p3;
wire   [0:0] tmp_97_fu_544_p3;
wire   [0:0] icmp_ln1494_fu_552_p2;
wire   [0:0] or_ln1495_fu_584_p2;
wire   [15:0] zext_ln1495_fu_580_p1;
wire   [0:0] tmp_101_fu_612_p3;
wire   [0:0] xor_ln1495_32_fu_620_p2;
wire   [10:0] tmp_102_fu_626_p3;
wire   [0:0] tmp_100_fu_598_p3;
wire   [0:0] icmp_ln1494_1_fu_606_p2;
wire   [0:0] or_ln1495_32_fu_638_p2;
wire   [15:0] zext_ln1495_32_fu_634_p1;
wire   [0:0] tmp_104_fu_666_p3;
wire   [0:0] xor_ln1495_33_fu_674_p2;
wire   [10:0] tmp_105_fu_680_p3;
wire   [0:0] tmp_103_fu_652_p3;
wire   [0:0] icmp_ln1494_2_fu_660_p2;
wire   [0:0] or_ln1495_33_fu_692_p2;
wire   [15:0] zext_ln1495_33_fu_688_p1;
wire   [0:0] tmp_107_fu_720_p3;
wire   [0:0] xor_ln1495_34_fu_728_p2;
wire   [10:0] tmp_108_fu_734_p3;
wire   [0:0] tmp_106_fu_706_p3;
wire   [0:0] icmp_ln1494_3_fu_714_p2;
wire   [0:0] or_ln1495_34_fu_746_p2;
wire   [15:0] zext_ln1495_34_fu_742_p1;
wire   [0:0] tmp_110_fu_774_p3;
wire   [0:0] xor_ln1495_35_fu_782_p2;
wire   [10:0] tmp_111_fu_788_p3;
wire   [0:0] tmp_109_fu_760_p3;
wire   [0:0] icmp_ln1494_4_fu_768_p2;
wire   [0:0] or_ln1495_35_fu_800_p2;
wire   [15:0] zext_ln1495_35_fu_796_p1;
wire   [0:0] tmp_113_fu_828_p3;
wire   [0:0] xor_ln1495_36_fu_836_p2;
wire   [10:0] tmp_114_fu_842_p3;
wire   [0:0] tmp_112_fu_814_p3;
wire   [0:0] icmp_ln1494_5_fu_822_p2;
wire   [0:0] or_ln1495_36_fu_854_p2;
wire   [15:0] zext_ln1495_36_fu_850_p1;
wire   [0:0] tmp_116_fu_882_p3;
wire   [0:0] xor_ln1495_37_fu_890_p2;
wire   [10:0] tmp_117_fu_896_p3;
wire   [0:0] tmp_115_fu_868_p3;
wire   [0:0] icmp_ln1494_6_fu_876_p2;
wire   [0:0] or_ln1495_37_fu_908_p2;
wire   [15:0] zext_ln1495_37_fu_904_p1;
wire   [0:0] tmp_119_fu_936_p3;
wire   [0:0] xor_ln1495_38_fu_944_p2;
wire   [10:0] tmp_120_fu_950_p3;
wire   [0:0] tmp_118_fu_922_p3;
wire   [0:0] icmp_ln1494_7_fu_930_p2;
wire   [0:0] or_ln1495_38_fu_962_p2;
wire   [15:0] zext_ln1495_38_fu_958_p1;
wire   [0:0] tmp_122_fu_990_p3;
wire   [0:0] xor_ln1495_39_fu_998_p2;
wire   [10:0] tmp_123_fu_1004_p3;
wire   [0:0] tmp_121_fu_976_p3;
wire   [0:0] icmp_ln1494_8_fu_984_p2;
wire   [0:0] or_ln1495_39_fu_1016_p2;
wire   [15:0] zext_ln1495_39_fu_1012_p1;
wire   [0:0] tmp_125_fu_1044_p3;
wire   [0:0] xor_ln1495_40_fu_1052_p2;
wire   [10:0] tmp_126_fu_1058_p3;
wire   [0:0] tmp_124_fu_1030_p3;
wire   [0:0] icmp_ln1494_9_fu_1038_p2;
wire   [0:0] or_ln1495_40_fu_1070_p2;
wire   [15:0] zext_ln1495_40_fu_1066_p1;
wire   [0:0] tmp_128_fu_1098_p3;
wire   [0:0] xor_ln1495_41_fu_1106_p2;
wire   [10:0] tmp_129_fu_1112_p3;
wire   [0:0] tmp_127_fu_1084_p3;
wire   [0:0] icmp_ln1494_10_fu_1092_p2;
wire   [0:0] or_ln1495_41_fu_1124_p2;
wire   [15:0] zext_ln1495_41_fu_1120_p1;
wire   [0:0] tmp_131_fu_1152_p3;
wire   [0:0] xor_ln1495_42_fu_1160_p2;
wire   [10:0] tmp_132_fu_1166_p3;
wire   [0:0] tmp_130_fu_1138_p3;
wire   [0:0] icmp_ln1494_11_fu_1146_p2;
wire   [0:0] or_ln1495_42_fu_1178_p2;
wire   [15:0] zext_ln1495_42_fu_1174_p1;
wire   [0:0] tmp_134_fu_1206_p3;
wire   [0:0] xor_ln1495_43_fu_1214_p2;
wire   [10:0] tmp_135_fu_1220_p3;
wire   [0:0] tmp_133_fu_1192_p3;
wire   [0:0] icmp_ln1494_12_fu_1200_p2;
wire   [0:0] or_ln1495_43_fu_1232_p2;
wire   [15:0] zext_ln1495_43_fu_1228_p1;
wire   [0:0] tmp_137_fu_1260_p3;
wire   [0:0] xor_ln1495_44_fu_1268_p2;
wire   [10:0] tmp_138_fu_1274_p3;
wire   [0:0] tmp_136_fu_1246_p3;
wire   [0:0] icmp_ln1494_13_fu_1254_p2;
wire   [0:0] or_ln1495_44_fu_1286_p2;
wire   [15:0] zext_ln1495_44_fu_1282_p1;
wire   [0:0] tmp_140_fu_1314_p3;
wire   [0:0] xor_ln1495_45_fu_1322_p2;
wire   [10:0] tmp_141_fu_1328_p3;
wire   [0:0] tmp_139_fu_1300_p3;
wire   [0:0] icmp_ln1494_14_fu_1308_p2;
wire   [0:0] or_ln1495_45_fu_1340_p2;
wire   [15:0] zext_ln1495_45_fu_1336_p1;
wire   [0:0] tmp_143_fu_1368_p3;
wire   [0:0] xor_ln1495_46_fu_1376_p2;
wire   [10:0] tmp_144_fu_1382_p3;
wire   [0:0] tmp_142_fu_1354_p3;
wire   [0:0] icmp_ln1494_15_fu_1362_p2;
wire   [0:0] or_ln1495_46_fu_1394_p2;
wire   [15:0] zext_ln1495_46_fu_1390_p1;
wire   [0:0] tmp_146_fu_1422_p3;
wire   [0:0] xor_ln1495_47_fu_1430_p2;
wire   [10:0] tmp_147_fu_1436_p3;
wire   [0:0] tmp_145_fu_1408_p3;
wire   [0:0] icmp_ln1494_16_fu_1416_p2;
wire   [0:0] or_ln1495_47_fu_1448_p2;
wire   [15:0] zext_ln1495_47_fu_1444_p1;
wire   [0:0] tmp_149_fu_1476_p3;
wire   [0:0] xor_ln1495_48_fu_1484_p2;
wire   [10:0] tmp_150_fu_1490_p3;
wire   [0:0] tmp_148_fu_1462_p3;
wire   [0:0] icmp_ln1494_17_fu_1470_p2;
wire   [0:0] or_ln1495_48_fu_1502_p2;
wire   [15:0] zext_ln1495_48_fu_1498_p1;
wire   [0:0] tmp_152_fu_1530_p3;
wire   [0:0] xor_ln1495_49_fu_1538_p2;
wire   [10:0] tmp_153_fu_1544_p3;
wire   [0:0] tmp_151_fu_1516_p3;
wire   [0:0] icmp_ln1494_18_fu_1524_p2;
wire   [0:0] or_ln1495_49_fu_1556_p2;
wire   [15:0] zext_ln1495_49_fu_1552_p1;
wire   [0:0] tmp_155_fu_1584_p3;
wire   [0:0] xor_ln1495_50_fu_1592_p2;
wire   [10:0] tmp_156_fu_1598_p3;
wire   [0:0] tmp_154_fu_1570_p3;
wire   [0:0] icmp_ln1494_19_fu_1578_p2;
wire   [0:0] or_ln1495_50_fu_1610_p2;
wire   [15:0] zext_ln1495_50_fu_1606_p1;
wire   [0:0] tmp_158_fu_1638_p3;
wire   [0:0] xor_ln1495_51_fu_1646_p2;
wire   [10:0] tmp_159_fu_1652_p3;
wire   [0:0] tmp_157_fu_1624_p3;
wire   [0:0] icmp_ln1494_20_fu_1632_p2;
wire   [0:0] or_ln1495_51_fu_1664_p2;
wire   [15:0] zext_ln1495_51_fu_1660_p1;
wire   [0:0] tmp_161_fu_1692_p3;
wire   [0:0] xor_ln1495_52_fu_1700_p2;
wire   [10:0] tmp_162_fu_1706_p3;
wire   [0:0] tmp_160_fu_1678_p3;
wire   [0:0] icmp_ln1494_21_fu_1686_p2;
wire   [0:0] or_ln1495_52_fu_1718_p2;
wire   [15:0] zext_ln1495_52_fu_1714_p1;
wire   [0:0] tmp_164_fu_1746_p3;
wire   [0:0] xor_ln1495_53_fu_1754_p2;
wire   [10:0] tmp_165_fu_1760_p3;
wire   [0:0] tmp_163_fu_1732_p3;
wire   [0:0] icmp_ln1494_22_fu_1740_p2;
wire   [0:0] or_ln1495_53_fu_1772_p2;
wire   [15:0] zext_ln1495_53_fu_1768_p1;
wire   [0:0] tmp_167_fu_1800_p3;
wire   [0:0] xor_ln1495_54_fu_1808_p2;
wire   [10:0] tmp_168_fu_1814_p3;
wire   [0:0] tmp_166_fu_1786_p3;
wire   [0:0] icmp_ln1494_23_fu_1794_p2;
wire   [0:0] or_ln1495_54_fu_1826_p2;
wire   [15:0] zext_ln1495_54_fu_1822_p1;
wire   [0:0] tmp_170_fu_1854_p3;
wire   [0:0] xor_ln1495_55_fu_1862_p2;
wire   [10:0] tmp_171_fu_1868_p3;
wire   [0:0] tmp_169_fu_1840_p3;
wire   [0:0] icmp_ln1494_24_fu_1848_p2;
wire   [0:0] or_ln1495_55_fu_1880_p2;
wire   [15:0] zext_ln1495_55_fu_1876_p1;
wire   [0:0] tmp_173_fu_1908_p3;
wire   [0:0] xor_ln1495_56_fu_1916_p2;
wire   [10:0] tmp_174_fu_1922_p3;
wire   [0:0] tmp_172_fu_1894_p3;
wire   [0:0] icmp_ln1494_25_fu_1902_p2;
wire   [0:0] or_ln1495_56_fu_1934_p2;
wire   [15:0] zext_ln1495_56_fu_1930_p1;
wire   [0:0] tmp_176_fu_1962_p3;
wire   [0:0] xor_ln1495_57_fu_1970_p2;
wire   [10:0] tmp_177_fu_1976_p3;
wire   [0:0] tmp_175_fu_1948_p3;
wire   [0:0] icmp_ln1494_26_fu_1956_p2;
wire   [0:0] or_ln1495_57_fu_1988_p2;
wire   [15:0] zext_ln1495_57_fu_1984_p1;
wire   [0:0] tmp_179_fu_2016_p3;
wire   [0:0] xor_ln1495_58_fu_2024_p2;
wire   [10:0] tmp_180_fu_2030_p3;
wire   [0:0] tmp_178_fu_2002_p3;
wire   [0:0] icmp_ln1494_27_fu_2010_p2;
wire   [0:0] or_ln1495_58_fu_2042_p2;
wire   [15:0] zext_ln1495_58_fu_2038_p1;
wire   [0:0] tmp_182_fu_2070_p3;
wire   [0:0] xor_ln1495_59_fu_2078_p2;
wire   [10:0] tmp_183_fu_2084_p3;
wire   [0:0] tmp_181_fu_2056_p3;
wire   [0:0] icmp_ln1494_28_fu_2064_p2;
wire   [0:0] or_ln1495_59_fu_2096_p2;
wire   [15:0] zext_ln1495_59_fu_2092_p1;
wire   [0:0] tmp_185_fu_2124_p3;
wire   [0:0] xor_ln1495_60_fu_2132_p2;
wire   [10:0] tmp_186_fu_2138_p3;
wire   [0:0] tmp_184_fu_2110_p3;
wire   [0:0] icmp_ln1494_29_fu_2118_p2;
wire   [0:0] or_ln1495_60_fu_2150_p2;
wire   [15:0] zext_ln1495_60_fu_2146_p1;
wire   [0:0] tmp_188_fu_2178_p3;
wire   [0:0] xor_ln1495_61_fu_2186_p2;
wire   [10:0] tmp_189_fu_2192_p3;
wire   [0:0] tmp_187_fu_2164_p3;
wire   [0:0] icmp_ln1494_30_fu_2172_p2;
wire   [0:0] or_ln1495_61_fu_2204_p2;
wire   [15:0] zext_ln1495_61_fu_2200_p1;
wire   [0:0] tmp_191_fu_2232_p3;
wire   [0:0] xor_ln1495_62_fu_2240_p2;
wire   [10:0] tmp_192_fu_2246_p3;
wire   [0:0] tmp_190_fu_2218_p3;
wire   [0:0] icmp_ln1494_31_fu_2226_p2;
wire   [0:0] or_ln1495_62_fu_2258_p2;
wire   [15:0] zext_ln1495_62_fu_2254_p1;
wire   [0:0] tmp_194_fu_2286_p3;
wire   [0:0] xor_ln1495_63_fu_2294_p2;
wire   [10:0] tmp_195_fu_2300_p3;
wire   [0:0] tmp_193_fu_2272_p3;
wire   [0:0] icmp_ln1494_32_fu_2280_p2;
wire   [0:0] or_ln1495_63_fu_2312_p2;
wire   [15:0] zext_ln1495_63_fu_2308_p1;
wire   [0:0] tmp_197_fu_2340_p3;
wire   [0:0] xor_ln1495_64_fu_2348_p2;
wire   [10:0] tmp_198_fu_2354_p3;
wire   [0:0] tmp_196_fu_2326_p3;
wire   [0:0] icmp_ln1494_33_fu_2334_p2;
wire   [0:0] or_ln1495_64_fu_2366_p2;
wire   [15:0] zext_ln1495_64_fu_2362_p1;
wire   [0:0] tmp_200_fu_2394_p3;
wire   [0:0] xor_ln1495_65_fu_2402_p2;
wire   [10:0] tmp_201_fu_2408_p3;
wire   [0:0] tmp_199_fu_2380_p3;
wire   [0:0] icmp_ln1494_34_fu_2388_p2;
wire   [0:0] or_ln1495_65_fu_2420_p2;
wire   [15:0] zext_ln1495_65_fu_2416_p1;
wire   [0:0] tmp_203_fu_2448_p3;
wire   [0:0] xor_ln1495_66_fu_2456_p2;
wire   [10:0] tmp_204_fu_2462_p3;
wire   [0:0] tmp_202_fu_2434_p3;
wire   [0:0] icmp_ln1494_35_fu_2442_p2;
wire   [0:0] or_ln1495_66_fu_2474_p2;
wire   [15:0] zext_ln1495_66_fu_2470_p1;
wire   [0:0] tmp_206_fu_2502_p3;
wire   [0:0] xor_ln1495_67_fu_2510_p2;
wire   [10:0] tmp_207_fu_2516_p3;
wire   [0:0] tmp_205_fu_2488_p3;
wire   [0:0] icmp_ln1494_36_fu_2496_p2;
wire   [0:0] or_ln1495_67_fu_2528_p2;
wire   [15:0] zext_ln1495_67_fu_2524_p1;
wire   [0:0] tmp_209_fu_2556_p3;
wire   [0:0] xor_ln1495_68_fu_2564_p2;
wire   [10:0] tmp_210_fu_2570_p3;
wire   [0:0] tmp_208_fu_2542_p3;
wire   [0:0] icmp_ln1494_37_fu_2550_p2;
wire   [0:0] or_ln1495_68_fu_2582_p2;
wire   [15:0] zext_ln1495_68_fu_2578_p1;
wire   [0:0] tmp_212_fu_2610_p3;
wire   [0:0] xor_ln1495_69_fu_2618_p2;
wire   [10:0] tmp_213_fu_2624_p3;
wire   [0:0] tmp_211_fu_2596_p3;
wire   [0:0] icmp_ln1494_38_fu_2604_p2;
wire   [0:0] or_ln1495_69_fu_2636_p2;
wire   [15:0] zext_ln1495_69_fu_2632_p1;
wire   [0:0] tmp_215_fu_2664_p3;
wire   [0:0] xor_ln1495_70_fu_2672_p2;
wire   [10:0] tmp_216_fu_2678_p3;
wire   [0:0] tmp_214_fu_2650_p3;
wire   [0:0] icmp_ln1494_39_fu_2658_p2;
wire   [0:0] or_ln1495_70_fu_2690_p2;
wire   [15:0] zext_ln1495_70_fu_2686_p1;
wire   [0:0] tmp_218_fu_2718_p3;
wire   [0:0] xor_ln1495_71_fu_2726_p2;
wire   [10:0] tmp_219_fu_2732_p3;
wire   [0:0] tmp_217_fu_2704_p3;
wire   [0:0] icmp_ln1494_40_fu_2712_p2;
wire   [0:0] or_ln1495_71_fu_2744_p2;
wire   [15:0] zext_ln1495_71_fu_2740_p1;
wire   [0:0] tmp_221_fu_2772_p3;
wire   [0:0] xor_ln1495_72_fu_2780_p2;
wire   [10:0] tmp_222_fu_2786_p3;
wire   [0:0] tmp_220_fu_2758_p3;
wire   [0:0] icmp_ln1494_41_fu_2766_p2;
wire   [0:0] or_ln1495_72_fu_2798_p2;
wire   [15:0] zext_ln1495_72_fu_2794_p1;
wire   [0:0] tmp_224_fu_2826_p3;
wire   [0:0] xor_ln1495_73_fu_2834_p2;
wire   [10:0] tmp_225_fu_2840_p3;
wire   [0:0] tmp_223_fu_2812_p3;
wire   [0:0] icmp_ln1494_42_fu_2820_p2;
wire   [0:0] or_ln1495_73_fu_2852_p2;
wire   [15:0] zext_ln1495_73_fu_2848_p1;
wire   [0:0] tmp_227_fu_2880_p3;
wire   [0:0] xor_ln1495_74_fu_2888_p2;
wire   [10:0] tmp_228_fu_2894_p3;
wire   [0:0] tmp_226_fu_2866_p3;
wire   [0:0] icmp_ln1494_43_fu_2874_p2;
wire   [0:0] or_ln1495_74_fu_2906_p2;
wire   [15:0] zext_ln1495_74_fu_2902_p1;
wire   [0:0] tmp_230_fu_2934_p3;
wire   [0:0] xor_ln1495_75_fu_2942_p2;
wire   [10:0] tmp_231_fu_2948_p3;
wire   [0:0] tmp_229_fu_2920_p3;
wire   [0:0] icmp_ln1494_44_fu_2928_p2;
wire   [0:0] or_ln1495_75_fu_2960_p2;
wire   [15:0] zext_ln1495_75_fu_2956_p1;
wire   [0:0] tmp_233_fu_2988_p3;
wire   [0:0] xor_ln1495_76_fu_2996_p2;
wire   [10:0] tmp_234_fu_3002_p3;
wire   [0:0] tmp_232_fu_2974_p3;
wire   [0:0] icmp_ln1494_45_fu_2982_p2;
wire   [0:0] or_ln1495_76_fu_3014_p2;
wire   [15:0] zext_ln1495_76_fu_3010_p1;
wire   [0:0] tmp_236_fu_3042_p3;
wire   [0:0] xor_ln1495_77_fu_3050_p2;
wire   [10:0] tmp_237_fu_3056_p3;
wire   [0:0] tmp_235_fu_3028_p3;
wire   [0:0] icmp_ln1494_46_fu_3036_p2;
wire   [0:0] or_ln1495_77_fu_3068_p2;
wire   [15:0] zext_ln1495_77_fu_3064_p1;
wire   [0:0] tmp_239_fu_3096_p3;
wire   [0:0] xor_ln1495_78_fu_3104_p2;
wire   [10:0] tmp_240_fu_3110_p3;
wire   [0:0] tmp_238_fu_3082_p3;
wire   [0:0] icmp_ln1494_47_fu_3090_p2;
wire   [0:0] or_ln1495_78_fu_3122_p2;
wire   [15:0] zext_ln1495_78_fu_3118_p1;
wire   [0:0] tmp_242_fu_3150_p3;
wire   [0:0] xor_ln1495_79_fu_3158_p2;
wire   [10:0] tmp_243_fu_3164_p3;
wire   [0:0] tmp_241_fu_3136_p3;
wire   [0:0] icmp_ln1494_48_fu_3144_p2;
wire   [0:0] or_ln1495_79_fu_3176_p2;
wire   [15:0] zext_ln1495_79_fu_3172_p1;
wire   [0:0] tmp_245_fu_3204_p3;
wire   [0:0] xor_ln1495_80_fu_3212_p2;
wire   [10:0] tmp_246_fu_3218_p3;
wire   [0:0] tmp_244_fu_3190_p3;
wire   [0:0] icmp_ln1494_49_fu_3198_p2;
wire   [0:0] or_ln1495_80_fu_3230_p2;
wire   [15:0] zext_ln1495_80_fu_3226_p1;
wire   [0:0] tmp_248_fu_3258_p3;
wire   [0:0] xor_ln1495_81_fu_3266_p2;
wire   [10:0] tmp_249_fu_3272_p3;
wire   [0:0] tmp_247_fu_3244_p3;
wire   [0:0] icmp_ln1494_50_fu_3252_p2;
wire   [0:0] or_ln1495_81_fu_3284_p2;
wire   [15:0] zext_ln1495_81_fu_3280_p1;
wire   [0:0] tmp_251_fu_3312_p3;
wire   [0:0] xor_ln1495_82_fu_3320_p2;
wire   [10:0] tmp_252_fu_3326_p3;
wire   [0:0] tmp_250_fu_3298_p3;
wire   [0:0] icmp_ln1494_51_fu_3306_p2;
wire   [0:0] or_ln1495_82_fu_3338_p2;
wire   [15:0] zext_ln1495_82_fu_3334_p1;
wire   [0:0] tmp_254_fu_3366_p3;
wire   [0:0] xor_ln1495_83_fu_3374_p2;
wire   [10:0] tmp_255_fu_3380_p3;
wire   [0:0] tmp_253_fu_3352_p3;
wire   [0:0] icmp_ln1494_52_fu_3360_p2;
wire   [0:0] or_ln1495_83_fu_3392_p2;
wire   [15:0] zext_ln1495_83_fu_3388_p1;
wire   [0:0] tmp_257_fu_3420_p3;
wire   [0:0] xor_ln1495_84_fu_3428_p2;
wire   [10:0] tmp_258_fu_3434_p3;
wire   [0:0] tmp_256_fu_3406_p3;
wire   [0:0] icmp_ln1494_53_fu_3414_p2;
wire   [0:0] or_ln1495_84_fu_3446_p2;
wire   [15:0] zext_ln1495_84_fu_3442_p1;
wire   [0:0] tmp_260_fu_3474_p3;
wire   [0:0] xor_ln1495_85_fu_3482_p2;
wire   [10:0] tmp_261_fu_3488_p3;
wire   [0:0] tmp_259_fu_3460_p3;
wire   [0:0] icmp_ln1494_54_fu_3468_p2;
wire   [0:0] or_ln1495_85_fu_3500_p2;
wire   [15:0] zext_ln1495_85_fu_3496_p1;
wire   [0:0] tmp_263_fu_3528_p3;
wire   [0:0] xor_ln1495_86_fu_3536_p2;
wire   [10:0] tmp_264_fu_3542_p3;
wire   [0:0] tmp_262_fu_3514_p3;
wire   [0:0] icmp_ln1494_55_fu_3522_p2;
wire   [0:0] or_ln1495_86_fu_3554_p2;
wire   [15:0] zext_ln1495_86_fu_3550_p1;
wire   [0:0] tmp_266_fu_3582_p3;
wire   [0:0] xor_ln1495_87_fu_3590_p2;
wire   [10:0] tmp_267_fu_3596_p3;
wire   [0:0] tmp_265_fu_3568_p3;
wire   [0:0] icmp_ln1494_56_fu_3576_p2;
wire   [0:0] or_ln1495_87_fu_3608_p2;
wire   [15:0] zext_ln1495_87_fu_3604_p1;
wire   [0:0] tmp_269_fu_3636_p3;
wire   [0:0] xor_ln1495_88_fu_3644_p2;
wire   [10:0] tmp_270_fu_3650_p3;
wire   [0:0] tmp_268_fu_3622_p3;
wire   [0:0] icmp_ln1494_57_fu_3630_p2;
wire   [0:0] or_ln1495_88_fu_3662_p2;
wire   [15:0] zext_ln1495_88_fu_3658_p1;
wire   [0:0] tmp_272_fu_3690_p3;
wire   [0:0] xor_ln1495_89_fu_3698_p2;
wire   [10:0] tmp_273_fu_3704_p3;
wire   [0:0] tmp_271_fu_3676_p3;
wire   [0:0] icmp_ln1494_58_fu_3684_p2;
wire   [0:0] or_ln1495_89_fu_3716_p2;
wire   [15:0] zext_ln1495_89_fu_3712_p1;
wire   [0:0] tmp_275_fu_3744_p3;
wire   [0:0] xor_ln1495_90_fu_3752_p2;
wire   [10:0] tmp_276_fu_3758_p3;
wire   [0:0] tmp_274_fu_3730_p3;
wire   [0:0] icmp_ln1494_59_fu_3738_p2;
wire   [0:0] or_ln1495_90_fu_3770_p2;
wire   [15:0] zext_ln1495_90_fu_3766_p1;
wire   [0:0] tmp_278_fu_3798_p3;
wire   [0:0] xor_ln1495_91_fu_3806_p2;
wire   [10:0] tmp_279_fu_3812_p3;
wire   [0:0] tmp_277_fu_3784_p3;
wire   [0:0] icmp_ln1494_60_fu_3792_p2;
wire   [0:0] or_ln1495_91_fu_3824_p2;
wire   [15:0] zext_ln1495_91_fu_3820_p1;
wire   [0:0] tmp_281_fu_3852_p3;
wire   [0:0] xor_ln1495_92_fu_3860_p2;
wire   [10:0] tmp_282_fu_3866_p3;
wire   [0:0] tmp_280_fu_3838_p3;
wire   [0:0] icmp_ln1494_61_fu_3846_p2;
wire   [0:0] or_ln1495_92_fu_3878_p2;
wire   [15:0] zext_ln1495_92_fu_3874_p1;
wire   [0:0] tmp_284_fu_3906_p3;
wire   [0:0] xor_ln1495_93_fu_3914_p2;
wire   [10:0] tmp_285_fu_3920_p3;
wire   [0:0] tmp_283_fu_3892_p3;
wire   [0:0] icmp_ln1494_62_fu_3900_p2;
wire   [0:0] or_ln1495_93_fu_3932_p2;
wire   [15:0] zext_ln1495_93_fu_3928_p1;
wire   [0:0] tmp_287_fu_3960_p3;
wire   [0:0] xor_ln1495_94_fu_3968_p2;
wire   [10:0] tmp_288_fu_3974_p3;
wire   [0:0] tmp_286_fu_3946_p3;
wire   [0:0] icmp_ln1494_63_fu_3954_p2;
wire   [0:0] or_ln1495_94_fu_3986_p2;
wire   [15:0] zext_ln1495_94_fu_3982_p1;
wire   [15:0] select_ln1495_fu_590_p3;
wire   [15:0] select_ln1495_32_fu_644_p3;
wire   [15:0] select_ln1495_33_fu_698_p3;
wire   [15:0] select_ln1495_34_fu_752_p3;
wire   [15:0] select_ln1495_35_fu_806_p3;
wire   [15:0] select_ln1495_36_fu_860_p3;
wire   [15:0] select_ln1495_37_fu_914_p3;
wire   [15:0] select_ln1495_38_fu_968_p3;
wire   [15:0] select_ln1495_39_fu_1022_p3;
wire   [15:0] select_ln1495_40_fu_1076_p3;
wire   [15:0] select_ln1495_41_fu_1130_p3;
wire   [15:0] select_ln1495_42_fu_1184_p3;
wire   [15:0] select_ln1495_43_fu_1238_p3;
wire   [15:0] select_ln1495_44_fu_1292_p3;
wire   [15:0] select_ln1495_45_fu_1346_p3;
wire   [15:0] select_ln1495_46_fu_1400_p3;
wire   [15:0] select_ln1495_47_fu_1454_p3;
wire   [15:0] select_ln1495_48_fu_1508_p3;
wire   [15:0] select_ln1495_49_fu_1562_p3;
wire   [15:0] select_ln1495_50_fu_1616_p3;
wire   [15:0] select_ln1495_51_fu_1670_p3;
wire   [15:0] select_ln1495_52_fu_1724_p3;
wire   [15:0] select_ln1495_53_fu_1778_p3;
wire   [15:0] select_ln1495_54_fu_1832_p3;
wire   [15:0] select_ln1495_55_fu_1886_p3;
wire   [15:0] select_ln1495_56_fu_1940_p3;
wire   [15:0] select_ln1495_57_fu_1994_p3;
wire   [15:0] select_ln1495_58_fu_2048_p3;
wire   [15:0] select_ln1495_59_fu_2102_p3;
wire   [15:0] select_ln1495_60_fu_2156_p3;
wire   [15:0] select_ln1495_61_fu_2210_p3;
wire   [15:0] select_ln1495_62_fu_2264_p3;
wire   [15:0] select_ln1495_63_fu_2318_p3;
wire   [15:0] select_ln1495_64_fu_2372_p3;
wire   [15:0] select_ln1495_65_fu_2426_p3;
wire   [15:0] select_ln1495_66_fu_2480_p3;
wire   [15:0] select_ln1495_67_fu_2534_p3;
wire   [15:0] select_ln1495_68_fu_2588_p3;
wire   [15:0] select_ln1495_69_fu_2642_p3;
wire   [15:0] select_ln1495_70_fu_2696_p3;
wire   [15:0] select_ln1495_71_fu_2750_p3;
wire   [15:0] select_ln1495_72_fu_2804_p3;
wire   [15:0] select_ln1495_73_fu_2858_p3;
wire   [15:0] select_ln1495_74_fu_2912_p3;
wire   [15:0] select_ln1495_75_fu_2966_p3;
wire   [15:0] select_ln1495_76_fu_3020_p3;
wire   [15:0] select_ln1495_77_fu_3074_p3;
wire   [15:0] select_ln1495_78_fu_3128_p3;
wire   [15:0] select_ln1495_79_fu_3182_p3;
wire   [15:0] select_ln1495_80_fu_3236_p3;
wire   [15:0] select_ln1495_81_fu_3290_p3;
wire   [15:0] select_ln1495_82_fu_3344_p3;
wire   [15:0] select_ln1495_83_fu_3398_p3;
wire   [15:0] select_ln1495_84_fu_3452_p3;
wire   [15:0] select_ln1495_85_fu_3506_p3;
wire   [15:0] select_ln1495_86_fu_3560_p3;
wire   [15:0] select_ln1495_87_fu_3614_p3;
wire   [15:0] select_ln1495_88_fu_3668_p3;
wire   [15:0] select_ln1495_89_fu_3722_p3;
wire   [15:0] select_ln1495_90_fu_3776_p3;
wire   [15:0] select_ln1495_91_fu_3830_p3;
wire   [15:0] select_ln1495_92_fu_3884_p3;
wire   [15:0] select_ln1495_93_fu_3938_p3;
wire   [15:0] select_ln1495_94_fu_3992_p3;

assign ap_ready = 1'b1;

assign ap_return_0 = select_ln1495_fu_590_p3;

assign ap_return_1 = select_ln1495_32_fu_644_p3;

assign ap_return_10 = select_ln1495_41_fu_1130_p3;

assign ap_return_11 = select_ln1495_42_fu_1184_p3;

assign ap_return_12 = select_ln1495_43_fu_1238_p3;

assign ap_return_13 = select_ln1495_44_fu_1292_p3;

assign ap_return_14 = select_ln1495_45_fu_1346_p3;

assign ap_return_15 = select_ln1495_46_fu_1400_p3;

assign ap_return_16 = select_ln1495_47_fu_1454_p3;

assign ap_return_17 = select_ln1495_48_fu_1508_p3;

assign ap_return_18 = select_ln1495_49_fu_1562_p3;

assign ap_return_19 = select_ln1495_50_fu_1616_p3;

assign ap_return_2 = select_ln1495_33_fu_698_p3;

assign ap_return_20 = select_ln1495_51_fu_1670_p3;

assign ap_return_21 = select_ln1495_52_fu_1724_p3;

assign ap_return_22 = select_ln1495_53_fu_1778_p3;

assign ap_return_23 = select_ln1495_54_fu_1832_p3;

assign ap_return_24 = select_ln1495_55_fu_1886_p3;

assign ap_return_25 = select_ln1495_56_fu_1940_p3;

assign ap_return_26 = select_ln1495_57_fu_1994_p3;

assign ap_return_27 = select_ln1495_58_fu_2048_p3;

assign ap_return_28 = select_ln1495_59_fu_2102_p3;

assign ap_return_29 = select_ln1495_60_fu_2156_p3;

assign ap_return_3 = select_ln1495_34_fu_752_p3;

assign ap_return_30 = select_ln1495_61_fu_2210_p3;

assign ap_return_31 = select_ln1495_62_fu_2264_p3;

assign ap_return_32 = select_ln1495_63_fu_2318_p3;

assign ap_return_33 = select_ln1495_64_fu_2372_p3;

assign ap_return_34 = select_ln1495_65_fu_2426_p3;

assign ap_return_35 = select_ln1495_66_fu_2480_p3;

assign ap_return_36 = select_ln1495_67_fu_2534_p3;

assign ap_return_37 = select_ln1495_68_fu_2588_p3;

assign ap_return_38 = select_ln1495_69_fu_2642_p3;

assign ap_return_39 = select_ln1495_70_fu_2696_p3;

assign ap_return_4 = select_ln1495_35_fu_806_p3;

assign ap_return_40 = select_ln1495_71_fu_2750_p3;

assign ap_return_41 = select_ln1495_72_fu_2804_p3;

assign ap_return_42 = select_ln1495_73_fu_2858_p3;

assign ap_return_43 = select_ln1495_74_fu_2912_p3;

assign ap_return_44 = select_ln1495_75_fu_2966_p3;

assign ap_return_45 = select_ln1495_76_fu_3020_p3;

assign ap_return_46 = select_ln1495_77_fu_3074_p3;

assign ap_return_47 = select_ln1495_78_fu_3128_p3;

assign ap_return_48 = select_ln1495_79_fu_3182_p3;

assign ap_return_49 = select_ln1495_80_fu_3236_p3;

assign ap_return_5 = select_ln1495_36_fu_860_p3;

assign ap_return_50 = select_ln1495_81_fu_3290_p3;

assign ap_return_51 = select_ln1495_82_fu_3344_p3;

assign ap_return_52 = select_ln1495_83_fu_3398_p3;

assign ap_return_53 = select_ln1495_84_fu_3452_p3;

assign ap_return_54 = select_ln1495_85_fu_3506_p3;

assign ap_return_55 = select_ln1495_86_fu_3560_p3;

assign ap_return_56 = select_ln1495_87_fu_3614_p3;

assign ap_return_57 = select_ln1495_88_fu_3668_p3;

assign ap_return_58 = select_ln1495_89_fu_3722_p3;

assign ap_return_59 = select_ln1495_90_fu_3776_p3;

assign ap_return_6 = select_ln1495_37_fu_914_p3;

assign ap_return_60 = select_ln1495_91_fu_3830_p3;

assign ap_return_61 = select_ln1495_92_fu_3884_p3;

assign ap_return_62 = select_ln1495_93_fu_3938_p3;

assign ap_return_63 = select_ln1495_94_fu_3992_p3;

assign ap_return_7 = select_ln1495_38_fu_968_p3;

assign ap_return_8 = select_ln1495_39_fu_1022_p3;

assign ap_return_9 = select_ln1495_40_fu_1076_p3;

assign icmp_ln1494_10_fu_1092_p2 = (((data_10_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_11_fu_1146_p2 = (((data_11_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_12_fu_1200_p2 = (((data_12_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_13_fu_1254_p2 = (((data_13_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_14_fu_1308_p2 = (((data_14_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_15_fu_1362_p2 = (((data_15_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_16_fu_1416_p2 = (((data_16_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_17_fu_1470_p2 = (((data_17_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_18_fu_1524_p2 = (((data_18_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_19_fu_1578_p2 = (((data_19_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_1_fu_606_p2 = (((data_1_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_20_fu_1632_p2 = (((data_20_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_21_fu_1686_p2 = (((data_21_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_22_fu_1740_p2 = (((data_22_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_23_fu_1794_p2 = (((data_23_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_24_fu_1848_p2 = (((data_24_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_25_fu_1902_p2 = (((data_25_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_26_fu_1956_p2 = (((data_26_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_27_fu_2010_p2 = (((data_27_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_28_fu_2064_p2 = (((data_28_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_29_fu_2118_p2 = (((data_29_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_2_fu_660_p2 = (((data_2_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_30_fu_2172_p2 = (((data_30_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_31_fu_2226_p2 = (((data_31_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_32_fu_2280_p2 = (((data_32_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_33_fu_2334_p2 = (((data_33_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_34_fu_2388_p2 = (((data_34_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_35_fu_2442_p2 = (((data_35_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_36_fu_2496_p2 = (((data_36_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_37_fu_2550_p2 = (((data_37_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_38_fu_2604_p2 = (((data_38_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_39_fu_2658_p2 = (((data_39_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_3_fu_714_p2 = (((data_3_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_40_fu_2712_p2 = (((data_40_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_41_fu_2766_p2 = (((data_41_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_42_fu_2820_p2 = (((data_42_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_43_fu_2874_p2 = (((data_43_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_44_fu_2928_p2 = (((data_44_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_45_fu_2982_p2 = (((data_45_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_46_fu_3036_p2 = (((data_46_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_47_fu_3090_p2 = (((data_47_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_48_fu_3144_p2 = (((data_48_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_49_fu_3198_p2 = (((data_49_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_4_fu_768_p2 = (((data_4_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_50_fu_3252_p2 = (((data_50_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_51_fu_3306_p2 = (((data_51_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_52_fu_3360_p2 = (((data_52_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_53_fu_3414_p2 = (((data_53_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_54_fu_3468_p2 = (((data_54_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_55_fu_3522_p2 = (((data_55_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_56_fu_3576_p2 = (((data_56_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_57_fu_3630_p2 = (((data_57_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_58_fu_3684_p2 = (((data_58_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_59_fu_3738_p2 = (((data_59_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_5_fu_822_p2 = (((data_5_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_60_fu_3792_p2 = (((data_60_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_61_fu_3846_p2 = (((data_61_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_62_fu_3900_p2 = (((data_62_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_63_fu_3954_p2 = (((data_63_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_6_fu_876_p2 = (((data_6_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_7_fu_930_p2 = (((data_7_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_8_fu_984_p2 = (((data_8_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_9_fu_1038_p2 = (((data_9_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign icmp_ln1494_fu_552_p2 = (((data_0_V_read) > (16'd1024)) ? 1'b1 : 1'b0);

assign or_ln1495_32_fu_638_p2 = (tmp_100_fu_598_p3 | icmp_ln1494_1_fu_606_p2);

assign or_ln1495_33_fu_692_p2 = (tmp_103_fu_652_p3 | icmp_ln1494_2_fu_660_p2);

assign or_ln1495_34_fu_746_p2 = (tmp_106_fu_706_p3 | icmp_ln1494_3_fu_714_p2);

assign or_ln1495_35_fu_800_p2 = (tmp_109_fu_760_p3 | icmp_ln1494_4_fu_768_p2);

assign or_ln1495_36_fu_854_p2 = (tmp_112_fu_814_p3 | icmp_ln1494_5_fu_822_p2);

assign or_ln1495_37_fu_908_p2 = (tmp_115_fu_868_p3 | icmp_ln1494_6_fu_876_p2);

assign or_ln1495_38_fu_962_p2 = (tmp_118_fu_922_p3 | icmp_ln1494_7_fu_930_p2);

assign or_ln1495_39_fu_1016_p2 = (tmp_121_fu_976_p3 | icmp_ln1494_8_fu_984_p2);

assign or_ln1495_40_fu_1070_p2 = (tmp_124_fu_1030_p3 | icmp_ln1494_9_fu_1038_p2);

assign or_ln1495_41_fu_1124_p2 = (tmp_127_fu_1084_p3 | icmp_ln1494_10_fu_1092_p2);

assign or_ln1495_42_fu_1178_p2 = (tmp_130_fu_1138_p3 | icmp_ln1494_11_fu_1146_p2);

assign or_ln1495_43_fu_1232_p2 = (tmp_133_fu_1192_p3 | icmp_ln1494_12_fu_1200_p2);

assign or_ln1495_44_fu_1286_p2 = (tmp_136_fu_1246_p3 | icmp_ln1494_13_fu_1254_p2);

assign or_ln1495_45_fu_1340_p2 = (tmp_139_fu_1300_p3 | icmp_ln1494_14_fu_1308_p2);

assign or_ln1495_46_fu_1394_p2 = (tmp_142_fu_1354_p3 | icmp_ln1494_15_fu_1362_p2);

assign or_ln1495_47_fu_1448_p2 = (tmp_145_fu_1408_p3 | icmp_ln1494_16_fu_1416_p2);

assign or_ln1495_48_fu_1502_p2 = (tmp_148_fu_1462_p3 | icmp_ln1494_17_fu_1470_p2);

assign or_ln1495_49_fu_1556_p2 = (tmp_151_fu_1516_p3 | icmp_ln1494_18_fu_1524_p2);

assign or_ln1495_50_fu_1610_p2 = (tmp_154_fu_1570_p3 | icmp_ln1494_19_fu_1578_p2);

assign or_ln1495_51_fu_1664_p2 = (tmp_157_fu_1624_p3 | icmp_ln1494_20_fu_1632_p2);

assign or_ln1495_52_fu_1718_p2 = (tmp_160_fu_1678_p3 | icmp_ln1494_21_fu_1686_p2);

assign or_ln1495_53_fu_1772_p2 = (tmp_163_fu_1732_p3 | icmp_ln1494_22_fu_1740_p2);

assign or_ln1495_54_fu_1826_p2 = (tmp_166_fu_1786_p3 | icmp_ln1494_23_fu_1794_p2);

assign or_ln1495_55_fu_1880_p2 = (tmp_169_fu_1840_p3 | icmp_ln1494_24_fu_1848_p2);

assign or_ln1495_56_fu_1934_p2 = (tmp_172_fu_1894_p3 | icmp_ln1494_25_fu_1902_p2);

assign or_ln1495_57_fu_1988_p2 = (tmp_175_fu_1948_p3 | icmp_ln1494_26_fu_1956_p2);

assign or_ln1495_58_fu_2042_p2 = (tmp_178_fu_2002_p3 | icmp_ln1494_27_fu_2010_p2);

assign or_ln1495_59_fu_2096_p2 = (tmp_181_fu_2056_p3 | icmp_ln1494_28_fu_2064_p2);

assign or_ln1495_60_fu_2150_p2 = (tmp_184_fu_2110_p3 | icmp_ln1494_29_fu_2118_p2);

assign or_ln1495_61_fu_2204_p2 = (tmp_187_fu_2164_p3 | icmp_ln1494_30_fu_2172_p2);

assign or_ln1495_62_fu_2258_p2 = (tmp_190_fu_2218_p3 | icmp_ln1494_31_fu_2226_p2);

assign or_ln1495_63_fu_2312_p2 = (tmp_193_fu_2272_p3 | icmp_ln1494_32_fu_2280_p2);

assign or_ln1495_64_fu_2366_p2 = (tmp_196_fu_2326_p3 | icmp_ln1494_33_fu_2334_p2);

assign or_ln1495_65_fu_2420_p2 = (tmp_199_fu_2380_p3 | icmp_ln1494_34_fu_2388_p2);

assign or_ln1495_66_fu_2474_p2 = (tmp_202_fu_2434_p3 | icmp_ln1494_35_fu_2442_p2);

assign or_ln1495_67_fu_2528_p2 = (tmp_205_fu_2488_p3 | icmp_ln1494_36_fu_2496_p2);

assign or_ln1495_68_fu_2582_p2 = (tmp_208_fu_2542_p3 | icmp_ln1494_37_fu_2550_p2);

assign or_ln1495_69_fu_2636_p2 = (tmp_211_fu_2596_p3 | icmp_ln1494_38_fu_2604_p2);

assign or_ln1495_70_fu_2690_p2 = (tmp_214_fu_2650_p3 | icmp_ln1494_39_fu_2658_p2);

assign or_ln1495_71_fu_2744_p2 = (tmp_217_fu_2704_p3 | icmp_ln1494_40_fu_2712_p2);

assign or_ln1495_72_fu_2798_p2 = (tmp_220_fu_2758_p3 | icmp_ln1494_41_fu_2766_p2);

assign or_ln1495_73_fu_2852_p2 = (tmp_223_fu_2812_p3 | icmp_ln1494_42_fu_2820_p2);

assign or_ln1495_74_fu_2906_p2 = (tmp_226_fu_2866_p3 | icmp_ln1494_43_fu_2874_p2);

assign or_ln1495_75_fu_2960_p2 = (tmp_229_fu_2920_p3 | icmp_ln1494_44_fu_2928_p2);

assign or_ln1495_76_fu_3014_p2 = (tmp_232_fu_2974_p3 | icmp_ln1494_45_fu_2982_p2);

assign or_ln1495_77_fu_3068_p2 = (tmp_235_fu_3028_p3 | icmp_ln1494_46_fu_3036_p2);

assign or_ln1495_78_fu_3122_p2 = (tmp_238_fu_3082_p3 | icmp_ln1494_47_fu_3090_p2);

assign or_ln1495_79_fu_3176_p2 = (tmp_241_fu_3136_p3 | icmp_ln1494_48_fu_3144_p2);

assign or_ln1495_80_fu_3230_p2 = (tmp_244_fu_3190_p3 | icmp_ln1494_49_fu_3198_p2);

assign or_ln1495_81_fu_3284_p2 = (tmp_247_fu_3244_p3 | icmp_ln1494_50_fu_3252_p2);

assign or_ln1495_82_fu_3338_p2 = (tmp_250_fu_3298_p3 | icmp_ln1494_51_fu_3306_p2);

assign or_ln1495_83_fu_3392_p2 = (tmp_253_fu_3352_p3 | icmp_ln1494_52_fu_3360_p2);

assign or_ln1495_84_fu_3446_p2 = (tmp_256_fu_3406_p3 | icmp_ln1494_53_fu_3414_p2);

assign or_ln1495_85_fu_3500_p2 = (tmp_259_fu_3460_p3 | icmp_ln1494_54_fu_3468_p2);

assign or_ln1495_86_fu_3554_p2 = (tmp_262_fu_3514_p3 | icmp_ln1494_55_fu_3522_p2);

assign or_ln1495_87_fu_3608_p2 = (tmp_265_fu_3568_p3 | icmp_ln1494_56_fu_3576_p2);

assign or_ln1495_88_fu_3662_p2 = (tmp_268_fu_3622_p3 | icmp_ln1494_57_fu_3630_p2);

assign or_ln1495_89_fu_3716_p2 = (tmp_271_fu_3676_p3 | icmp_ln1494_58_fu_3684_p2);

assign or_ln1495_90_fu_3770_p2 = (tmp_274_fu_3730_p3 | icmp_ln1494_59_fu_3738_p2);

assign or_ln1495_91_fu_3824_p2 = (tmp_277_fu_3784_p3 | icmp_ln1494_60_fu_3792_p2);

assign or_ln1495_92_fu_3878_p2 = (tmp_280_fu_3838_p3 | icmp_ln1494_61_fu_3846_p2);

assign or_ln1495_93_fu_3932_p2 = (tmp_283_fu_3892_p3 | icmp_ln1494_62_fu_3900_p2);

assign or_ln1495_94_fu_3986_p2 = (tmp_286_fu_3946_p3 | icmp_ln1494_63_fu_3954_p2);

assign or_ln1495_fu_584_p2 = (tmp_97_fu_544_p3 | icmp_ln1494_fu_552_p2);

assign select_ln1495_32_fu_644_p3 = ((or_ln1495_32_fu_638_p2[0:0] == 1'b1) ? zext_ln1495_32_fu_634_p1 : data_1_V_read);

assign select_ln1495_33_fu_698_p3 = ((or_ln1495_33_fu_692_p2[0:0] == 1'b1) ? zext_ln1495_33_fu_688_p1 : data_2_V_read);

assign select_ln1495_34_fu_752_p3 = ((or_ln1495_34_fu_746_p2[0:0] == 1'b1) ? zext_ln1495_34_fu_742_p1 : data_3_V_read);

assign select_ln1495_35_fu_806_p3 = ((or_ln1495_35_fu_800_p2[0:0] == 1'b1) ? zext_ln1495_35_fu_796_p1 : data_4_V_read);

assign select_ln1495_36_fu_860_p3 = ((or_ln1495_36_fu_854_p2[0:0] == 1'b1) ? zext_ln1495_36_fu_850_p1 : data_5_V_read);

assign select_ln1495_37_fu_914_p3 = ((or_ln1495_37_fu_908_p2[0:0] == 1'b1) ? zext_ln1495_37_fu_904_p1 : data_6_V_read);

assign select_ln1495_38_fu_968_p3 = ((or_ln1495_38_fu_962_p2[0:0] == 1'b1) ? zext_ln1495_38_fu_958_p1 : data_7_V_read);

assign select_ln1495_39_fu_1022_p3 = ((or_ln1495_39_fu_1016_p2[0:0] == 1'b1) ? zext_ln1495_39_fu_1012_p1 : data_8_V_read);

assign select_ln1495_40_fu_1076_p3 = ((or_ln1495_40_fu_1070_p2[0:0] == 1'b1) ? zext_ln1495_40_fu_1066_p1 : data_9_V_read);

assign select_ln1495_41_fu_1130_p3 = ((or_ln1495_41_fu_1124_p2[0:0] == 1'b1) ? zext_ln1495_41_fu_1120_p1 : data_10_V_read);

assign select_ln1495_42_fu_1184_p3 = ((or_ln1495_42_fu_1178_p2[0:0] == 1'b1) ? zext_ln1495_42_fu_1174_p1 : data_11_V_read);

assign select_ln1495_43_fu_1238_p3 = ((or_ln1495_43_fu_1232_p2[0:0] == 1'b1) ? zext_ln1495_43_fu_1228_p1 : data_12_V_read);

assign select_ln1495_44_fu_1292_p3 = ((or_ln1495_44_fu_1286_p2[0:0] == 1'b1) ? zext_ln1495_44_fu_1282_p1 : data_13_V_read);

assign select_ln1495_45_fu_1346_p3 = ((or_ln1495_45_fu_1340_p2[0:0] == 1'b1) ? zext_ln1495_45_fu_1336_p1 : data_14_V_read);

assign select_ln1495_46_fu_1400_p3 = ((or_ln1495_46_fu_1394_p2[0:0] == 1'b1) ? zext_ln1495_46_fu_1390_p1 : data_15_V_read);

assign select_ln1495_47_fu_1454_p3 = ((or_ln1495_47_fu_1448_p2[0:0] == 1'b1) ? zext_ln1495_47_fu_1444_p1 : data_16_V_read);

assign select_ln1495_48_fu_1508_p3 = ((or_ln1495_48_fu_1502_p2[0:0] == 1'b1) ? zext_ln1495_48_fu_1498_p1 : data_17_V_read);

assign select_ln1495_49_fu_1562_p3 = ((or_ln1495_49_fu_1556_p2[0:0] == 1'b1) ? zext_ln1495_49_fu_1552_p1 : data_18_V_read);

assign select_ln1495_50_fu_1616_p3 = ((or_ln1495_50_fu_1610_p2[0:0] == 1'b1) ? zext_ln1495_50_fu_1606_p1 : data_19_V_read);

assign select_ln1495_51_fu_1670_p3 = ((or_ln1495_51_fu_1664_p2[0:0] == 1'b1) ? zext_ln1495_51_fu_1660_p1 : data_20_V_read);

assign select_ln1495_52_fu_1724_p3 = ((or_ln1495_52_fu_1718_p2[0:0] == 1'b1) ? zext_ln1495_52_fu_1714_p1 : data_21_V_read);

assign select_ln1495_53_fu_1778_p3 = ((or_ln1495_53_fu_1772_p2[0:0] == 1'b1) ? zext_ln1495_53_fu_1768_p1 : data_22_V_read);

assign select_ln1495_54_fu_1832_p3 = ((or_ln1495_54_fu_1826_p2[0:0] == 1'b1) ? zext_ln1495_54_fu_1822_p1 : data_23_V_read);

assign select_ln1495_55_fu_1886_p3 = ((or_ln1495_55_fu_1880_p2[0:0] == 1'b1) ? zext_ln1495_55_fu_1876_p1 : data_24_V_read);

assign select_ln1495_56_fu_1940_p3 = ((or_ln1495_56_fu_1934_p2[0:0] == 1'b1) ? zext_ln1495_56_fu_1930_p1 : data_25_V_read);

assign select_ln1495_57_fu_1994_p3 = ((or_ln1495_57_fu_1988_p2[0:0] == 1'b1) ? zext_ln1495_57_fu_1984_p1 : data_26_V_read);

assign select_ln1495_58_fu_2048_p3 = ((or_ln1495_58_fu_2042_p2[0:0] == 1'b1) ? zext_ln1495_58_fu_2038_p1 : data_27_V_read);

assign select_ln1495_59_fu_2102_p3 = ((or_ln1495_59_fu_2096_p2[0:0] == 1'b1) ? zext_ln1495_59_fu_2092_p1 : data_28_V_read);

assign select_ln1495_60_fu_2156_p3 = ((or_ln1495_60_fu_2150_p2[0:0] == 1'b1) ? zext_ln1495_60_fu_2146_p1 : data_29_V_read);

assign select_ln1495_61_fu_2210_p3 = ((or_ln1495_61_fu_2204_p2[0:0] == 1'b1) ? zext_ln1495_61_fu_2200_p1 : data_30_V_read);

assign select_ln1495_62_fu_2264_p3 = ((or_ln1495_62_fu_2258_p2[0:0] == 1'b1) ? zext_ln1495_62_fu_2254_p1 : data_31_V_read);

assign select_ln1495_63_fu_2318_p3 = ((or_ln1495_63_fu_2312_p2[0:0] == 1'b1) ? zext_ln1495_63_fu_2308_p1 : data_32_V_read);

assign select_ln1495_64_fu_2372_p3 = ((or_ln1495_64_fu_2366_p2[0:0] == 1'b1) ? zext_ln1495_64_fu_2362_p1 : data_33_V_read);

assign select_ln1495_65_fu_2426_p3 = ((or_ln1495_65_fu_2420_p2[0:0] == 1'b1) ? zext_ln1495_65_fu_2416_p1 : data_34_V_read);

assign select_ln1495_66_fu_2480_p3 = ((or_ln1495_66_fu_2474_p2[0:0] == 1'b1) ? zext_ln1495_66_fu_2470_p1 : data_35_V_read);

assign select_ln1495_67_fu_2534_p3 = ((or_ln1495_67_fu_2528_p2[0:0] == 1'b1) ? zext_ln1495_67_fu_2524_p1 : data_36_V_read);

assign select_ln1495_68_fu_2588_p3 = ((or_ln1495_68_fu_2582_p2[0:0] == 1'b1) ? zext_ln1495_68_fu_2578_p1 : data_37_V_read);

assign select_ln1495_69_fu_2642_p3 = ((or_ln1495_69_fu_2636_p2[0:0] == 1'b1) ? zext_ln1495_69_fu_2632_p1 : data_38_V_read);

assign select_ln1495_70_fu_2696_p3 = ((or_ln1495_70_fu_2690_p2[0:0] == 1'b1) ? zext_ln1495_70_fu_2686_p1 : data_39_V_read);

assign select_ln1495_71_fu_2750_p3 = ((or_ln1495_71_fu_2744_p2[0:0] == 1'b1) ? zext_ln1495_71_fu_2740_p1 : data_40_V_read);

assign select_ln1495_72_fu_2804_p3 = ((or_ln1495_72_fu_2798_p2[0:0] == 1'b1) ? zext_ln1495_72_fu_2794_p1 : data_41_V_read);

assign select_ln1495_73_fu_2858_p3 = ((or_ln1495_73_fu_2852_p2[0:0] == 1'b1) ? zext_ln1495_73_fu_2848_p1 : data_42_V_read);

assign select_ln1495_74_fu_2912_p3 = ((or_ln1495_74_fu_2906_p2[0:0] == 1'b1) ? zext_ln1495_74_fu_2902_p1 : data_43_V_read);

assign select_ln1495_75_fu_2966_p3 = ((or_ln1495_75_fu_2960_p2[0:0] == 1'b1) ? zext_ln1495_75_fu_2956_p1 : data_44_V_read);

assign select_ln1495_76_fu_3020_p3 = ((or_ln1495_76_fu_3014_p2[0:0] == 1'b1) ? zext_ln1495_76_fu_3010_p1 : data_45_V_read);

assign select_ln1495_77_fu_3074_p3 = ((or_ln1495_77_fu_3068_p2[0:0] == 1'b1) ? zext_ln1495_77_fu_3064_p1 : data_46_V_read);

assign select_ln1495_78_fu_3128_p3 = ((or_ln1495_78_fu_3122_p2[0:0] == 1'b1) ? zext_ln1495_78_fu_3118_p1 : data_47_V_read);

assign select_ln1495_79_fu_3182_p3 = ((or_ln1495_79_fu_3176_p2[0:0] == 1'b1) ? zext_ln1495_79_fu_3172_p1 : data_48_V_read);

assign select_ln1495_80_fu_3236_p3 = ((or_ln1495_80_fu_3230_p2[0:0] == 1'b1) ? zext_ln1495_80_fu_3226_p1 : data_49_V_read);

assign select_ln1495_81_fu_3290_p3 = ((or_ln1495_81_fu_3284_p2[0:0] == 1'b1) ? zext_ln1495_81_fu_3280_p1 : data_50_V_read);

assign select_ln1495_82_fu_3344_p3 = ((or_ln1495_82_fu_3338_p2[0:0] == 1'b1) ? zext_ln1495_82_fu_3334_p1 : data_51_V_read);

assign select_ln1495_83_fu_3398_p3 = ((or_ln1495_83_fu_3392_p2[0:0] == 1'b1) ? zext_ln1495_83_fu_3388_p1 : data_52_V_read);

assign select_ln1495_84_fu_3452_p3 = ((or_ln1495_84_fu_3446_p2[0:0] == 1'b1) ? zext_ln1495_84_fu_3442_p1 : data_53_V_read);

assign select_ln1495_85_fu_3506_p3 = ((or_ln1495_85_fu_3500_p2[0:0] == 1'b1) ? zext_ln1495_85_fu_3496_p1 : data_54_V_read);

assign select_ln1495_86_fu_3560_p3 = ((or_ln1495_86_fu_3554_p2[0:0] == 1'b1) ? zext_ln1495_86_fu_3550_p1 : data_55_V_read);

assign select_ln1495_87_fu_3614_p3 = ((or_ln1495_87_fu_3608_p2[0:0] == 1'b1) ? zext_ln1495_87_fu_3604_p1 : data_56_V_read);

assign select_ln1495_88_fu_3668_p3 = ((or_ln1495_88_fu_3662_p2[0:0] == 1'b1) ? zext_ln1495_88_fu_3658_p1 : data_57_V_read);

assign select_ln1495_89_fu_3722_p3 = ((or_ln1495_89_fu_3716_p2[0:0] == 1'b1) ? zext_ln1495_89_fu_3712_p1 : data_58_V_read);

assign select_ln1495_90_fu_3776_p3 = ((or_ln1495_90_fu_3770_p2[0:0] == 1'b1) ? zext_ln1495_90_fu_3766_p1 : data_59_V_read);

assign select_ln1495_91_fu_3830_p3 = ((or_ln1495_91_fu_3824_p2[0:0] == 1'b1) ? zext_ln1495_91_fu_3820_p1 : data_60_V_read);

assign select_ln1495_92_fu_3884_p3 = ((or_ln1495_92_fu_3878_p2[0:0] == 1'b1) ? zext_ln1495_92_fu_3874_p1 : data_61_V_read);

assign select_ln1495_93_fu_3938_p3 = ((or_ln1495_93_fu_3932_p2[0:0] == 1'b1) ? zext_ln1495_93_fu_3928_p1 : data_62_V_read);

assign select_ln1495_94_fu_3992_p3 = ((or_ln1495_94_fu_3986_p2[0:0] == 1'b1) ? zext_ln1495_94_fu_3982_p1 : data_63_V_read);

assign select_ln1495_fu_590_p3 = ((or_ln1495_fu_584_p2[0:0] == 1'b1) ? zext_ln1495_fu_580_p1 : data_0_V_read);

assign tmp_100_fu_598_p3 = data_1_V_read[32'd15];

assign tmp_101_fu_612_p3 = data_1_V_read[32'd15];

assign tmp_102_fu_626_p3 = {{xor_ln1495_32_fu_620_p2}, {10'd0}};

assign tmp_103_fu_652_p3 = data_2_V_read[32'd15];

assign tmp_104_fu_666_p3 = data_2_V_read[32'd15];

assign tmp_105_fu_680_p3 = {{xor_ln1495_33_fu_674_p2}, {10'd0}};

assign tmp_106_fu_706_p3 = data_3_V_read[32'd15];

assign tmp_107_fu_720_p3 = data_3_V_read[32'd15];

assign tmp_108_fu_734_p3 = {{xor_ln1495_34_fu_728_p2}, {10'd0}};

assign tmp_109_fu_760_p3 = data_4_V_read[32'd15];

assign tmp_110_fu_774_p3 = data_4_V_read[32'd15];

assign tmp_111_fu_788_p3 = {{xor_ln1495_35_fu_782_p2}, {10'd0}};

assign tmp_112_fu_814_p3 = data_5_V_read[32'd15];

assign tmp_113_fu_828_p3 = data_5_V_read[32'd15];

assign tmp_114_fu_842_p3 = {{xor_ln1495_36_fu_836_p2}, {10'd0}};

assign tmp_115_fu_868_p3 = data_6_V_read[32'd15];

assign tmp_116_fu_882_p3 = data_6_V_read[32'd15];

assign tmp_117_fu_896_p3 = {{xor_ln1495_37_fu_890_p2}, {10'd0}};

assign tmp_118_fu_922_p3 = data_7_V_read[32'd15];

assign tmp_119_fu_936_p3 = data_7_V_read[32'd15];

assign tmp_120_fu_950_p3 = {{xor_ln1495_38_fu_944_p2}, {10'd0}};

assign tmp_121_fu_976_p3 = data_8_V_read[32'd15];

assign tmp_122_fu_990_p3 = data_8_V_read[32'd15];

assign tmp_123_fu_1004_p3 = {{xor_ln1495_39_fu_998_p2}, {10'd0}};

assign tmp_124_fu_1030_p3 = data_9_V_read[32'd15];

assign tmp_125_fu_1044_p3 = data_9_V_read[32'd15];

assign tmp_126_fu_1058_p3 = {{xor_ln1495_40_fu_1052_p2}, {10'd0}};

assign tmp_127_fu_1084_p3 = data_10_V_read[32'd15];

assign tmp_128_fu_1098_p3 = data_10_V_read[32'd15];

assign tmp_129_fu_1112_p3 = {{xor_ln1495_41_fu_1106_p2}, {10'd0}};

assign tmp_130_fu_1138_p3 = data_11_V_read[32'd15];

assign tmp_131_fu_1152_p3 = data_11_V_read[32'd15];

assign tmp_132_fu_1166_p3 = {{xor_ln1495_42_fu_1160_p2}, {10'd0}};

assign tmp_133_fu_1192_p3 = data_12_V_read[32'd15];

assign tmp_134_fu_1206_p3 = data_12_V_read[32'd15];

assign tmp_135_fu_1220_p3 = {{xor_ln1495_43_fu_1214_p2}, {10'd0}};

assign tmp_136_fu_1246_p3 = data_13_V_read[32'd15];

assign tmp_137_fu_1260_p3 = data_13_V_read[32'd15];

assign tmp_138_fu_1274_p3 = {{xor_ln1495_44_fu_1268_p2}, {10'd0}};

assign tmp_139_fu_1300_p3 = data_14_V_read[32'd15];

assign tmp_140_fu_1314_p3 = data_14_V_read[32'd15];

assign tmp_141_fu_1328_p3 = {{xor_ln1495_45_fu_1322_p2}, {10'd0}};

assign tmp_142_fu_1354_p3 = data_15_V_read[32'd15];

assign tmp_143_fu_1368_p3 = data_15_V_read[32'd15];

assign tmp_144_fu_1382_p3 = {{xor_ln1495_46_fu_1376_p2}, {10'd0}};

assign tmp_145_fu_1408_p3 = data_16_V_read[32'd15];

assign tmp_146_fu_1422_p3 = data_16_V_read[32'd15];

assign tmp_147_fu_1436_p3 = {{xor_ln1495_47_fu_1430_p2}, {10'd0}};

assign tmp_148_fu_1462_p3 = data_17_V_read[32'd15];

assign tmp_149_fu_1476_p3 = data_17_V_read[32'd15];

assign tmp_150_fu_1490_p3 = {{xor_ln1495_48_fu_1484_p2}, {10'd0}};

assign tmp_151_fu_1516_p3 = data_18_V_read[32'd15];

assign tmp_152_fu_1530_p3 = data_18_V_read[32'd15];

assign tmp_153_fu_1544_p3 = {{xor_ln1495_49_fu_1538_p2}, {10'd0}};

assign tmp_154_fu_1570_p3 = data_19_V_read[32'd15];

assign tmp_155_fu_1584_p3 = data_19_V_read[32'd15];

assign tmp_156_fu_1598_p3 = {{xor_ln1495_50_fu_1592_p2}, {10'd0}};

assign tmp_157_fu_1624_p3 = data_20_V_read[32'd15];

assign tmp_158_fu_1638_p3 = data_20_V_read[32'd15];

assign tmp_159_fu_1652_p3 = {{xor_ln1495_51_fu_1646_p2}, {10'd0}};

assign tmp_160_fu_1678_p3 = data_21_V_read[32'd15];

assign tmp_161_fu_1692_p3 = data_21_V_read[32'd15];

assign tmp_162_fu_1706_p3 = {{xor_ln1495_52_fu_1700_p2}, {10'd0}};

assign tmp_163_fu_1732_p3 = data_22_V_read[32'd15];

assign tmp_164_fu_1746_p3 = data_22_V_read[32'd15];

assign tmp_165_fu_1760_p3 = {{xor_ln1495_53_fu_1754_p2}, {10'd0}};

assign tmp_166_fu_1786_p3 = data_23_V_read[32'd15];

assign tmp_167_fu_1800_p3 = data_23_V_read[32'd15];

assign tmp_168_fu_1814_p3 = {{xor_ln1495_54_fu_1808_p2}, {10'd0}};

assign tmp_169_fu_1840_p3 = data_24_V_read[32'd15];

assign tmp_170_fu_1854_p3 = data_24_V_read[32'd15];

assign tmp_171_fu_1868_p3 = {{xor_ln1495_55_fu_1862_p2}, {10'd0}};

assign tmp_172_fu_1894_p3 = data_25_V_read[32'd15];

assign tmp_173_fu_1908_p3 = data_25_V_read[32'd15];

assign tmp_174_fu_1922_p3 = {{xor_ln1495_56_fu_1916_p2}, {10'd0}};

assign tmp_175_fu_1948_p3 = data_26_V_read[32'd15];

assign tmp_176_fu_1962_p3 = data_26_V_read[32'd15];

assign tmp_177_fu_1976_p3 = {{xor_ln1495_57_fu_1970_p2}, {10'd0}};

assign tmp_178_fu_2002_p3 = data_27_V_read[32'd15];

assign tmp_179_fu_2016_p3 = data_27_V_read[32'd15];

assign tmp_180_fu_2030_p3 = {{xor_ln1495_58_fu_2024_p2}, {10'd0}};

assign tmp_181_fu_2056_p3 = data_28_V_read[32'd15];

assign tmp_182_fu_2070_p3 = data_28_V_read[32'd15];

assign tmp_183_fu_2084_p3 = {{xor_ln1495_59_fu_2078_p2}, {10'd0}};

assign tmp_184_fu_2110_p3 = data_29_V_read[32'd15];

assign tmp_185_fu_2124_p3 = data_29_V_read[32'd15];

assign tmp_186_fu_2138_p3 = {{xor_ln1495_60_fu_2132_p2}, {10'd0}};

assign tmp_187_fu_2164_p3 = data_30_V_read[32'd15];

assign tmp_188_fu_2178_p3 = data_30_V_read[32'd15];

assign tmp_189_fu_2192_p3 = {{xor_ln1495_61_fu_2186_p2}, {10'd0}};

assign tmp_190_fu_2218_p3 = data_31_V_read[32'd15];

assign tmp_191_fu_2232_p3 = data_31_V_read[32'd15];

assign tmp_192_fu_2246_p3 = {{xor_ln1495_62_fu_2240_p2}, {10'd0}};

assign tmp_193_fu_2272_p3 = data_32_V_read[32'd15];

assign tmp_194_fu_2286_p3 = data_32_V_read[32'd15];

assign tmp_195_fu_2300_p3 = {{xor_ln1495_63_fu_2294_p2}, {10'd0}};

assign tmp_196_fu_2326_p3 = data_33_V_read[32'd15];

assign tmp_197_fu_2340_p3 = data_33_V_read[32'd15];

assign tmp_198_fu_2354_p3 = {{xor_ln1495_64_fu_2348_p2}, {10'd0}};

assign tmp_199_fu_2380_p3 = data_34_V_read[32'd15];

assign tmp_200_fu_2394_p3 = data_34_V_read[32'd15];

assign tmp_201_fu_2408_p3 = {{xor_ln1495_65_fu_2402_p2}, {10'd0}};

assign tmp_202_fu_2434_p3 = data_35_V_read[32'd15];

assign tmp_203_fu_2448_p3 = data_35_V_read[32'd15];

assign tmp_204_fu_2462_p3 = {{xor_ln1495_66_fu_2456_p2}, {10'd0}};

assign tmp_205_fu_2488_p3 = data_36_V_read[32'd15];

assign tmp_206_fu_2502_p3 = data_36_V_read[32'd15];

assign tmp_207_fu_2516_p3 = {{xor_ln1495_67_fu_2510_p2}, {10'd0}};

assign tmp_208_fu_2542_p3 = data_37_V_read[32'd15];

assign tmp_209_fu_2556_p3 = data_37_V_read[32'd15];

assign tmp_210_fu_2570_p3 = {{xor_ln1495_68_fu_2564_p2}, {10'd0}};

assign tmp_211_fu_2596_p3 = data_38_V_read[32'd15];

assign tmp_212_fu_2610_p3 = data_38_V_read[32'd15];

assign tmp_213_fu_2624_p3 = {{xor_ln1495_69_fu_2618_p2}, {10'd0}};

assign tmp_214_fu_2650_p3 = data_39_V_read[32'd15];

assign tmp_215_fu_2664_p3 = data_39_V_read[32'd15];

assign tmp_216_fu_2678_p3 = {{xor_ln1495_70_fu_2672_p2}, {10'd0}};

assign tmp_217_fu_2704_p3 = data_40_V_read[32'd15];

assign tmp_218_fu_2718_p3 = data_40_V_read[32'd15];

assign tmp_219_fu_2732_p3 = {{xor_ln1495_71_fu_2726_p2}, {10'd0}};

assign tmp_220_fu_2758_p3 = data_41_V_read[32'd15];

assign tmp_221_fu_2772_p3 = data_41_V_read[32'd15];

assign tmp_222_fu_2786_p3 = {{xor_ln1495_72_fu_2780_p2}, {10'd0}};

assign tmp_223_fu_2812_p3 = data_42_V_read[32'd15];

assign tmp_224_fu_2826_p3 = data_42_V_read[32'd15];

assign tmp_225_fu_2840_p3 = {{xor_ln1495_73_fu_2834_p2}, {10'd0}};

assign tmp_226_fu_2866_p3 = data_43_V_read[32'd15];

assign tmp_227_fu_2880_p3 = data_43_V_read[32'd15];

assign tmp_228_fu_2894_p3 = {{xor_ln1495_74_fu_2888_p2}, {10'd0}};

assign tmp_229_fu_2920_p3 = data_44_V_read[32'd15];

assign tmp_230_fu_2934_p3 = data_44_V_read[32'd15];

assign tmp_231_fu_2948_p3 = {{xor_ln1495_75_fu_2942_p2}, {10'd0}};

assign tmp_232_fu_2974_p3 = data_45_V_read[32'd15];

assign tmp_233_fu_2988_p3 = data_45_V_read[32'd15];

assign tmp_234_fu_3002_p3 = {{xor_ln1495_76_fu_2996_p2}, {10'd0}};

assign tmp_235_fu_3028_p3 = data_46_V_read[32'd15];

assign tmp_236_fu_3042_p3 = data_46_V_read[32'd15];

assign tmp_237_fu_3056_p3 = {{xor_ln1495_77_fu_3050_p2}, {10'd0}};

assign tmp_238_fu_3082_p3 = data_47_V_read[32'd15];

assign tmp_239_fu_3096_p3 = data_47_V_read[32'd15];

assign tmp_240_fu_3110_p3 = {{xor_ln1495_78_fu_3104_p2}, {10'd0}};

assign tmp_241_fu_3136_p3 = data_48_V_read[32'd15];

assign tmp_242_fu_3150_p3 = data_48_V_read[32'd15];

assign tmp_243_fu_3164_p3 = {{xor_ln1495_79_fu_3158_p2}, {10'd0}};

assign tmp_244_fu_3190_p3 = data_49_V_read[32'd15];

assign tmp_245_fu_3204_p3 = data_49_V_read[32'd15];

assign tmp_246_fu_3218_p3 = {{xor_ln1495_80_fu_3212_p2}, {10'd0}};

assign tmp_247_fu_3244_p3 = data_50_V_read[32'd15];

assign tmp_248_fu_3258_p3 = data_50_V_read[32'd15];

assign tmp_249_fu_3272_p3 = {{xor_ln1495_81_fu_3266_p2}, {10'd0}};

assign tmp_250_fu_3298_p3 = data_51_V_read[32'd15];

assign tmp_251_fu_3312_p3 = data_51_V_read[32'd15];

assign tmp_252_fu_3326_p3 = {{xor_ln1495_82_fu_3320_p2}, {10'd0}};

assign tmp_253_fu_3352_p3 = data_52_V_read[32'd15];

assign tmp_254_fu_3366_p3 = data_52_V_read[32'd15];

assign tmp_255_fu_3380_p3 = {{xor_ln1495_83_fu_3374_p2}, {10'd0}};

assign tmp_256_fu_3406_p3 = data_53_V_read[32'd15];

assign tmp_257_fu_3420_p3 = data_53_V_read[32'd15];

assign tmp_258_fu_3434_p3 = {{xor_ln1495_84_fu_3428_p2}, {10'd0}};

assign tmp_259_fu_3460_p3 = data_54_V_read[32'd15];

assign tmp_260_fu_3474_p3 = data_54_V_read[32'd15];

assign tmp_261_fu_3488_p3 = {{xor_ln1495_85_fu_3482_p2}, {10'd0}};

assign tmp_262_fu_3514_p3 = data_55_V_read[32'd15];

assign tmp_263_fu_3528_p3 = data_55_V_read[32'd15];

assign tmp_264_fu_3542_p3 = {{xor_ln1495_86_fu_3536_p2}, {10'd0}};

assign tmp_265_fu_3568_p3 = data_56_V_read[32'd15];

assign tmp_266_fu_3582_p3 = data_56_V_read[32'd15];

assign tmp_267_fu_3596_p3 = {{xor_ln1495_87_fu_3590_p2}, {10'd0}};

assign tmp_268_fu_3622_p3 = data_57_V_read[32'd15];

assign tmp_269_fu_3636_p3 = data_57_V_read[32'd15];

assign tmp_270_fu_3650_p3 = {{xor_ln1495_88_fu_3644_p2}, {10'd0}};

assign tmp_271_fu_3676_p3 = data_58_V_read[32'd15];

assign tmp_272_fu_3690_p3 = data_58_V_read[32'd15];

assign tmp_273_fu_3704_p3 = {{xor_ln1495_89_fu_3698_p2}, {10'd0}};

assign tmp_274_fu_3730_p3 = data_59_V_read[32'd15];

assign tmp_275_fu_3744_p3 = data_59_V_read[32'd15];

assign tmp_276_fu_3758_p3 = {{xor_ln1495_90_fu_3752_p2}, {10'd0}};

assign tmp_277_fu_3784_p3 = data_60_V_read[32'd15];

assign tmp_278_fu_3798_p3 = data_60_V_read[32'd15];

assign tmp_279_fu_3812_p3 = {{xor_ln1495_91_fu_3806_p2}, {10'd0}};

assign tmp_280_fu_3838_p3 = data_61_V_read[32'd15];

assign tmp_281_fu_3852_p3 = data_61_V_read[32'd15];

assign tmp_282_fu_3866_p3 = {{xor_ln1495_92_fu_3860_p2}, {10'd0}};

assign tmp_283_fu_3892_p3 = data_62_V_read[32'd15];

assign tmp_284_fu_3906_p3 = data_62_V_read[32'd15];

assign tmp_285_fu_3920_p3 = {{xor_ln1495_93_fu_3914_p2}, {10'd0}};

assign tmp_286_fu_3946_p3 = data_63_V_read[32'd15];

assign tmp_287_fu_3960_p3 = data_63_V_read[32'd15];

assign tmp_288_fu_3974_p3 = {{xor_ln1495_94_fu_3968_p2}, {10'd0}};

assign tmp_97_fu_544_p3 = data_0_V_read[32'd15];

assign tmp_98_fu_558_p3 = data_0_V_read[32'd15];

assign tmp_99_fu_572_p3 = {{xor_ln1495_fu_566_p2}, {10'd0}};

assign xor_ln1495_32_fu_620_p2 = (tmp_101_fu_612_p3 ^ 1'd1);

assign xor_ln1495_33_fu_674_p2 = (tmp_104_fu_666_p3 ^ 1'd1);

assign xor_ln1495_34_fu_728_p2 = (tmp_107_fu_720_p3 ^ 1'd1);

assign xor_ln1495_35_fu_782_p2 = (tmp_110_fu_774_p3 ^ 1'd1);

assign xor_ln1495_36_fu_836_p2 = (tmp_113_fu_828_p3 ^ 1'd1);

assign xor_ln1495_37_fu_890_p2 = (tmp_116_fu_882_p3 ^ 1'd1);

assign xor_ln1495_38_fu_944_p2 = (tmp_119_fu_936_p3 ^ 1'd1);

assign xor_ln1495_39_fu_998_p2 = (tmp_122_fu_990_p3 ^ 1'd1);

assign xor_ln1495_40_fu_1052_p2 = (tmp_125_fu_1044_p3 ^ 1'd1);

assign xor_ln1495_41_fu_1106_p2 = (tmp_128_fu_1098_p3 ^ 1'd1);

assign xor_ln1495_42_fu_1160_p2 = (tmp_131_fu_1152_p3 ^ 1'd1);

assign xor_ln1495_43_fu_1214_p2 = (tmp_134_fu_1206_p3 ^ 1'd1);

assign xor_ln1495_44_fu_1268_p2 = (tmp_137_fu_1260_p3 ^ 1'd1);

assign xor_ln1495_45_fu_1322_p2 = (tmp_140_fu_1314_p3 ^ 1'd1);

assign xor_ln1495_46_fu_1376_p2 = (tmp_143_fu_1368_p3 ^ 1'd1);

assign xor_ln1495_47_fu_1430_p2 = (tmp_146_fu_1422_p3 ^ 1'd1);

assign xor_ln1495_48_fu_1484_p2 = (tmp_149_fu_1476_p3 ^ 1'd1);

assign xor_ln1495_49_fu_1538_p2 = (tmp_152_fu_1530_p3 ^ 1'd1);

assign xor_ln1495_50_fu_1592_p2 = (tmp_155_fu_1584_p3 ^ 1'd1);

assign xor_ln1495_51_fu_1646_p2 = (tmp_158_fu_1638_p3 ^ 1'd1);

assign xor_ln1495_52_fu_1700_p2 = (tmp_161_fu_1692_p3 ^ 1'd1);

assign xor_ln1495_53_fu_1754_p2 = (tmp_164_fu_1746_p3 ^ 1'd1);

assign xor_ln1495_54_fu_1808_p2 = (tmp_167_fu_1800_p3 ^ 1'd1);

assign xor_ln1495_55_fu_1862_p2 = (tmp_170_fu_1854_p3 ^ 1'd1);

assign xor_ln1495_56_fu_1916_p2 = (tmp_173_fu_1908_p3 ^ 1'd1);

assign xor_ln1495_57_fu_1970_p2 = (tmp_176_fu_1962_p3 ^ 1'd1);

assign xor_ln1495_58_fu_2024_p2 = (tmp_179_fu_2016_p3 ^ 1'd1);

assign xor_ln1495_59_fu_2078_p2 = (tmp_182_fu_2070_p3 ^ 1'd1);

assign xor_ln1495_60_fu_2132_p2 = (tmp_185_fu_2124_p3 ^ 1'd1);

assign xor_ln1495_61_fu_2186_p2 = (tmp_188_fu_2178_p3 ^ 1'd1);

assign xor_ln1495_62_fu_2240_p2 = (tmp_191_fu_2232_p3 ^ 1'd1);

assign xor_ln1495_63_fu_2294_p2 = (tmp_194_fu_2286_p3 ^ 1'd1);

assign xor_ln1495_64_fu_2348_p2 = (tmp_197_fu_2340_p3 ^ 1'd1);

assign xor_ln1495_65_fu_2402_p2 = (tmp_200_fu_2394_p3 ^ 1'd1);

assign xor_ln1495_66_fu_2456_p2 = (tmp_203_fu_2448_p3 ^ 1'd1);

assign xor_ln1495_67_fu_2510_p2 = (tmp_206_fu_2502_p3 ^ 1'd1);

assign xor_ln1495_68_fu_2564_p2 = (tmp_209_fu_2556_p3 ^ 1'd1);

assign xor_ln1495_69_fu_2618_p2 = (tmp_212_fu_2610_p3 ^ 1'd1);

assign xor_ln1495_70_fu_2672_p2 = (tmp_215_fu_2664_p3 ^ 1'd1);

assign xor_ln1495_71_fu_2726_p2 = (tmp_218_fu_2718_p3 ^ 1'd1);

assign xor_ln1495_72_fu_2780_p2 = (tmp_221_fu_2772_p3 ^ 1'd1);

assign xor_ln1495_73_fu_2834_p2 = (tmp_224_fu_2826_p3 ^ 1'd1);

assign xor_ln1495_74_fu_2888_p2 = (tmp_227_fu_2880_p3 ^ 1'd1);

assign xor_ln1495_75_fu_2942_p2 = (tmp_230_fu_2934_p3 ^ 1'd1);

assign xor_ln1495_76_fu_2996_p2 = (tmp_233_fu_2988_p3 ^ 1'd1);

assign xor_ln1495_77_fu_3050_p2 = (tmp_236_fu_3042_p3 ^ 1'd1);

assign xor_ln1495_78_fu_3104_p2 = (tmp_239_fu_3096_p3 ^ 1'd1);

assign xor_ln1495_79_fu_3158_p2 = (tmp_242_fu_3150_p3 ^ 1'd1);

assign xor_ln1495_80_fu_3212_p2 = (tmp_245_fu_3204_p3 ^ 1'd1);

assign xor_ln1495_81_fu_3266_p2 = (tmp_248_fu_3258_p3 ^ 1'd1);

assign xor_ln1495_82_fu_3320_p2 = (tmp_251_fu_3312_p3 ^ 1'd1);

assign xor_ln1495_83_fu_3374_p2 = (tmp_254_fu_3366_p3 ^ 1'd1);

assign xor_ln1495_84_fu_3428_p2 = (tmp_257_fu_3420_p3 ^ 1'd1);

assign xor_ln1495_85_fu_3482_p2 = (tmp_260_fu_3474_p3 ^ 1'd1);

assign xor_ln1495_86_fu_3536_p2 = (tmp_263_fu_3528_p3 ^ 1'd1);

assign xor_ln1495_87_fu_3590_p2 = (tmp_266_fu_3582_p3 ^ 1'd1);

assign xor_ln1495_88_fu_3644_p2 = (tmp_269_fu_3636_p3 ^ 1'd1);

assign xor_ln1495_89_fu_3698_p2 = (tmp_272_fu_3690_p3 ^ 1'd1);

assign xor_ln1495_90_fu_3752_p2 = (tmp_275_fu_3744_p3 ^ 1'd1);

assign xor_ln1495_91_fu_3806_p2 = (tmp_278_fu_3798_p3 ^ 1'd1);

assign xor_ln1495_92_fu_3860_p2 = (tmp_281_fu_3852_p3 ^ 1'd1);

assign xor_ln1495_93_fu_3914_p2 = (tmp_284_fu_3906_p3 ^ 1'd1);

assign xor_ln1495_94_fu_3968_p2 = (tmp_287_fu_3960_p3 ^ 1'd1);

assign xor_ln1495_fu_566_p2 = (tmp_98_fu_558_p3 ^ 1'd1);

assign zext_ln1495_32_fu_634_p1 = tmp_102_fu_626_p3;

assign zext_ln1495_33_fu_688_p1 = tmp_105_fu_680_p3;

assign zext_ln1495_34_fu_742_p1 = tmp_108_fu_734_p3;

assign zext_ln1495_35_fu_796_p1 = tmp_111_fu_788_p3;

assign zext_ln1495_36_fu_850_p1 = tmp_114_fu_842_p3;

assign zext_ln1495_37_fu_904_p1 = tmp_117_fu_896_p3;

assign zext_ln1495_38_fu_958_p1 = tmp_120_fu_950_p3;

assign zext_ln1495_39_fu_1012_p1 = tmp_123_fu_1004_p3;

assign zext_ln1495_40_fu_1066_p1 = tmp_126_fu_1058_p3;

assign zext_ln1495_41_fu_1120_p1 = tmp_129_fu_1112_p3;

assign zext_ln1495_42_fu_1174_p1 = tmp_132_fu_1166_p3;

assign zext_ln1495_43_fu_1228_p1 = tmp_135_fu_1220_p3;

assign zext_ln1495_44_fu_1282_p1 = tmp_138_fu_1274_p3;

assign zext_ln1495_45_fu_1336_p1 = tmp_141_fu_1328_p3;

assign zext_ln1495_46_fu_1390_p1 = tmp_144_fu_1382_p3;

assign zext_ln1495_47_fu_1444_p1 = tmp_147_fu_1436_p3;

assign zext_ln1495_48_fu_1498_p1 = tmp_150_fu_1490_p3;

assign zext_ln1495_49_fu_1552_p1 = tmp_153_fu_1544_p3;

assign zext_ln1495_50_fu_1606_p1 = tmp_156_fu_1598_p3;

assign zext_ln1495_51_fu_1660_p1 = tmp_159_fu_1652_p3;

assign zext_ln1495_52_fu_1714_p1 = tmp_162_fu_1706_p3;

assign zext_ln1495_53_fu_1768_p1 = tmp_165_fu_1760_p3;

assign zext_ln1495_54_fu_1822_p1 = tmp_168_fu_1814_p3;

assign zext_ln1495_55_fu_1876_p1 = tmp_171_fu_1868_p3;

assign zext_ln1495_56_fu_1930_p1 = tmp_174_fu_1922_p3;

assign zext_ln1495_57_fu_1984_p1 = tmp_177_fu_1976_p3;

assign zext_ln1495_58_fu_2038_p1 = tmp_180_fu_2030_p3;

assign zext_ln1495_59_fu_2092_p1 = tmp_183_fu_2084_p3;

assign zext_ln1495_60_fu_2146_p1 = tmp_186_fu_2138_p3;

assign zext_ln1495_61_fu_2200_p1 = tmp_189_fu_2192_p3;

assign zext_ln1495_62_fu_2254_p1 = tmp_192_fu_2246_p3;

assign zext_ln1495_63_fu_2308_p1 = tmp_195_fu_2300_p3;

assign zext_ln1495_64_fu_2362_p1 = tmp_198_fu_2354_p3;

assign zext_ln1495_65_fu_2416_p1 = tmp_201_fu_2408_p3;

assign zext_ln1495_66_fu_2470_p1 = tmp_204_fu_2462_p3;

assign zext_ln1495_67_fu_2524_p1 = tmp_207_fu_2516_p3;

assign zext_ln1495_68_fu_2578_p1 = tmp_210_fu_2570_p3;

assign zext_ln1495_69_fu_2632_p1 = tmp_213_fu_2624_p3;

assign zext_ln1495_70_fu_2686_p1 = tmp_216_fu_2678_p3;

assign zext_ln1495_71_fu_2740_p1 = tmp_219_fu_2732_p3;

assign zext_ln1495_72_fu_2794_p1 = tmp_222_fu_2786_p3;

assign zext_ln1495_73_fu_2848_p1 = tmp_225_fu_2840_p3;

assign zext_ln1495_74_fu_2902_p1 = tmp_228_fu_2894_p3;

assign zext_ln1495_75_fu_2956_p1 = tmp_231_fu_2948_p3;

assign zext_ln1495_76_fu_3010_p1 = tmp_234_fu_3002_p3;

assign zext_ln1495_77_fu_3064_p1 = tmp_237_fu_3056_p3;

assign zext_ln1495_78_fu_3118_p1 = tmp_240_fu_3110_p3;

assign zext_ln1495_79_fu_3172_p1 = tmp_243_fu_3164_p3;

assign zext_ln1495_80_fu_3226_p1 = tmp_246_fu_3218_p3;

assign zext_ln1495_81_fu_3280_p1 = tmp_249_fu_3272_p3;

assign zext_ln1495_82_fu_3334_p1 = tmp_252_fu_3326_p3;

assign zext_ln1495_83_fu_3388_p1 = tmp_255_fu_3380_p3;

assign zext_ln1495_84_fu_3442_p1 = tmp_258_fu_3434_p3;

assign zext_ln1495_85_fu_3496_p1 = tmp_261_fu_3488_p3;

assign zext_ln1495_86_fu_3550_p1 = tmp_264_fu_3542_p3;

assign zext_ln1495_87_fu_3604_p1 = tmp_267_fu_3596_p3;

assign zext_ln1495_88_fu_3658_p1 = tmp_270_fu_3650_p3;

assign zext_ln1495_89_fu_3712_p1 = tmp_273_fu_3704_p3;

assign zext_ln1495_90_fu_3766_p1 = tmp_276_fu_3758_p3;

assign zext_ln1495_91_fu_3820_p1 = tmp_279_fu_3812_p3;

assign zext_ln1495_92_fu_3874_p1 = tmp_282_fu_3866_p3;

assign zext_ln1495_93_fu_3928_p1 = tmp_285_fu_3920_p3;

assign zext_ln1495_94_fu_3982_p1 = tmp_288_fu_3974_p3;

assign zext_ln1495_fu_580_p1 = tmp_99_fu_572_p3;

endmodule //relu_max_ap_fixed_ap_fixed_1_relu1_config5_s
