//////////////////////////////////////////////////////////////////////////////
// HLS generated design for Tiny Darknet neural network (https://pjreddie.com/darknet/tiny-darknet/)
// IEEE FP16 is used.
// Pairs of layers are fused. Separate buffers for weights of each layer. Double buffering for activations. 
//////////////////////////////////////////////////////////////////////////////

// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

//////////////////////////////////////////////////////////////////////////////
// Abridged for VTR by: Daniel Rauch
//////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ps 

module td_fused_top_Block_entry_proc_proc392 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        tmp,
        ap_return
);

parameter    ap_ST_fsm_state1 = 1'd1;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
input  [15:0] tmp;
output  [15:0] ap_return;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg[15:0] ap_return;

reg    ap_done_reg;
  reg   [0:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    ap_block_state1;
reg   [15:0] ap_return_preg;
reg   [0:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 1'd1;
#0 ap_return_preg = 16'd0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_return_preg <= 16'd0;
    end else begin
        if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_return_preg <= tmp;
        end
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_return = tmp;
    end else begin
        ap_return = ap_return_preg;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (ap_done_reg == 1'b1));
end

endmodule //td_fused_top_Block_entry_proc_proc392
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_Block_entry_proc_proc397 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        tmp,
        ap_return
);

parameter    ap_ST_fsm_state1 = 1'd1;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
input  [15:0] tmp;
output  [15:0] ap_return;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg[15:0] ap_return;

reg    ap_done_reg;
  reg   [0:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    ap_block_state1;
reg   [15:0] ap_return_preg;
reg   [0:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 1'd1;
#0 ap_return_preg = 16'd0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_return_preg <= 16'd0;
    end else begin
        if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_return_preg <= tmp;
        end
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_return = tmp;
    end else begin
        ap_return = ap_return_preg;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (ap_done_reg == 1'b1));
end

endmodule //td_fused_top_Block_entry_proc_proc397
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_Block_entry_proc_proc403 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        tmp,
        ap_return
);

parameter    ap_ST_fsm_state1 = 1'd1;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
input  [15:0] tmp;
output  [15:0] ap_return;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg[15:0] ap_return;

reg    ap_done_reg;
  reg   [0:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    ap_block_state1;
reg   [15:0] ap_return_preg;
reg   [0:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 1'd1;
#0 ap_return_preg = 16'd0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_return_preg <= 16'd0;
    end else begin
        if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_return_preg <= tmp;
        end
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_return = tmp;
    end else begin
        ap_return = ap_return_preg;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (ap_done_reg == 1'b1));
end

endmodule //td_fused_top_Block_entry_proc_proc403
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_Block_entry_proc_proc408 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        tmp,
        ap_return
);

parameter    ap_ST_fsm_state1 = 1'd1;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
input  [15:0] tmp;
output  [15:0] ap_return;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg[15:0] ap_return;

reg    ap_done_reg;
  reg   [0:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    ap_block_state1;
reg   [15:0] ap_return_preg;
reg   [0:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 1'd1;
#0 ap_return_preg = 16'd0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_return_preg <= 16'd0;
    end else begin
        if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_return_preg <= tmp;
        end
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_return = tmp;
    end else begin
        ap_return = ap_return_preg;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (ap_done_reg == 1'b1));
end

endmodule //td_fused_top_Block_entry_proc_proc408
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_Block_entry_proc_proc413 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        tmp,
        ap_return
);

parameter    ap_ST_fsm_state1 = 1'd1;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
input  [15:0] tmp;
output  [15:0] ap_return;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg[15:0] ap_return;

reg    ap_done_reg;
  reg   [0:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    ap_block_state1;
reg   [15:0] ap_return_preg;
reg   [0:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 1'd1;
#0 ap_return_preg = 16'd0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_return_preg <= 16'd0;
    end else begin
        if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_return_preg <= tmp;
        end
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_return = tmp;
    end else begin
        ap_return = ap_return_preg;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (ap_done_reg == 1'b1));
end

endmodule //td_fused_top_Block_entry_proc_proc413
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_Block_entry_proc_proc419 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        tmp,
        ap_return
);

parameter    ap_ST_fsm_state1 = 1'd1;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
input  [15:0] tmp;
output  [15:0] ap_return;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg[15:0] ap_return;

reg    ap_done_reg;
  reg   [0:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    ap_block_state1;
reg   [15:0] ap_return_preg;
reg   [0:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 1'd1;
#0 ap_return_preg = 16'd0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_return_preg <= 16'd0;
    end else begin
        if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_return_preg <= tmp;
        end
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_return = tmp;
    end else begin
        ap_return = ap_return_preg;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (ap_done_reg == 1'b1));
end

endmodule //td_fused_top_Block_entry_proc_proc419
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_Block_entry_proc_proc424 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        tmp,
        ap_return
);

parameter    ap_ST_fsm_state1 = 1'd1;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
input  [15:0] tmp;
output  [15:0] ap_return;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg[15:0] ap_return;

reg    ap_done_reg;
  reg   [0:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    ap_block_state1;
reg   [15:0] ap_return_preg;
reg   [0:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 1'd1;
#0 ap_return_preg = 16'd0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_return_preg <= 16'd0;
    end else begin
        if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_return_preg <= tmp;
        end
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_return = tmp;
    end else begin
        ap_return = ap_return_preg;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (ap_done_reg == 1'b1));
end

endmodule //td_fused_top_Block_entry_proc_proc424
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_Block_entry_proc_proc429 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        tmp,
        ap_return
);

parameter    ap_ST_fsm_state1 = 1'd1;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
input  [15:0] tmp;
output  [15:0] ap_return;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg[15:0] ap_return;

reg    ap_done_reg;
  reg   [0:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    ap_block_state1;
reg   [15:0] ap_return_preg;
reg   [0:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 1'd1;
#0 ap_return_preg = 16'd0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_return_preg <= 16'd0;
    end else begin
        if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_return_preg <= tmp;
        end
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_return = tmp;
    end else begin
        ap_return = ap_return_preg;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (ap_done_reg == 1'b1));
end

endmodule //td_fused_top_Block_entry_proc_proc429
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_Block_entry_proc_proc435 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        tmp,
        ap_return
);

parameter    ap_ST_fsm_state1 = 1'd1;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
input  [15:0] tmp;
output  [15:0] ap_return;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg[15:0] ap_return;

reg    ap_done_reg;
  reg   [0:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    ap_block_state1;
reg   [15:0] ap_return_preg;
reg   [0:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 1'd1;
#0 ap_return_preg = 16'd0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_return_preg <= 16'd0;
    end else begin
        if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_return_preg <= tmp;
        end
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_return = tmp;
    end else begin
        ap_return = ap_return_preg;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (ap_done_reg == 1'b1));
end

endmodule //td_fused_top_Block_entry_proc_proc435
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_Block_entry_proc_proc441 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        tmp,
        ap_return
);

parameter    ap_ST_fsm_state1 = 1'd1;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
input  [15:0] tmp;
output  [15:0] ap_return;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg[15:0] ap_return;

reg    ap_done_reg;
  reg   [0:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    ap_block_state1;
reg   [15:0] ap_return_preg;
reg   [0:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 1'd1;
#0 ap_return_preg = 16'd0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_return_preg <= 16'd0;
    end else begin
        if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_return_preg <= tmp;
        end
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_return = tmp;
    end else begin
        ap_return = ap_return_preg;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (ap_done_reg == 1'b1));
end

endmodule //td_fused_top_Block_entry_proc_proc441
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_Block_entry_proc_proc446 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        tmp,
        ap_return
);

parameter    ap_ST_fsm_state1 = 1'd1;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
input  [15:0] tmp;
output  [15:0] ap_return;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg[15:0] ap_return;

reg    ap_done_reg;
  reg   [0:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    ap_block_state1;
reg   [15:0] ap_return_preg;
reg   [0:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 1'd1;
#0 ap_return_preg = 16'd0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_return_preg <= 16'd0;
    end else begin
        if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_return_preg <= tmp;
        end
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_return = tmp;
    end else begin
        ap_return = ap_return_preg;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (ap_done_reg == 1'b1));
end

endmodule //td_fused_top_Block_entry_proc_proc446
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_Block_entry_proc_proc (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        tmp,
        ap_return
);

parameter    ap_ST_fsm_state1 = 1'd1;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
input  [15:0] tmp;
output  [15:0] ap_return;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg[15:0] ap_return;

reg    ap_done_reg;
  reg   [0:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    ap_block_state1;
reg   [15:0] ap_return_preg;
reg   [0:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 1'd1;
#0 ap_return_preg = 16'd0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_return_preg <= 16'd0;
    end else begin
        if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_return_preg <= tmp;
        end
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_return = tmp;
    end else begin
        ap_return = ap_return_preg;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (ap_done_reg == 1'b1));
end

endmodule //td_fused_top_Block_entry_proc_proc
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37360_accum1_out_0_memcore_ram (addr0, ce0, d0, we0, q0, addr1, ce1, d1, we1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 3;
parameter MEM_SIZE = 8;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
input clk;

reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];




always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1) 
            ram[addr1] <= d1; 
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37360_accum1_out_0_memcore(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    q0,
    address1,
    ce1,
    we1,
    d1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd8;
parameter AddressWidth = 32'd3;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;



td_fused_top_dataflow_in_loop_TOP_LOOP37360_accum1_out_0_memcore_ram td_fused_top_dataflow_in_loop_TOP_LOOP37360_accum1_out_0_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_dataflow_in_loop_TOP_LOOP37360_accum1_out_0
#(parameter
    DataWidth    = 16,
    AddressRange = 32,
    AddressWidth = 3,
    BufferCount  = 2,
    MemLatency   = 1,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire                    i_we0,
    input  wire [AddressWidth-1:0] i_address0,
    input  wire [DataWidth-1:0]    i_d0,
    output wire [DataWidth-1:0]    i_q0,
    input  wire                    i_ce1,
    input  wire                    i_we1,
    input  wire [AddressWidth-1:0] i_address1,
    input  wire [DataWidth-1:0]    i_d1,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire                    t_we0,
    input  wire [AddressWidth-1:0] t_address0,
    input  wire [DataWidth-1:0]    t_d0,
    output wire [DataWidth-1:0]    t_q0,
    input  wire                    t_ce1,
    input  wire                    t_we1,
    input  wire [AddressWidth-1:0] t_address1,
    input  wire [DataWidth-1:0]    t_d1
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth-1:0]   prev_iptr    = 1'b0; // previous initiator index
reg  [IndexWidth-1:0]   prev_tptr    = 1'b0; // previous target index
reg  [DataWidth-1:0]    reg_q0      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid0    = 1'b0; // buffer has valid data
reg  [DataWidth-1:0]    reg_q1      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid1    = 1'b0; // buffer has valid data
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
// buffer signals
wire [BufferCount-1:0] buf_ce0;
wire [BufferCount-1:0] buf_we0;
wire [AddressWidth-1:0] buf_a0_0, buf_a0_1;
wire [DataWidth-1:0] buf_d0_0, buf_d0_1;
wire [DataWidth-1:0] buf_q0_0, buf_q0_1;
wire [BufferCount-1:0] buf_ce1;
wire [BufferCount-1:0] buf_we1;
wire [AddressWidth-1:0] buf_a1_0, buf_a1_1;
wire [DataWidth-1:0] buf_d1_0, buf_d1_1;
//------------------------Instantiation------------------
//genvar i;
        td_fused_top_dataflow_in_loop_TOP_LOOP37360_accum1_out_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP37360_accum1_out_0_memcore_U_0 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_0 ),
            .ce0      ( buf_ce0[ 0 ] ),
            .we0      ( buf_we0[ 0 ] ),
            .d0       ( buf_d0_0 ),
            .q0       ( buf_q0_0 ),
            .address1 ( buf_a1_0 ),
            .ce1      ( buf_ce1[ 0 ] ),
            .we1      ( buf_we1[ 0 ] ),
            .d1       ( buf_d1_0 )
        );
        td_fused_top_dataflow_in_loop_TOP_LOOP37360_accum1_out_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP37360_accum1_out_0_memcore_U_1 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_1 ),
            .ce0      ( buf_ce0[ 1 ] ),
            .we0      ( buf_we0[ 1 ] ),
            .d0       ( buf_d0_1 ),
            .q0       ( buf_q0_1 ),
            .address1 ( buf_a1_1 ),
            .ce1      ( buf_ce1[ 1 ] ),
            .we1      ( buf_we1[ 1 ] ),
            .d1       ( buf_d1_1 )
        );

//++++++++++++++++++++++++buffer signals+++++++++++++++++
        assign buf_ce0[ 0 ] = (tptr ==  0  && empty_n) ? t_ce0
                             : (iptr ==  0 ) ? i_ce0 : 1'b0;
        assign buf_a0_0  = (tptr ==  0  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 0 ] = (tptr ==  0  && empty_n)  ? t_we0
                             : (iptr ==  0 ) ? i_we0 : 1'b0;
        assign buf_d0_0  = (tptr ==  0  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 0 ] = (tptr ==  0  && empty_n) ? t_ce1
                             : (iptr ==  0 ) ? i_ce1 : 1'b0;
        assign buf_a1_0  = (tptr ==  0  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 0 ] = (tptr ==  0  && empty_n)  ? t_we1
                             : (iptr ==  0 ) ? i_we1 : 1'b0;
        assign buf_d1_0  = (tptr ==  0  && empty_n) ? t_d1       : i_d1;
        assign buf_ce0[ 1 ] = (tptr ==  1  && empty_n) ? t_ce0
                             : (iptr ==  1 ) ? i_ce0 : 1'b0;
        assign buf_a0_1  = (tptr ==  1  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 1 ] = (tptr ==  1  && empty_n)  ? t_we0
                             : (iptr ==  1 ) ? i_we0 : 1'b0;
        assign buf_d0_1  = (tptr ==  1  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 1 ] = (tptr ==  1  && empty_n) ? t_ce1
                             : (iptr ==  1 ) ? i_ce1 : 1'b0;
        assign buf_a1_1  = (tptr ==  1  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 1 ] = (tptr ==  1  && empty_n)  ? t_we1
                             : (iptr ==  1 ) ? i_we1 : 1'b0;
        assign buf_d1_1  = (tptr ==  1  && empty_n) ? t_d1       : i_d1;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//------------------------Body---------------------------
assign i_q0      = (prev_iptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign t_q0      = reg_valid0 ? reg_q0 : (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// prev_iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_iptr <= 1'b0;
    else begin
        prev_iptr <= iptr;
    end
end

// prev_tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_tptr <= 1'b0;
    else begin
        prev_tptr <= tptr;
    end
end

// reg_q0 and reg_valid0
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q0     <= 1'b0;
        reg_valid0 <= 1'b0;
    end else if (!t_ce0 && !reg_valid0) begin
        reg_q0     <= (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
        reg_valid0 <= 1'b1;
    end else if (t_ce0) begin
        reg_valid0 <= 1'b0;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37360_ifmap_vec_0_0_memcore_ram (addr0, ce0, d0, we0, q0, addr1, ce1, d1, we1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 8;
parameter MEM_SIZE = 256;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
input clk;

reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];




always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1) 
            ram[addr1] <= d1; 
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37360_ifmap_vec_0_0_memcore(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    q0,
    address1,
    ce1,
    we1,
    d1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd256;
parameter AddressWidth = 32'd8;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;



td_fused_top_dataflow_in_loop_TOP_LOOP37360_ifmap_vec_0_0_memcore_ram td_fused_top_dataflow_in_loop_TOP_LOOP37360_ifmap_vec_0_0_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_dataflow_in_loop_TOP_LOOP37360_ifmap_vec_0_0
#(parameter
    DataWidth    = 16,
    AddressRange = 32,
    AddressWidth = 8,
    BufferCount  = 2,
    MemLatency   = 1,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire                    i_we0,
    input  wire [AddressWidth-1:0] i_address0,
    input  wire [DataWidth-1:0]    i_d0,
    output wire [DataWidth-1:0]    i_q0,
    input  wire                    i_ce1,
    input  wire                    i_we1,
    input  wire [AddressWidth-1:0] i_address1,
    input  wire [DataWidth-1:0]    i_d1,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire                    t_we0,
    input  wire [AddressWidth-1:0] t_address0,
    input  wire [DataWidth-1:0]    t_d0,
    output wire [DataWidth-1:0]    t_q0,
    input  wire                    t_ce1,
    input  wire                    t_we1,
    input  wire [AddressWidth-1:0] t_address1,
    input  wire [DataWidth-1:0]    t_d1
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth-1:0]   prev_iptr    = 1'b0; // previous initiator index
reg  [IndexWidth-1:0]   prev_tptr    = 1'b0; // previous target index
reg  [DataWidth-1:0]    reg_q0      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid0    = 1'b0; // buffer has valid data
reg  [DataWidth-1:0]    reg_q1      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid1    = 1'b0; // buffer has valid data
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
// buffer signals
wire [BufferCount-1:0] buf_ce0;
wire [BufferCount-1:0] buf_we0;
wire [AddressWidth-1:0] buf_a0_0, buf_a0_1;
wire [DataWidth-1:0] buf_d0_0, buf_d0_1;
wire [DataWidth-1:0] buf_q0_0, buf_q0_1;
wire [BufferCount-1:0] buf_ce1;
wire [BufferCount-1:0] buf_we1;
wire [AddressWidth-1:0] buf_a1_0, buf_a1_1;
wire [DataWidth-1:0] buf_d1_0, buf_d1_1;
//------------------------Instantiation------------------
//genvar i;
        td_fused_top_dataflow_in_loop_TOP_LOOP37360_ifmap_vec_0_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP37360_ifmap_vec_0_0_memcore_U_0 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_0 ),
            .ce0      ( buf_ce0[ 0 ] ),
            .we0      ( buf_we0[ 0 ] ),
            .d0       ( buf_d0_0 ),
            .q0       ( buf_q0_0 ),
            .address1 ( buf_a1_0 ),
            .ce1      ( buf_ce1[ 0 ] ),
            .we1      ( buf_we1[ 0 ] ),
            .d1       ( buf_d1_0 )
        );
        td_fused_top_dataflow_in_loop_TOP_LOOP37360_ifmap_vec_0_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP37360_ifmap_vec_0_0_memcore_U_1 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_1 ),
            .ce0      ( buf_ce0[ 1 ] ),
            .we0      ( buf_we0[ 1 ] ),
            .d0       ( buf_d0_1 ),
            .q0       ( buf_q0_1 ),
            .address1 ( buf_a1_1 ),
            .ce1      ( buf_ce1[ 1 ] ),
            .we1      ( buf_we1[ 1 ] ),
            .d1       ( buf_d1_1 )
        );

//++++++++++++++++++++++++buffer signals+++++++++++++++++
        assign buf_ce0[ 0 ] = (tptr ==  0  && empty_n) ? t_ce0
                             : (iptr ==  0 ) ? i_ce0 : 1'b0;
        assign buf_a0_0  = (tptr ==  0  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 0 ] = (tptr ==  0  && empty_n)  ? t_we0
                             : (iptr ==  0 ) ? i_we0 : 1'b0;
        assign buf_d0_0  = (tptr ==  0  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 0 ] = (tptr ==  0  && empty_n) ? t_ce1
                             : (iptr ==  0 ) ? i_ce1 : 1'b0;
        assign buf_a1_0  = (tptr ==  0  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 0 ] = (tptr ==  0  && empty_n)  ? t_we1
                             : (iptr ==  0 ) ? i_we1 : 1'b0;
        assign buf_d1_0  = (tptr ==  0  && empty_n) ? t_d1       : i_d1;
        assign buf_ce0[ 1 ] = (tptr ==  1  && empty_n) ? t_ce0
                             : (iptr ==  1 ) ? i_ce0 : 1'b0;
        assign buf_a0_1  = (tptr ==  1  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 1 ] = (tptr ==  1  && empty_n)  ? t_we0
                             : (iptr ==  1 ) ? i_we0 : 1'b0;
        assign buf_d0_1  = (tptr ==  1  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 1 ] = (tptr ==  1  && empty_n) ? t_ce1
                             : (iptr ==  1 ) ? i_ce1 : 1'b0;
        assign buf_a1_1  = (tptr ==  1  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 1 ] = (tptr ==  1  && empty_n)  ? t_we1
                             : (iptr ==  1 ) ? i_we1 : 1'b0;
        assign buf_d1_1  = (tptr ==  1  && empty_n) ? t_d1       : i_d1;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//------------------------Body---------------------------
assign i_q0      = (prev_iptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign t_q0      = reg_valid0 ? reg_q0 : (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// prev_iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_iptr <= 1'b0;
    else begin
        prev_iptr <= iptr;
    end
end

// prev_tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_tptr <= 1'b0;
    else begin
        prev_tptr <= tptr;
    end
end

// reg_q0 and reg_valid0
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q0     <= 1'b0;
        reg_valid0 <= 1'b0;
    end else if (!t_ce0 && !reg_valid0) begin
        reg_q0     <= (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
        reg_valid0 <= 1'b1;
    end else if (t_ce0) begin
        reg_valid0 <= 1'b0;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37360_products_0_memcore_ram (addr0, ce0, d0, we0, q0, addr1, ce1, q1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 8;
parameter MEM_SIZE = 256;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
output reg[DWIDTH-1:0] q1;
input clk;

reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];




always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        q1 <= ram[addr1];
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37360_products_0_memcore(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    q0,
    address1,
    ce1,
    q1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd256;
parameter AddressWidth = 32'd8;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
output[DataWidth - 1:0] q1;



td_fused_top_dataflow_in_loop_TOP_LOOP37360_products_0_memcore_ram td_fused_top_dataflow_in_loop_TOP_LOOP37360_products_0_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .q1( q1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_dataflow_in_loop_TOP_LOOP37360_products_0
#(parameter
    DataWidth    = 16,
    AddressRange = 32,
    AddressWidth = 8,
    BufferCount  = 2,
    MemLatency   = 1,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire                    i_we0,
    input  wire [AddressWidth-1:0] i_address0,
    input  wire [DataWidth-1:0]    i_d0,
    output wire [DataWidth-1:0]    i_q0,
    input  wire                    i_ce1,
    input  wire [AddressWidth-1:0] i_address1,
    output wire [DataWidth-1:0]    i_q1,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire                    t_we0,
    input  wire [AddressWidth-1:0] t_address0,
    input  wire [DataWidth-1:0]    t_d0,
    output wire [DataWidth-1:0]    t_q0,
    input  wire                    t_ce1,
    input  wire [AddressWidth-1:0] t_address1,
    output wire [DataWidth-1:0]    t_q1
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth-1:0]   prev_iptr    = 1'b0; // previous initiator index
reg  [IndexWidth-1:0]   prev_tptr    = 1'b0; // previous target index
reg  [DataWidth-1:0]    reg_q0      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid0    = 1'b0; // buffer has valid data
reg  [DataWidth-1:0]    reg_q1      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid1    = 1'b0; // buffer has valid data
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
// buffer signals
wire [BufferCount-1:0] buf_ce0;
wire [BufferCount-1:0] buf_we0;
wire [AddressWidth-1:0] buf_a0_0, buf_a0_1;
wire [DataWidth-1:0] buf_d0_0, buf_d0_1;
wire [DataWidth-1:0] buf_q0_0, buf_q0_1;
wire [BufferCount-1:0] buf_ce1;
wire [AddressWidth-1:0] buf_a1_0, buf_a1_1;
wire [DataWidth-1:0] buf_q1_0, buf_q1_1;
//------------------------Instantiation------------------
//genvar i;
        td_fused_top_dataflow_in_loop_TOP_LOOP37360_products_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP37360_products_0_memcore_U_0 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_0 ),
            .ce0      ( buf_ce0[ 0 ] ),
            .we0      ( buf_we0[ 0 ] ),
            .d0       ( buf_d0_0 ),
            .q0       ( buf_q0_0 ),
            .address1 ( buf_a1_0 ),
            .ce1      ( buf_ce1[ 0 ] ),
            .q1       ( buf_q1_0 )
        );
        td_fused_top_dataflow_in_loop_TOP_LOOP37360_products_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP37360_products_0_memcore_U_1 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_1 ),
            .ce0      ( buf_ce0[ 1 ] ),
            .we0      ( buf_we0[ 1 ] ),
            .d0       ( buf_d0_1 ),
            .q0       ( buf_q0_1 ),
            .address1 ( buf_a1_1 ),
            .ce1      ( buf_ce1[ 1 ] ),
            .q1       ( buf_q1_1 )
        );

//++++++++++++++++++++++++buffer signals+++++++++++++++++
        assign buf_ce0[ 0 ] = (tptr ==  0  && empty_n) ? t_ce0
                             : (iptr ==  0 ) ? i_ce0 : 1'b0;
        assign buf_a0_0  = (tptr ==  0  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 0 ] = (tptr ==  0  && empty_n)  ? t_we0
                             : (iptr ==  0 ) ? i_we0 : 1'b0;
        assign buf_d0_0  = (tptr ==  0  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 0 ] = (tptr ==  0  && empty_n) ? t_ce1
                             : (iptr ==  0 ) ? i_ce1 : 1'b0;
        assign buf_a1_0  = (tptr ==  0  && empty_n) ?  t_address1 : i_address1;
        assign buf_ce0[ 1 ] = (tptr ==  1  && empty_n) ? t_ce0
                             : (iptr ==  1 ) ? i_ce0 : 1'b0;
        assign buf_a0_1  = (tptr ==  1  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 1 ] = (tptr ==  1  && empty_n)  ? t_we0
                             : (iptr ==  1 ) ? i_we0 : 1'b0;
        assign buf_d0_1  = (tptr ==  1  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 1 ] = (tptr ==  1  && empty_n) ? t_ce1
                             : (iptr ==  1 ) ? i_ce1 : 1'b0;
        assign buf_a1_1  = (tptr ==  1  && empty_n) ?  t_address1 : i_address1;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//------------------------Body---------------------------
assign i_q0      = (prev_iptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign t_q0      = reg_valid0 ? reg_q0 : (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign i_q1      = (prev_iptr == 1'b1 ? buf_q1_1 : buf_q1_0);
assign t_q1      = reg_valid1 ? reg_q1 : (prev_tptr == 1'b1 ? buf_q1_1 : buf_q1_0);

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// prev_iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_iptr <= 1'b0;
    else begin
        prev_iptr <= iptr;
    end
end

// prev_tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_tptr <= 1'b0;
    else begin
        prev_tptr <= tptr;
    end
end

// reg_q0 and reg_valid0
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q0     <= 1'b0;
        reg_valid0 <= 1'b0;
    end else if (!t_ce0 && !reg_valid0) begin
        reg_q0     <= (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
        reg_valid0 <= 1'b1;
    end else if (t_ce0) begin
        reg_valid0 <= 1'b0;
    end
end

// reg_q1 and reg_valid1
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q1     <= 1'b0;
        reg_valid1 <= 1'b0;
    end else if (!t_ce1 && !reg_valid1) begin
        reg_q1     <= (prev_tptr == 1'b1 ? buf_q1_1 : buf_q1_0);
        reg_valid1 <= 1'b1;
    end else if (t_ce1) begin
        reg_valid1 <= 1'b0;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_dataflow_in_loop_TOP_LOOP37360 (
        ap_clk,
        ap_rst,
        in_data_address0,
        in_data_ce0,
        in_data_d0,
        in_data_q0,
        in_data_we0,
        in_data_address1,
        in_data_ce1,
        in_data_d1,
        in_data_q1,
        in_data_we1,
        filter_data_address0,
        filter_data_ce0,
        filter_data_d0,
        filter_data_q0,
        filter_data_we0,
        filter_data_address1,
        filter_data_ce1,
        filter_data_d1,
        filter_data_q1,
        filter_data_we1,
        adjustments_address0,
        adjustments_ce0,
        adjustments_d0,
        adjustments_q0,
        adjustments_we0,
        adjustments_address1,
        adjustments_ce1,
        adjustments_d1,
        adjustments_q1,
        adjustments_we1,
        out_data_address0,
        out_data_ce0,
        out_data_d0,
        out_data_q0,
        out_data_we0,
        out_data_address1,
        out_data_ce1,
        out_data_d1,
        out_data_q1,
        out_data_we1,
        ap_start,
        in_data_empty_n,
        in_data_read,
        out_data_full_n,
        out_data_write,
        ap_done,
        ap_ready,
        ap_idle,
        ap_continue
);


input   ap_clk;
input   ap_rst;
output  [13:0] in_data_address0;
output   in_data_ce0;
output  [63:0] in_data_d0;
input  [63:0] in_data_q0;
output   in_data_we0;
output  [13:0] in_data_address1;
output   in_data_ce1;
output  [63:0] in_data_d1;
input  [63:0] in_data_q1;
output   in_data_we1;
output  [13:0] filter_data_address0;
output   filter_data_ce0;
output  [15:0] filter_data_d0;
input  [15:0] filter_data_q0;
output   filter_data_we0;
output  [13:0] filter_data_address1;
output   filter_data_ce1;
output  [15:0] filter_data_d1;
input  [15:0] filter_data_q1;
output   filter_data_we1;
output  [5:0] adjustments_address0;
output   adjustments_ce0;
output  [47:0] adjustments_d0;
input  [47:0] adjustments_q0;
output   adjustments_we0;
output  [5:0] adjustments_address1;
output   adjustments_ce1;
output  [47:0] adjustments_d1;
input  [47:0] adjustments_q1;
output   adjustments_we1;
output  [11:0] out_data_address0;
output   out_data_ce0;
output  [63:0] out_data_d0;
input  [63:0] out_data_q0;
output   out_data_we0;
output  [11:0] out_data_address1;
output   out_data_ce1;
output  [63:0] out_data_d1;
input  [63:0] out_data_q1;
output   out_data_we1;
input   ap_start;
input   in_data_empty_n;
output   in_data_read;
input   out_data_full_n;
output   out_data_write;
output   ap_done;
output   ap_ready;
output   ap_idle;
input   ap_continue;

wire   [15:0] ifmap_vec_0_0_i_q0;
wire   [15:0] ifmap_vec_0_0_t_q0;
wire   [15:0] weight_vecs_0_0_0_i_q0;
wire   [15:0] weight_vecs_0_0_0_t_q0;
wire   [15:0] products_0_i_q0;
wire   [15:0] products_0_i_q1;
wire   [15:0] products_0_t_q0;
wire   [15:0] products_0_t_q1;
wire   [15:0] accum1_out_0_i_q0;
wire   [15:0] accum1_out_0_t_q0;
wire    tdf9_get_next_ijk_U0_ap_start;
wire    tdf9_get_next_ijk_U0_ap_done;
wire    tdf9_get_next_ijk_U0_ap_continue;
wire    tdf9_get_next_ijk_U0_ap_idle;
wire    tdf9_get_next_ijk_U0_ap_ready;
wire    tdf9_get_next_ijk_U0_start_out;
wire    tdf9_get_next_ijk_U0_start_write;
wire   [15:0] tdf9_get_next_ijk_U0_indices_0_din;
wire    tdf9_get_next_ijk_U0_indices_0_write;
wire   [15:0] tdf9_get_next_ijk_U0_indices_1_din;
wire    tdf9_get_next_ijk_U0_indices_1_write;
wire   [5:0] tdf9_get_next_ijk_U0_indices_2_out_din;
wire    tdf9_get_next_ijk_U0_indices_2_out_write;
wire   [5:0] tdf9_get_next_ijk_U0_indices_2_out1_din;
wire    tdf9_get_next_ijk_U0_indices_2_out1_write;
wire    tdf9_readInputs_U0_ap_start;
wire    tdf9_readInputs_U0_ap_done;
wire    tdf9_readInputs_U0_ap_continue;
wire    tdf9_readInputs_U0_ap_idle;
wire    tdf9_readInputs_U0_ap_ready;
wire   [13:0] tdf9_readInputs_U0_in_data_address0;
wire    tdf9_readInputs_U0_in_data_ce0;
wire    tdf9_readInputs_U0_indices_01_read;
wire    tdf9_readInputs_U0_indices_12_read;
wire   [7:0] tdf9_readInputs_U0_ifmap_vec_0_0_address0;
wire    tdf9_readInputs_U0_ifmap_vec_0_0_ce0;
wire    tdf9_readInputs_U0_ifmap_vec_0_0_we0;
wire   [15:0] tdf9_readInputs_U0_ifmap_vec_0_0_d0;
wire   [7:0] tdf9_readInputs_U0_ifmap_vec_0_0_address1;
wire    tdf9_readInputs_U0_ifmap_vec_0_0_ce1;
wire    tdf9_readInputs_U0_ifmap_vec_0_0_we1;
wire   [15:0] tdf9_readInputs_U0_ifmap_vec_0_0_d1;
wire   [3:0] tdf9_readInputs_U0_indices_01_out_din;
wire    tdf9_readInputs_U0_indices_01_out_write;
wire   [7:0] tdf9_readInputs_U0_indices_12_out_din;
wire    tdf9_readInputs_U0_indices_12_out_write;
wire    tdf9_readInputs_U0_in_data_full_n;
wire    tdf9_readInputs_U0_in_data_write;
wire    ap_channel_done_ifmap_vec_0_0;
wire    tdf9_readInputs_U0_ifmap_vec_0_0_full_n;
wire    tdf9_readFilters62_U0_ap_start;
wire    tdf9_readFilters62_U0_ap_done;
wire    tdf9_readFilters62_U0_ap_continue;
wire    tdf9_readFilters62_U0_ap_idle;
wire    tdf9_readFilters62_U0_ap_ready;
wire   [13:0] tdf9_readFilters62_U0_filter_data_address0;
wire    tdf9_readFilters62_U0_filter_data_ce0;
wire    tdf9_readFilters62_U0_indices_23_read;
wire   [7:0] tdf9_readFilters62_U0_weight_vecs_0_0_0_address0;
wire    tdf9_readFilters62_U0_weight_vecs_0_0_0_ce0;
wire    tdf9_readFilters62_U0_weight_vecs_0_0_0_we0;
wire   [15:0] tdf9_readFilters62_U0_weight_vecs_0_0_0_d0;
wire    ap_channel_done_weight_vecs_0_0_0;
wire    tdf9_readFilters62_U0_weight_vecs_0_0_0_full_n;
wire    tdf9_dot_product_U0_ap_start;
wire    tdf9_dot_product_U0_ap_done;
wire    tdf9_dot_product_U0_ap_continue;
wire    tdf9_dot_product_U0_ap_idle;
wire    tdf9_dot_product_U0_ap_ready;
wire   [7:0] tdf9_dot_product_U0_ifmap_vec_0_0_address0;
wire    tdf9_dot_product_U0_ifmap_vec_0_0_ce0;
wire   [7:0] tdf9_dot_product_U0_weight_vecs_0_0_0_address0;
wire    tdf9_dot_product_U0_weight_vecs_0_0_0_ce0;
wire   [7:0] tdf9_dot_product_U0_products_0_address0;
wire    tdf9_dot_product_U0_products_0_ce0;
wire    tdf9_dot_product_U0_products_0_we0;
wire   [15:0] tdf9_dot_product_U0_products_0_d0;
wire    ap_channel_done_products_0;
wire    tdf9_dot_product_U0_products_0_full_n;
wire    tdf9_accum_1_U0_ap_start;
wire    tdf9_accum_1_U0_ap_done;
wire    tdf9_accum_1_U0_ap_continue;
wire    tdf9_accum_1_U0_ap_idle;
wire    tdf9_accum_1_U0_ap_ready;
wire   [7:0] tdf9_accum_1_U0_accum_in_0_address0;
wire    tdf9_accum_1_U0_accum_in_0_ce0;
wire   [7:0] tdf9_accum_1_U0_accum_in_0_address1;
wire    tdf9_accum_1_U0_accum_in_0_ce1;
wire   [2:0] tdf9_accum_1_U0_accum_out_address0;
wire    tdf9_accum_1_U0_accum_out_ce0;
wire    tdf9_accum_1_U0_accum_out_we0;
wire   [15:0] tdf9_accum_1_U0_accum_out_d0;
wire   [2:0] tdf9_accum_1_U0_accum_out_address1;
wire    tdf9_accum_1_U0_accum_out_ce1;
wire    tdf9_accum_1_U0_accum_out_we1;
wire   [15:0] tdf9_accum_1_U0_accum_out_d1;
wire    ap_channel_done_accum1_out_0;
wire    tdf9_accum_1_U0_accum_out_full_n;
wire    tdf9_accum_2_U0_ap_start;
wire    tdf9_accum_2_U0_ap_done;
wire    tdf9_accum_2_U0_ap_continue;
wire    tdf9_accum_2_U0_ap_idle;
wire    tdf9_accum_2_U0_ap_ready;
wire   [15:0] tdf9_accum_2_U0_accum_in_2;
wire    tdf9_accum_2_U0_accum_in_2_ap_vld;
wire   [2:0] tdf9_accum_2_U0_accum_in_address0;
wire    tdf9_accum_2_U0_accum_in_ce0;
wire    ap_channel_done_tmp_channel;
wire    tmp_channel_full_n;
wire    Block_entry_proc_proc429_U0_ap_start;
wire    Block_entry_proc_proc429_U0_ap_done;
wire    Block_entry_proc_proc429_U0_ap_continue;
wire    Block_entry_proc_proc429_U0_ap_idle;
wire    Block_entry_proc_proc429_U0_ap_ready;
wire   [15:0] Block_entry_proc_proc429_U0_ap_return;
wire    ap_channel_done_sums_0;
wire    sums_0_full_n;
wire    tdf9_adjust_U0_ap_start;
wire    tdf9_adjust_U0_ap_done;
wire    tdf9_adjust_U0_ap_continue;
wire    tdf9_adjust_U0_ap_idle;
wire    tdf9_adjust_U0_ap_ready;
wire   [5:0] tdf9_adjust_U0_adjustments_address0;
wire    tdf9_adjust_U0_adjustments_ce0;
wire    tdf9_adjust_U0_indices_23_read;
wire   [15:0] tdf9_adjust_U0_ap_return;
wire    ap_channel_done_outputs_0;
wire    outputs_0_full_n;
wire    tdf9_writeOutputs_unaligned_U0_ap_start;
wire    tdf9_writeOutputs_unaligned_U0_ap_done;
wire    tdf9_writeOutputs_unaligned_U0_ap_continue;
wire    tdf9_writeOutputs_unaligned_U0_ap_idle;
wire    tdf9_writeOutputs_unaligned_U0_ap_ready;
wire    tdf9_writeOutputs_unaligned_U0_indices_01_read;
wire    tdf9_writeOutputs_unaligned_U0_indices_12_read;
wire   [11:0] tdf9_writeOutputs_unaligned_U0_out_data_address1;
wire    tdf9_writeOutputs_unaligned_U0_out_data_ce1;
wire    tdf9_writeOutputs_unaligned_U0_out_data_we1;
wire   [63:0] tdf9_writeOutputs_unaligned_U0_out_data_d1;
wire    tdf9_writeOutputs_unaligned_U0_out_data_full_n;
wire    tdf9_writeOutputs_unaligned_U0_out_data_write;
wire    ap_sync_continue;
wire    ifmap_vec_0_0_i_full_n;
wire    ifmap_vec_0_0_t_empty_n;
wire    weight_vecs_0_0_0_i_full_n;
wire    weight_vecs_0_0_0_t_empty_n;
wire    products_0_i_full_n;
wire    products_0_t_empty_n;
wire   [15:0] products_0_t_d1;
wire    products_0_t_we1;
wire    accum1_out_0_i_full_n;
wire    accum1_out_0_t_empty_n;
wire    indices_01_c_full_n;
wire   [15:0] indices_01_c_dout;
wire    indices_01_c_empty_n;
wire    indices_12_c_full_n;
wire   [15:0] indices_12_c_dout;
wire    indices_12_c_empty_n;
wire    indices_23_c_full_n;
wire   [5:0] indices_23_c_dout;
wire    indices_23_c_empty_n;
wire    indices_23_c1_full_n;
wire   [5:0] indices_23_c1_dout;
wire    indices_23_c1_empty_n;
wire    indices_01_c2_full_n;
wire   [3:0] indices_01_c2_dout;
wire    indices_01_c2_empty_n;
wire    indices_12_c3_full_n;
wire   [7:0] indices_12_c3_dout;
wire    indices_12_c3_empty_n;
wire   [15:0] tmp_channel_dout;
wire    tmp_channel_empty_n;
wire   [15:0] sums_0_dout;
wire    sums_0_empty_n;
wire   [15:0] outputs_0_dout;
wire    outputs_0_empty_n;
wire    ap_sync_done;
wire    ap_sync_ready;
reg    ap_sync_reg_tdf9_get_next_ijk_U0_ap_ready;
wire    ap_sync_tdf9_get_next_ijk_U0_ap_ready;
reg    ap_sync_reg_tdf9_readInputs_U0_ap_ready;
wire    ap_sync_tdf9_readInputs_U0_ap_ready;
wire   [0:0] start_for_tdf9_readFilters62_U0_din;
wire    start_for_tdf9_readFilters62_U0_full_n;
wire   [0:0] start_for_tdf9_readFilters62_U0_dout;
wire    start_for_tdf9_readFilters62_U0_empty_n;
wire    tdf9_readInputs_U0_start_full_n;
wire    tdf9_readInputs_U0_start_write;
wire    tdf9_readFilters62_U0_start_full_n;
wire    tdf9_readFilters62_U0_start_write;
wire    tdf9_dot_product_U0_start_full_n;
wire    tdf9_dot_product_U0_start_write;
wire    tdf9_accum_1_U0_start_full_n;
wire    tdf9_accum_1_U0_start_write;
wire    tdf9_accum_2_U0_start_full_n;
wire    tdf9_accum_2_U0_start_write;
wire    Block_entry_proc_proc429_U0_start_full_n;
wire    Block_entry_proc_proc429_U0_start_write;
wire    tdf9_adjust_U0_start_full_n;
wire    tdf9_adjust_U0_start_write;
wire    tdf9_writeOutputs_unaligned_U0_start_full_n;
wire    tdf9_writeOutputs_unaligned_U0_start_write;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_sync_reg_tdf9_get_next_ijk_U0_ap_ready = 1'b0;
#0 ap_sync_reg_tdf9_readInputs_U0_ap_ready = 1'b0;
end

td_fused_top_dataflow_in_loop_TOP_LOOP37360_ifmap_vec_0_0 #(
    .DataWidth( 16 ),
    .AddressRange( 256 ),
    .AddressWidth( 8 ))
ifmap_vec_0_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf9_readInputs_U0_ap_done),
    .i_full_n(ifmap_vec_0_0_i_full_n),
    .i_ce0(tdf9_readInputs_U0_ifmap_vec_0_0_ce0),
    .i_we0(tdf9_readInputs_U0_ifmap_vec_0_0_we0),
    .i_address0(tdf9_readInputs_U0_ifmap_vec_0_0_address0),
    .i_d0(tdf9_readInputs_U0_ifmap_vec_0_0_d0),
    .i_q0(ifmap_vec_0_0_i_q0),
    .i_ce1(tdf9_readInputs_U0_ifmap_vec_0_0_ce1),
    .i_we1(tdf9_readInputs_U0_ifmap_vec_0_0_we1),
    .i_address1(tdf9_readInputs_U0_ifmap_vec_0_0_address1),
    .i_d1(tdf9_readInputs_U0_ifmap_vec_0_0_d1),
    .t_ce(1'b1),
    .t_read(tdf9_dot_product_U0_ap_ready),
    .t_empty_n(ifmap_vec_0_0_t_empty_n),
    .t_ce0(tdf9_dot_product_U0_ifmap_vec_0_0_ce0),
    .t_we0(1'b0),
    .t_address0(tdf9_dot_product_U0_ifmap_vec_0_0_address0),
    .t_d0(16'd0),
    .t_q0(ifmap_vec_0_0_t_q0),
    .t_ce1(1'b0),
    .t_we1(1'b0),
    .t_address1(8'd0),
    .t_d1(16'd0)
);

td_fused_top_dataflow_in_loop_TOP_LOOP37360_weight_vecs_0_0_0 #(
    .DataWidth( 16 ),
    .AddressRange( 256 ),
    .AddressWidth( 8 ))
weight_vecs_0_0_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf9_readFilters62_U0_ap_done),
    .i_full_n(weight_vecs_0_0_0_i_full_n),
    .i_ce0(tdf9_readFilters62_U0_weight_vecs_0_0_0_ce0),
    .i_we0(tdf9_readFilters62_U0_weight_vecs_0_0_0_we0),
    .i_address0(tdf9_readFilters62_U0_weight_vecs_0_0_0_address0),
    .i_d0(tdf9_readFilters62_U0_weight_vecs_0_0_0_d0),
    .i_q0(weight_vecs_0_0_0_i_q0),
    .t_ce(1'b1),
    .t_read(tdf9_dot_product_U0_ap_ready),
    .t_empty_n(weight_vecs_0_0_0_t_empty_n),
    .t_ce0(tdf9_dot_product_U0_weight_vecs_0_0_0_ce0),
    .t_we0(1'b0),
    .t_address0(tdf9_dot_product_U0_weight_vecs_0_0_0_address0),
    .t_d0(16'd0),
    .t_q0(weight_vecs_0_0_0_t_q0)
);

td_fused_top_dataflow_in_loop_TOP_LOOP37360_products_0 #(
    .DataWidth( 16 ),
    .AddressRange( 256 ),
    .AddressWidth( 8 ))
products_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf9_dot_product_U0_ap_done),
    .i_full_n(products_0_i_full_n),
    .i_ce0(tdf9_dot_product_U0_products_0_ce0),
    .i_we0(tdf9_dot_product_U0_products_0_we0),
    .i_address0(tdf9_dot_product_U0_products_0_address0),
    .i_d0(tdf9_dot_product_U0_products_0_d0),
    .i_q0(products_0_i_q0),
    .i_ce1(1'b0),
    .i_address1(8'd0),
    .i_q1(products_0_i_q1),
    .t_ce(1'b1),
    .t_read(tdf9_accum_1_U0_ap_ready),
    .t_empty_n(products_0_t_empty_n),
    .t_ce0(tdf9_accum_1_U0_accum_in_0_ce0),
    .t_we0(1'b0),
    .t_address0(tdf9_accum_1_U0_accum_in_0_address0),
    .t_d0(16'd0),
    .t_q0(products_0_t_q0),
    .t_ce1(tdf9_accum_1_U0_accum_in_0_ce1),
    .t_address1(tdf9_accum_1_U0_accum_in_0_address1),
    .t_q1(products_0_t_q1)
);

td_fused_top_dataflow_in_loop_TOP_LOOP37360_accum1_out_0 #(
    .DataWidth( 16 ),
    .AddressRange( 8 ),
    .AddressWidth( 3 ))
accum1_out_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf9_accum_1_U0_ap_done),
    .i_full_n(accum1_out_0_i_full_n),
    .i_ce0(tdf9_accum_1_U0_accum_out_ce0),
    .i_we0(tdf9_accum_1_U0_accum_out_we0),
    .i_address0(tdf9_accum_1_U0_accum_out_address0),
    .i_d0(tdf9_accum_1_U0_accum_out_d0),
    .i_q0(accum1_out_0_i_q0),
    .i_ce1(tdf9_accum_1_U0_accum_out_ce1),
    .i_we1(tdf9_accum_1_U0_accum_out_we1),
    .i_address1(tdf9_accum_1_U0_accum_out_address1),
    .i_d1(tdf9_accum_1_U0_accum_out_d1),
    .t_ce(1'b1),
    .t_read(tdf9_accum_2_U0_ap_ready),
    .t_empty_n(accum1_out_0_t_empty_n),
    .t_ce0(tdf9_accum_2_U0_accum_in_ce0),
    .t_we0(1'b0),
    .t_address0(tdf9_accum_2_U0_accum_in_address0),
    .t_d0(16'd0),
    .t_q0(accum1_out_0_t_q0),
    .t_ce1(1'b0),
    .t_we1(1'b0),
    .t_address1(3'd0),
    .t_d1(16'd0)
);

td_fused_top_tdf9_get_next_ijk tdf9_get_next_ijk_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf9_get_next_ijk_U0_ap_start),
    .start_full_n(start_for_tdf9_readFilters62_U0_full_n),
    .ap_done(tdf9_get_next_ijk_U0_ap_done),
    .ap_continue(tdf9_get_next_ijk_U0_ap_continue),
    .ap_idle(tdf9_get_next_ijk_U0_ap_idle),
    .ap_ready(tdf9_get_next_ijk_U0_ap_ready),
    .start_out(tdf9_get_next_ijk_U0_start_out),
    .start_write(tdf9_get_next_ijk_U0_start_write),
    .indices_0_din(tdf9_get_next_ijk_U0_indices_0_din),
    .indices_0_full_n(indices_01_c_full_n),
    .indices_0_write(tdf9_get_next_ijk_U0_indices_0_write),
    .indices_1_din(tdf9_get_next_ijk_U0_indices_1_din),
    .indices_1_full_n(indices_12_c_full_n),
    .indices_1_write(tdf9_get_next_ijk_U0_indices_1_write),
    .indices_2_out_din(tdf9_get_next_ijk_U0_indices_2_out_din),
    .indices_2_out_full_n(indices_23_c_full_n),
    .indices_2_out_write(tdf9_get_next_ijk_U0_indices_2_out_write),
    .indices_2_out1_din(tdf9_get_next_ijk_U0_indices_2_out1_din),
    .indices_2_out1_full_n(indices_23_c1_full_n),
    .indices_2_out1_write(tdf9_get_next_ijk_U0_indices_2_out1_write)
);

td_fused_top_tdf9_readInputs tdf9_readInputs_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf9_readInputs_U0_ap_start),
    .ap_done(tdf9_readInputs_U0_ap_done),
    .ap_continue(tdf9_readInputs_U0_ap_continue),
    .ap_idle(tdf9_readInputs_U0_ap_idle),
    .ap_ready(tdf9_readInputs_U0_ap_ready),
    .in_data_address0(tdf9_readInputs_U0_in_data_address0),
    .in_data_ce0(tdf9_readInputs_U0_in_data_ce0),
    .in_data_q0(in_data_q0),
    .indices_01_dout(indices_01_c_dout),
    .indices_01_empty_n(indices_01_c_empty_n),
    .indices_01_read(tdf9_readInputs_U0_indices_01_read),
    .indices_12_dout(indices_12_c_dout),
    .indices_12_empty_n(indices_12_c_empty_n),
    .indices_12_read(tdf9_readInputs_U0_indices_12_read),
    .ifmap_vec_0_0_address0(tdf9_readInputs_U0_ifmap_vec_0_0_address0),
    .ifmap_vec_0_0_ce0(tdf9_readInputs_U0_ifmap_vec_0_0_ce0),
    .ifmap_vec_0_0_we0(tdf9_readInputs_U0_ifmap_vec_0_0_we0),
    .ifmap_vec_0_0_d0(tdf9_readInputs_U0_ifmap_vec_0_0_d0),
    .ifmap_vec_0_0_address1(tdf9_readInputs_U0_ifmap_vec_0_0_address1),
    .ifmap_vec_0_0_ce1(tdf9_readInputs_U0_ifmap_vec_0_0_ce1),
    .ifmap_vec_0_0_we1(tdf9_readInputs_U0_ifmap_vec_0_0_we1),
    .ifmap_vec_0_0_d1(tdf9_readInputs_U0_ifmap_vec_0_0_d1),
    .indices_01_out_din(tdf9_readInputs_U0_indices_01_out_din),
    .indices_01_out_full_n(indices_01_c2_full_n),
    .indices_01_out_write(tdf9_readInputs_U0_indices_01_out_write),
    .indices_12_out_din(tdf9_readInputs_U0_indices_12_out_din),
    .indices_12_out_full_n(indices_12_c3_full_n),
    .indices_12_out_write(tdf9_readInputs_U0_indices_12_out_write)
);

td_fused_top_tdf9_readFilters62 tdf9_readFilters62_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf9_readFilters62_U0_ap_start),
    .ap_done(tdf9_readFilters62_U0_ap_done),
    .ap_continue(tdf9_readFilters62_U0_ap_continue),
    .ap_idle(tdf9_readFilters62_U0_ap_idle),
    .ap_ready(tdf9_readFilters62_U0_ap_ready),
    .filter_data_address0(tdf9_readFilters62_U0_filter_data_address0),
    .filter_data_ce0(tdf9_readFilters62_U0_filter_data_ce0),
    .filter_data_q0(filter_data_q0),
    .indices_23_dout(indices_23_c_dout),
    .indices_23_empty_n(indices_23_c_empty_n),
    .indices_23_read(tdf9_readFilters62_U0_indices_23_read),
    .weight_vecs_0_0_0_address0(tdf9_readFilters62_U0_weight_vecs_0_0_0_address0),
    .weight_vecs_0_0_0_ce0(tdf9_readFilters62_U0_weight_vecs_0_0_0_ce0),
    .weight_vecs_0_0_0_we0(tdf9_readFilters62_U0_weight_vecs_0_0_0_we0),
    .weight_vecs_0_0_0_d0(tdf9_readFilters62_U0_weight_vecs_0_0_0_d0)
);

td_fused_top_tdf9_dot_product tdf9_dot_product_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf9_dot_product_U0_ap_start),
    .ap_done(tdf9_dot_product_U0_ap_done),
    .ap_continue(tdf9_dot_product_U0_ap_continue),
    .ap_idle(tdf9_dot_product_U0_ap_idle),
    .ap_ready(tdf9_dot_product_U0_ap_ready),
    .ifmap_vec_0_0_address0(tdf9_dot_product_U0_ifmap_vec_0_0_address0),
    .ifmap_vec_0_0_ce0(tdf9_dot_product_U0_ifmap_vec_0_0_ce0),
    .ifmap_vec_0_0_q0(ifmap_vec_0_0_t_q0),
    .weight_vecs_0_0_0_address0(tdf9_dot_product_U0_weight_vecs_0_0_0_address0),
    .weight_vecs_0_0_0_ce0(tdf9_dot_product_U0_weight_vecs_0_0_0_ce0),
    .weight_vecs_0_0_0_q0(weight_vecs_0_0_0_t_q0),
    .products_0_address0(tdf9_dot_product_U0_products_0_address0),
    .products_0_ce0(tdf9_dot_product_U0_products_0_ce0),
    .products_0_we0(tdf9_dot_product_U0_products_0_we0),
    .products_0_d0(tdf9_dot_product_U0_products_0_d0)
);

td_fused_top_tdf9_accum_1 tdf9_accum_1_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf9_accum_1_U0_ap_start),
    .ap_done(tdf9_accum_1_U0_ap_done),
    .ap_continue(tdf9_accum_1_U0_ap_continue),
    .ap_idle(tdf9_accum_1_U0_ap_idle),
    .ap_ready(tdf9_accum_1_U0_ap_ready),
    .accum_in_0_address0(tdf9_accum_1_U0_accum_in_0_address0),
    .accum_in_0_ce0(tdf9_accum_1_U0_accum_in_0_ce0),
    .accum_in_0_q0(products_0_t_q0),
    .accum_in_0_address1(tdf9_accum_1_U0_accum_in_0_address1),
    .accum_in_0_ce1(tdf9_accum_1_U0_accum_in_0_ce1),
    .accum_in_0_q1(products_0_t_q1),
    .accum_out_address0(tdf9_accum_1_U0_accum_out_address0),
    .accum_out_ce0(tdf9_accum_1_U0_accum_out_ce0),
    .accum_out_we0(tdf9_accum_1_U0_accum_out_we0),
    .accum_out_d0(tdf9_accum_1_U0_accum_out_d0),
    .accum_out_address1(tdf9_accum_1_U0_accum_out_address1),
    .accum_out_ce1(tdf9_accum_1_U0_accum_out_ce1),
    .accum_out_we1(tdf9_accum_1_U0_accum_out_we1),
    .accum_out_d1(tdf9_accum_1_U0_accum_out_d1)
);

td_fused_top_tdf9_accum_2 tdf9_accum_2_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf9_accum_2_U0_ap_start),
    .ap_done(tdf9_accum_2_U0_ap_done),
    .ap_continue(tdf9_accum_2_U0_ap_continue),
    .ap_idle(tdf9_accum_2_U0_ap_idle),
    .ap_ready(tdf9_accum_2_U0_ap_ready),
    .accum_in_2(tdf9_accum_2_U0_accum_in_2),
    .accum_in_2_ap_vld(tdf9_accum_2_U0_accum_in_2_ap_vld),
    .accum_in_address0(tdf9_accum_2_U0_accum_in_address0),
    .accum_in_ce0(tdf9_accum_2_U0_accum_in_ce0),
    .accum_in_q0(accum1_out_0_t_q0)
);

td_fused_top_Block_entry_proc_proc429 Block_entry_proc_proc429_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(Block_entry_proc_proc429_U0_ap_start),
    .ap_done(Block_entry_proc_proc429_U0_ap_done),
    .ap_continue(Block_entry_proc_proc429_U0_ap_continue),
    .ap_idle(Block_entry_proc_proc429_U0_ap_idle),
    .ap_ready(Block_entry_proc_proc429_U0_ap_ready),
    .tmp(tmp_channel_dout),
    .ap_return(Block_entry_proc_proc429_U0_ap_return)
);

td_fused_top_tdf9_adjust tdf9_adjust_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf9_adjust_U0_ap_start),
    .ap_done(tdf9_adjust_U0_ap_done),
    .ap_continue(tdf9_adjust_U0_ap_continue),
    .ap_idle(tdf9_adjust_U0_ap_idle),
    .ap_ready(tdf9_adjust_U0_ap_ready),
    .sums_read(sums_0_dout),
    .adjustments_address0(tdf9_adjust_U0_adjustments_address0),
    .adjustments_ce0(tdf9_adjust_U0_adjustments_ce0),
    .adjustments_q0(adjustments_q0),
    .indices_23_dout(indices_23_c1_dout),
    .indices_23_empty_n(indices_23_c1_empty_n),
    .indices_23_read(tdf9_adjust_U0_indices_23_read),
    .ap_return(tdf9_adjust_U0_ap_return)
);

td_fused_top_tdf9_writeOutputs_unaligned tdf9_writeOutputs_unaligned_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf9_writeOutputs_unaligned_U0_ap_start),
    .ap_done(tdf9_writeOutputs_unaligned_U0_ap_done),
    .ap_continue(tdf9_writeOutputs_unaligned_U0_ap_continue),
    .ap_idle(tdf9_writeOutputs_unaligned_U0_ap_idle),
    .ap_ready(tdf9_writeOutputs_unaligned_U0_ap_ready),
    .indices_01_dout(indices_01_c2_dout),
    .indices_01_empty_n(indices_01_c2_empty_n),
    .indices_01_read(tdf9_writeOutputs_unaligned_U0_indices_01_read),
    .indices_12_dout(indices_12_c3_dout),
    .indices_12_empty_n(indices_12_c3_empty_n),
    .indices_12_read(tdf9_writeOutputs_unaligned_U0_indices_12_read),
    .p_read(outputs_0_dout),
    .out_data_address1(tdf9_writeOutputs_unaligned_U0_out_data_address1),
    .out_data_ce1(tdf9_writeOutputs_unaligned_U0_out_data_ce1),
    .out_data_we1(tdf9_writeOutputs_unaligned_U0_out_data_we1),
    .out_data_d1(tdf9_writeOutputs_unaligned_U0_out_data_d1)
);

td_fused_top_fifo_w16_d2_S_x6 indices_01_c_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(indices_01_c_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf9_readInputs_U0_indices_01_read),
    .if_dout(indices_01_c_dout),
    .if_full_n(indices_01_c_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf9_get_next_ijk_U0_indices_0_write),
    .if_din(tdf9_get_next_ijk_U0_indices_0_din)
);

td_fused_top_fifo_w16_d2_S_x6 indices_12_c_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(indices_12_c_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf9_readInputs_U0_indices_12_read),
    .if_dout(indices_12_c_dout),
    .if_full_n(indices_12_c_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf9_get_next_ijk_U0_indices_1_write),
    .if_din(tdf9_get_next_ijk_U0_indices_1_din)
);

td_fused_top_fifo_w6_d2_S indices_23_c_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(indices_23_c_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf9_readFilters62_U0_indices_23_read),
    .if_dout(indices_23_c_dout),
    .if_full_n(indices_23_c_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf9_get_next_ijk_U0_indices_2_out_write),
    .if_din(tdf9_get_next_ijk_U0_indices_2_out_din)
);

td_fused_top_fifo_w6_d7_S_x indices_23_c1_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(indices_23_c1_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf9_adjust_U0_indices_23_read),
    .if_dout(indices_23_c1_dout),
    .if_full_n(indices_23_c1_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf9_get_next_ijk_U0_indices_2_out1_write),
    .if_din(tdf9_get_next_ijk_U0_indices_2_out1_din)
);

td_fused_top_fifo_w4_d7_S_x indices_01_c2_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(indices_01_c2_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf9_writeOutputs_unaligned_U0_indices_01_read),
    .if_dout(indices_01_c2_dout),
    .if_full_n(indices_01_c2_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf9_readInputs_U0_indices_01_out_write),
    .if_din(tdf9_readInputs_U0_indices_01_out_din)
);

td_fused_top_fifo_w8_d7_S_x indices_12_c3_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(indices_12_c3_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf9_writeOutputs_unaligned_U0_indices_12_read),
    .if_dout(indices_12_c3_dout),
    .if_full_n(indices_12_c3_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf9_readInputs_U0_indices_12_out_write),
    .if_din(tdf9_readInputs_U0_indices_12_out_din)
);

td_fused_top_fifo_w16_d2_S_x6 tmp_channel_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(tmp_channel_empty_n),
    .if_read_ce(1'b1),
    .if_read(Block_entry_proc_proc429_U0_ap_ready),
    .if_dout(tmp_channel_dout),
    .if_full_n(tmp_channel_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf9_accum_2_U0_ap_done),
    .if_din(tdf9_accum_2_U0_accum_in_2)
);

td_fused_top_fifo_w16_d2_S_x6 sums_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(sums_0_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf9_adjust_U0_ap_ready),
    .if_dout(sums_0_dout),
    .if_full_n(sums_0_full_n),
    .if_write_ce(1'b1),
    .if_write(Block_entry_proc_proc429_U0_ap_done),
    .if_din(Block_entry_proc_proc429_U0_ap_return)
);

td_fused_top_fifo_w16_d2_S_x6 outputs_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(outputs_0_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf9_writeOutputs_unaligned_U0_ap_ready),
    .if_dout(outputs_0_dout),
    .if_full_n(outputs_0_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf9_adjust_U0_ap_done),
    .if_din(tdf9_adjust_U0_ap_return)
);

td_fused_top_start_for_tdf9_readFilters62_U0 start_for_tdf9_readFilters62_U0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(start_for_tdf9_readFilters62_U0_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf9_readFilters62_U0_ap_ready),
    .if_dout(start_for_tdf9_readFilters62_U0_dout),
    .if_full_n(start_for_tdf9_readFilters62_U0_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf9_get_next_ijk_U0_start_write),
    .if_din(start_for_tdf9_readFilters62_U0_din)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_sync_reg_tdf9_get_next_ijk_U0_ap_ready <= 1'b0;
    end else begin
        if (((ap_sync_ready & ap_start) == 1'b1)) begin
            ap_sync_reg_tdf9_get_next_ijk_U0_ap_ready <= 1'b0;
        end else begin
            ap_sync_reg_tdf9_get_next_ijk_U0_ap_ready <= ap_sync_tdf9_get_next_ijk_U0_ap_ready;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_sync_reg_tdf9_readInputs_U0_ap_ready <= 1'b0;
    end else begin
        if (((ap_sync_ready & ap_start) == 1'b1)) begin
            ap_sync_reg_tdf9_readInputs_U0_ap_ready <= 1'b0;
        end else begin
            ap_sync_reg_tdf9_readInputs_U0_ap_ready <= ap_sync_tdf9_readInputs_U0_ap_ready;
        end
    end
end

assign Block_entry_proc_proc429_U0_ap_continue = sums_0_full_n;

assign Block_entry_proc_proc429_U0_ap_start = tmp_channel_empty_n;

assign Block_entry_proc_proc429_U0_start_full_n = 1'b1;

assign Block_entry_proc_proc429_U0_start_write = 1'b0;

assign adjustments_address0 = tdf9_adjust_U0_adjustments_address0;

assign adjustments_address1 = 6'd0;

assign adjustments_ce0 = tdf9_adjust_U0_adjustments_ce0;

assign adjustments_ce1 = 1'b0;

assign adjustments_d0 = 48'd0;

assign adjustments_d1 = 48'd0;

assign adjustments_we0 = 1'b0;

assign adjustments_we1 = 1'b0;

assign ap_channel_done_accum1_out_0 = tdf9_accum_1_U0_ap_done;

assign ap_channel_done_ifmap_vec_0_0 = tdf9_readInputs_U0_ap_done;

assign ap_channel_done_outputs_0 = tdf9_adjust_U0_ap_done;

assign ap_channel_done_products_0 = tdf9_dot_product_U0_ap_done;

assign ap_channel_done_sums_0 = Block_entry_proc_proc429_U0_ap_done;

assign ap_channel_done_tmp_channel = tdf9_accum_2_U0_ap_done;

assign ap_channel_done_weight_vecs_0_0_0 = tdf9_readFilters62_U0_ap_done;

assign ap_done = tdf9_writeOutputs_unaligned_U0_ap_done;

assign ap_idle = (tdf9_writeOutputs_unaligned_U0_ap_idle & tdf9_readInputs_U0_ap_idle & tdf9_readFilters62_U0_ap_idle & tdf9_get_next_ijk_U0_ap_idle & tdf9_dot_product_U0_ap_idle & tdf9_adjust_U0_ap_idle & tdf9_accum_2_U0_ap_idle & tdf9_accum_1_U0_ap_idle & (outputs_0_empty_n ^ 1'b1) & (sums_0_empty_n ^ 1'b1) & (tmp_channel_empty_n ^ 1'b1) & (products_0_t_empty_n ^ 1'b1) & (weight_vecs_0_0_0_t_empty_n ^ 1'b1) & (ifmap_vec_0_0_t_empty_n ^ 1'b1) & (1'b1 ^ accum1_out_0_t_empty_n) & Block_entry_proc_proc429_U0_ap_idle);

assign ap_ready = ap_sync_ready;

assign ap_sync_continue = ap_continue;

assign ap_sync_done = tdf9_writeOutputs_unaligned_U0_ap_done;

assign ap_sync_ready = (ap_sync_tdf9_readInputs_U0_ap_ready & ap_sync_tdf9_get_next_ijk_U0_ap_ready);

assign ap_sync_tdf9_get_next_ijk_U0_ap_ready = (tdf9_get_next_ijk_U0_ap_ready | ap_sync_reg_tdf9_get_next_ijk_U0_ap_ready);

assign ap_sync_tdf9_readInputs_U0_ap_ready = (tdf9_readInputs_U0_ap_ready | ap_sync_reg_tdf9_readInputs_U0_ap_ready);

assign filter_data_address0 = tdf9_readFilters62_U0_filter_data_address0;

assign filter_data_address1 = 14'd0;

assign filter_data_ce0 = tdf9_readFilters62_U0_filter_data_ce0;

assign filter_data_ce1 = 1'b0;

assign filter_data_d0 = 16'd0;

assign filter_data_d1 = 16'd0;

assign filter_data_we0 = 1'b0;

assign filter_data_we1 = 1'b0;

assign in_data_address0 = tdf9_readInputs_U0_in_data_address0;

assign in_data_address1 = 14'd0;

assign in_data_ce0 = tdf9_readInputs_U0_in_data_ce0;

assign in_data_ce1 = 1'b0;

assign in_data_d0 = 64'd0;

assign in_data_d1 = 64'd0;

assign in_data_read = tdf9_readInputs_U0_in_data_write;

assign in_data_we0 = 1'b0;

assign in_data_we1 = 1'b0;

assign out_data_address0 = 12'd0;

assign out_data_address1 = tdf9_writeOutputs_unaligned_U0_out_data_address1;

assign out_data_ce0 = 1'b0;

assign out_data_ce1 = tdf9_writeOutputs_unaligned_U0_out_data_ce1;

assign out_data_d0 = 64'd0;

assign out_data_d1 = tdf9_writeOutputs_unaligned_U0_out_data_d1;

assign out_data_we0 = 1'b0;

assign out_data_we1 = tdf9_writeOutputs_unaligned_U0_out_data_we1;

assign out_data_write = tdf9_writeOutputs_unaligned_U0_out_data_write;

assign products_0_t_d1 = 16'd0;

assign products_0_t_we1 = 1'b0;

assign start_for_tdf9_readFilters62_U0_din = 1'b1;

assign tdf9_accum_1_U0_accum_out_full_n = accum1_out_0_i_full_n;

assign tdf9_accum_1_U0_ap_continue = accum1_out_0_i_full_n;

assign tdf9_accum_1_U0_ap_start = products_0_t_empty_n;

assign tdf9_accum_1_U0_start_full_n = 1'b1;

assign tdf9_accum_1_U0_start_write = 1'b0;

assign tdf9_accum_2_U0_ap_continue = tmp_channel_full_n;

assign tdf9_accum_2_U0_ap_start = accum1_out_0_t_empty_n;

assign tdf9_accum_2_U0_start_full_n = 1'b1;

assign tdf9_accum_2_U0_start_write = 1'b0;

assign tdf9_adjust_U0_ap_continue = outputs_0_full_n;

assign tdf9_adjust_U0_ap_start = sums_0_empty_n;

assign tdf9_adjust_U0_start_full_n = 1'b1;

assign tdf9_adjust_U0_start_write = 1'b0;

assign tdf9_dot_product_U0_ap_continue = products_0_i_full_n;

assign tdf9_dot_product_U0_ap_start = (weight_vecs_0_0_0_t_empty_n & ifmap_vec_0_0_t_empty_n);

assign tdf9_dot_product_U0_products_0_full_n = products_0_i_full_n;

assign tdf9_dot_product_U0_start_full_n = 1'b1;

assign tdf9_dot_product_U0_start_write = 1'b0;

assign tdf9_get_next_ijk_U0_ap_continue = 1'b1;

assign tdf9_get_next_ijk_U0_ap_start = ((ap_sync_reg_tdf9_get_next_ijk_U0_ap_ready ^ 1'b1) & ap_start);

assign tdf9_readFilters62_U0_ap_continue = weight_vecs_0_0_0_i_full_n;

assign tdf9_readFilters62_U0_ap_start = start_for_tdf9_readFilters62_U0_empty_n;

assign tdf9_readFilters62_U0_start_full_n = 1'b1;

assign tdf9_readFilters62_U0_start_write = 1'b0;

assign tdf9_readFilters62_U0_weight_vecs_0_0_0_full_n = weight_vecs_0_0_0_i_full_n;

assign tdf9_readInputs_U0_ap_continue = ifmap_vec_0_0_i_full_n;

assign tdf9_readInputs_U0_ap_start = ((ap_sync_reg_tdf9_readInputs_U0_ap_ready ^ 1'b1) & ap_start);

assign tdf9_readInputs_U0_ifmap_vec_0_0_full_n = ifmap_vec_0_0_i_full_n;

assign tdf9_readInputs_U0_in_data_full_n = in_data_empty_n;

assign tdf9_readInputs_U0_in_data_write = 1'b0;

assign tdf9_readInputs_U0_start_full_n = 1'b1;

assign tdf9_readInputs_U0_start_write = 1'b0;

assign tdf9_writeOutputs_unaligned_U0_ap_continue = ap_continue;

assign tdf9_writeOutputs_unaligned_U0_ap_start = outputs_0_empty_n;

assign tdf9_writeOutputs_unaligned_U0_out_data_full_n = out_data_full_n;

assign tdf9_writeOutputs_unaligned_U0_out_data_write = 1'b0;

assign tdf9_writeOutputs_unaligned_U0_start_full_n = 1'b1;

assign tdf9_writeOutputs_unaligned_U0_start_write = 1'b0;

endmodule //td_fused_top_dataflow_in_loop_TOP_LOOP37360
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37360_weight_vecs_0_0_0_memcore_ram (addr0, ce0, d0, we0, q0, addr1, ce1, d1, we1, q1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 9;
parameter MEM_SIZE = 512;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
output reg[DWIDTH-1:0] q1;
input clk;

reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];




always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1) 
            ram[addr1] <= d1; 
        q1 <= ram[addr1];
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37360_weight_vecs_0_0_0_memcore(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    q0,
    address1,
    ce1,
    we1,
    d1,
    q1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd512;
parameter AddressWidth = 32'd9;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;
output[DataWidth - 1:0] q1;



td_fused_top_dataflow_in_loop_TOP_LOOP37360_weight_vecs_0_0_0_memcore_ram td_fused_top_dataflow_in_loop_TOP_LOOP37360_weight_vecs_0_0_0_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 ),
    .q1( q1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_dataflow_in_loop_TOP_LOOP37360_weight_vecs_0_0_0
#(parameter
    DataWidth    = 16,
    AddressRange = 32,
    AddressWidth = 8,
    BufferCount  = 2,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire                    i_we0,
    input  wire [AddressWidth-1:0] i_address0,
    input  wire [DataWidth-1:0]    i_d0,
    output wire [DataWidth-1:0]    i_q0,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire                    t_we0,
    input  wire [AddressWidth-1:0] t_address0,
    input  wire [DataWidth-1:0]    t_d0,
    output wire [DataWidth-1:0]    t_q0
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
wire [AddressWidth+IndexWidth-1:0]   memcore_iaddr;
wire [AddressWidth+IndexWidth-1:0]   memcore_taddr;

//------------------------Instantiation------------------
assign memcore_iaddr = {i_address0, iptr};
assign memcore_taddr = {t_address0, tptr};
td_fused_top_dataflow_in_loop_TOP_LOOP37360_weight_vecs_0_0_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP37360_weight_vecs_0_0_0_memcore_U (
    .reset    ( reset ),
    .clk      ( clk ),
    .address0 ( memcore_iaddr ),
    .ce0      ( i_ce0 ),
    .we0      ( i_we0),
    .d0       ( i_d0 ),
    .q0       ( i_q0 ),
    .address1 ( memcore_taddr ),
    .ce1      ( t_ce0 ),
    .we1      ( t_we0),
    .d1       ( t_d0 ),
    .q1       ( t_q0 )

);

//------------------------Body---------------------------

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37454_accum1_out_0_memcore_ram (addr0, ce0, d0, we0, q0, addr1, ce1, d1, we1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 3;
parameter MEM_SIZE = 8;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
input clk;

reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];




always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1) 
            ram[addr1] <= d1; 
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37454_accum1_out_0_memcore(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    q0,
    address1,
    ce1,
    we1,
    d1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd8;
parameter AddressWidth = 32'd3;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;



td_fused_top_dataflow_in_loop_TOP_LOOP37454_accum1_out_0_memcore_ram td_fused_top_dataflow_in_loop_TOP_LOOP37454_accum1_out_0_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_dataflow_in_loop_TOP_LOOP37454_accum1_out_0
#(parameter
    DataWidth    = 16,
    AddressRange = 32,
    AddressWidth = 3,
    BufferCount  = 2,
    MemLatency   = 1,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire                    i_we0,
    input  wire [AddressWidth-1:0] i_address0,
    input  wire [DataWidth-1:0]    i_d0,
    output wire [DataWidth-1:0]    i_q0,
    input  wire                    i_ce1,
    input  wire                    i_we1,
    input  wire [AddressWidth-1:0] i_address1,
    input  wire [DataWidth-1:0]    i_d1,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire                    t_we0,
    input  wire [AddressWidth-1:0] t_address0,
    input  wire [DataWidth-1:0]    t_d0,
    output wire [DataWidth-1:0]    t_q0,
    input  wire                    t_ce1,
    input  wire                    t_we1,
    input  wire [AddressWidth-1:0] t_address1,
    input  wire [DataWidth-1:0]    t_d1
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth-1:0]   prev_iptr    = 1'b0; // previous initiator index
reg  [IndexWidth-1:0]   prev_tptr    = 1'b0; // previous target index
reg  [DataWidth-1:0]    reg_q0      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid0    = 1'b0; // buffer has valid data
reg  [DataWidth-1:0]    reg_q1      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid1    = 1'b0; // buffer has valid data
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
// buffer signals
wire [BufferCount-1:0] buf_ce0;
wire [BufferCount-1:0] buf_we0;
wire [AddressWidth-1:0] buf_a0_0, buf_a0_1;
wire [DataWidth-1:0] buf_d0_0, buf_d0_1;
wire [DataWidth-1:0] buf_q0_0, buf_q0_1;
wire [BufferCount-1:0] buf_ce1;
wire [BufferCount-1:0] buf_we1;
wire [AddressWidth-1:0] buf_a1_0, buf_a1_1;
wire [DataWidth-1:0] buf_d1_0, buf_d1_1;
//------------------------Instantiation------------------
//genvar i;
        td_fused_top_dataflow_in_loop_TOP_LOOP37454_accum1_out_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP37454_accum1_out_0_memcore_U_0 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_0 ),
            .ce0      ( buf_ce0[ 0 ] ),
            .we0      ( buf_we0[ 0 ] ),
            .d0       ( buf_d0_0 ),
            .q0       ( buf_q0_0 ),
            .address1 ( buf_a1_0 ),
            .ce1      ( buf_ce1[ 0 ] ),
            .we1      ( buf_we1[ 0 ] ),
            .d1       ( buf_d1_0 )
        );
        td_fused_top_dataflow_in_loop_TOP_LOOP37454_accum1_out_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP37454_accum1_out_0_memcore_U_1 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_1 ),
            .ce0      ( buf_ce0[ 1 ] ),
            .we0      ( buf_we0[ 1 ] ),
            .d0       ( buf_d0_1 ),
            .q0       ( buf_q0_1 ),
            .address1 ( buf_a1_1 ),
            .ce1      ( buf_ce1[ 1 ] ),
            .we1      ( buf_we1[ 1 ] ),
            .d1       ( buf_d1_1 )
        );

//++++++++++++++++++++++++buffer signals+++++++++++++++++
        assign buf_ce0[ 0 ] = (tptr ==  0  && empty_n) ? t_ce0
                             : (iptr ==  0 ) ? i_ce0 : 1'b0;
        assign buf_a0_0  = (tptr ==  0  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 0 ] = (tptr ==  0  && empty_n)  ? t_we0
                             : (iptr ==  0 ) ? i_we0 : 1'b0;
        assign buf_d0_0  = (tptr ==  0  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 0 ] = (tptr ==  0  && empty_n) ? t_ce1
                             : (iptr ==  0 ) ? i_ce1 : 1'b0;
        assign buf_a1_0  = (tptr ==  0  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 0 ] = (tptr ==  0  && empty_n)  ? t_we1
                             : (iptr ==  0 ) ? i_we1 : 1'b0;
        assign buf_d1_0  = (tptr ==  0  && empty_n) ? t_d1       : i_d1;
        assign buf_ce0[ 1 ] = (tptr ==  1  && empty_n) ? t_ce0
                             : (iptr ==  1 ) ? i_ce0 : 1'b0;
        assign buf_a0_1  = (tptr ==  1  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 1 ] = (tptr ==  1  && empty_n)  ? t_we0
                             : (iptr ==  1 ) ? i_we0 : 1'b0;
        assign buf_d0_1  = (tptr ==  1  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 1 ] = (tptr ==  1  && empty_n) ? t_ce1
                             : (iptr ==  1 ) ? i_ce1 : 1'b0;
        assign buf_a1_1  = (tptr ==  1  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 1 ] = (tptr ==  1  && empty_n)  ? t_we1
                             : (iptr ==  1 ) ? i_we1 : 1'b0;
        assign buf_d1_1  = (tptr ==  1  && empty_n) ? t_d1       : i_d1;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//------------------------Body---------------------------
assign i_q0      = (prev_iptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign t_q0      = reg_valid0 ? reg_q0 : (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// prev_iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_iptr <= 1'b0;
    else begin
        prev_iptr <= iptr;
    end
end

// prev_tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_tptr <= 1'b0;
    else begin
        prev_tptr <= tptr;
    end
end

// reg_q0 and reg_valid0
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q0     <= 1'b0;
        reg_valid0 <= 1'b0;
    end else if (!t_ce0 && !reg_valid0) begin
        reg_q0     <= (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
        reg_valid0 <= 1'b1;
    end else if (t_ce0) begin
        reg_valid0 <= 1'b0;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37454_ifmap_vec_memcore_ram (addr0, ce0, d0, we0, q0, addr1, ce1, d1, we1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 9;
parameter MEM_SIZE = 288;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
input clk;

reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];




always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1) 
            ram[addr1] <= d1; 
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37454_ifmap_vec_memcore(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    q0,
    address1,
    ce1,
    we1,
    d1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd288;
parameter AddressWidth = 32'd9;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;



td_fused_top_dataflow_in_loop_TOP_LOOP37454_ifmap_vec_memcore_ram td_fused_top_dataflow_in_loop_TOP_LOOP37454_ifmap_vec_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_dataflow_in_loop_TOP_LOOP37454_ifmap_vec
#(parameter
    DataWidth    = 16,
    AddressRange = 32,
    AddressWidth = 9,
    BufferCount  = 2,
    MemLatency   = 1,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire                    i_we0,
    input  wire [AddressWidth-1:0] i_address0,
    input  wire [DataWidth-1:0]    i_d0,
    output wire [DataWidth-1:0]    i_q0,
    input  wire                    i_ce1,
    input  wire                    i_we1,
    input  wire [AddressWidth-1:0] i_address1,
    input  wire [DataWidth-1:0]    i_d1,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire                    t_we0,
    input  wire [AddressWidth-1:0] t_address0,
    input  wire [DataWidth-1:0]    t_d0,
    output wire [DataWidth-1:0]    t_q0,
    input  wire                    t_ce1,
    input  wire                    t_we1,
    input  wire [AddressWidth-1:0] t_address1,
    input  wire [DataWidth-1:0]    t_d1
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth-1:0]   prev_iptr    = 1'b0; // previous initiator index
reg  [IndexWidth-1:0]   prev_tptr    = 1'b0; // previous target index
reg  [DataWidth-1:0]    reg_q0      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid0    = 1'b0; // buffer has valid data
reg  [DataWidth-1:0]    reg_q1      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid1    = 1'b0; // buffer has valid data
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
// buffer signals
wire [BufferCount-1:0] buf_ce0;
wire [BufferCount-1:0] buf_we0;
wire [AddressWidth-1:0] buf_a0_0, buf_a0_1;
wire [DataWidth-1:0] buf_d0_0, buf_d0_1;
wire [DataWidth-1:0] buf_q0_0, buf_q0_1;
wire [BufferCount-1:0] buf_ce1;
wire [BufferCount-1:0] buf_we1;
wire [AddressWidth-1:0] buf_a1_0, buf_a1_1;
wire [DataWidth-1:0] buf_d1_0, buf_d1_1;
//------------------------Instantiation------------------
//genvar i;
        td_fused_top_dataflow_in_loop_TOP_LOOP37454_ifmap_vec_memcore td_fused_top_dataflow_in_loop_TOP_LOOP37454_ifmap_vec_memcore_U_0 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_0 ),
            .ce0      ( buf_ce0[ 0 ] ),
            .we0      ( buf_we0[ 0 ] ),
            .d0       ( buf_d0_0 ),
            .q0       ( buf_q0_0 ),
            .address1 ( buf_a1_0 ),
            .ce1      ( buf_ce1[ 0 ] ),
            .we1      ( buf_we1[ 0 ] ),
            .d1       ( buf_d1_0 )
        );
        td_fused_top_dataflow_in_loop_TOP_LOOP37454_ifmap_vec_memcore td_fused_top_dataflow_in_loop_TOP_LOOP37454_ifmap_vec_memcore_U_1 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_1 ),
            .ce0      ( buf_ce0[ 1 ] ),
            .we0      ( buf_we0[ 1 ] ),
            .d0       ( buf_d0_1 ),
            .q0       ( buf_q0_1 ),
            .address1 ( buf_a1_1 ),
            .ce1      ( buf_ce1[ 1 ] ),
            .we1      ( buf_we1[ 1 ] ),
            .d1       ( buf_d1_1 )
        );

//++++++++++++++++++++++++buffer signals+++++++++++++++++
        assign buf_ce0[ 0 ] = (tptr ==  0  && empty_n) ? t_ce0
                             : (iptr ==  0 ) ? i_ce0 : 1'b0;
        assign buf_a0_0  = (tptr ==  0  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 0 ] = (tptr ==  0  && empty_n)  ? t_we0
                             : (iptr ==  0 ) ? i_we0 : 1'b0;
        assign buf_d0_0  = (tptr ==  0  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 0 ] = (tptr ==  0  && empty_n) ? t_ce1
                             : (iptr ==  0 ) ? i_ce1 : 1'b0;
        assign buf_a1_0  = (tptr ==  0  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 0 ] = (tptr ==  0  && empty_n)  ? t_we1
                             : (iptr ==  0 ) ? i_we1 : 1'b0;
        assign buf_d1_0  = (tptr ==  0  && empty_n) ? t_d1       : i_d1;
        assign buf_ce0[ 1 ] = (tptr ==  1  && empty_n) ? t_ce0
                             : (iptr ==  1 ) ? i_ce0 : 1'b0;
        assign buf_a0_1  = (tptr ==  1  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 1 ] = (tptr ==  1  && empty_n)  ? t_we0
                             : (iptr ==  1 ) ? i_we0 : 1'b0;
        assign buf_d0_1  = (tptr ==  1  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 1 ] = (tptr ==  1  && empty_n) ? t_ce1
                             : (iptr ==  1 ) ? i_ce1 : 1'b0;
        assign buf_a1_1  = (tptr ==  1  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 1 ] = (tptr ==  1  && empty_n)  ? t_we1
                             : (iptr ==  1 ) ? i_we1 : 1'b0;
        assign buf_d1_1  = (tptr ==  1  && empty_n) ? t_d1       : i_d1;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//------------------------Body---------------------------
assign i_q0      = (prev_iptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign t_q0      = reg_valid0 ? reg_q0 : (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// prev_iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_iptr <= 1'b0;
    else begin
        prev_iptr <= iptr;
    end
end

// prev_tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_tptr <= 1'b0;
    else begin
        prev_tptr <= tptr;
    end
end

// reg_q0 and reg_valid0
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q0     <= 1'b0;
        reg_valid0 <= 1'b0;
    end else if (!t_ce0 && !reg_valid0) begin
        reg_q0     <= (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
        reg_valid0 <= 1'b1;
    end else if (t_ce0) begin
        reg_valid0 <= 1'b0;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37454_products_0_memcore_ram (addr0, ce0, d0, we0, q0, addr1, ce1, q1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 9;
parameter MEM_SIZE = 288;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
output reg[DWIDTH-1:0] q1;
input clk;

reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];




always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        q1 <= ram[addr1];
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37454_products_0_memcore(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    q0,
    address1,
    ce1,
    q1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd288;
parameter AddressWidth = 32'd9;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
output[DataWidth - 1:0] q1;



td_fused_top_dataflow_in_loop_TOP_LOOP37454_products_0_memcore_ram td_fused_top_dataflow_in_loop_TOP_LOOP37454_products_0_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .q1( q1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_dataflow_in_loop_TOP_LOOP37454_products_0
#(parameter
    DataWidth    = 16,
    AddressRange = 32,
    AddressWidth = 9,
    BufferCount  = 2,
    MemLatency   = 1,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire                    i_we0,
    input  wire [AddressWidth-1:0] i_address0,
    input  wire [DataWidth-1:0]    i_d0,
    output wire [DataWidth-1:0]    i_q0,
    input  wire                    i_ce1,
    input  wire [AddressWidth-1:0] i_address1,
    output wire [DataWidth-1:0]    i_q1,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire                    t_we0,
    input  wire [AddressWidth-1:0] t_address0,
    input  wire [DataWidth-1:0]    t_d0,
    output wire [DataWidth-1:0]    t_q0,
    input  wire                    t_ce1,
    input  wire [AddressWidth-1:0] t_address1,
    output wire [DataWidth-1:0]    t_q1
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth-1:0]   prev_iptr    = 1'b0; // previous initiator index
reg  [IndexWidth-1:0]   prev_tptr    = 1'b0; // previous target index
reg  [DataWidth-1:0]    reg_q0      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid0    = 1'b0; // buffer has valid data
reg  [DataWidth-1:0]    reg_q1      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid1    = 1'b0; // buffer has valid data
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
// buffer signals
wire [BufferCount-1:0] buf_ce0;
wire [BufferCount-1:0] buf_we0;
wire [AddressWidth-1:0] buf_a0_0, buf_a0_1;
wire [DataWidth-1:0] buf_d0_0, buf_d0_1;
wire [DataWidth-1:0] buf_q0_0, buf_q0_1;
wire [BufferCount-1:0] buf_ce1;
wire [AddressWidth-1:0] buf_a1_0, buf_a1_1;
wire [DataWidth-1:0] buf_q1_0, buf_q1_1;
//------------------------Instantiation------------------
//genvar i;
        td_fused_top_dataflow_in_loop_TOP_LOOP37454_products_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP37454_products_0_memcore_U_0 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_0 ),
            .ce0      ( buf_ce0[ 0 ] ),
            .we0      ( buf_we0[ 0 ] ),
            .d0       ( buf_d0_0 ),
            .q0       ( buf_q0_0 ),
            .address1 ( buf_a1_0 ),
            .ce1      ( buf_ce1[ 0 ] ),
            .q1       ( buf_q1_0 )
        );
        td_fused_top_dataflow_in_loop_TOP_LOOP37454_products_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP37454_products_0_memcore_U_1 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_1 ),
            .ce0      ( buf_ce0[ 1 ] ),
            .we0      ( buf_we0[ 1 ] ),
            .d0       ( buf_d0_1 ),
            .q0       ( buf_q0_1 ),
            .address1 ( buf_a1_1 ),
            .ce1      ( buf_ce1[ 1 ] ),
            .q1       ( buf_q1_1 )
        );

//++++++++++++++++++++++++buffer signals+++++++++++++++++
        assign buf_ce0[ 0 ] = (tptr ==  0  && empty_n) ? t_ce0
                             : (iptr ==  0 ) ? i_ce0 : 1'b0;
        assign buf_a0_0  = (tptr ==  0  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 0 ] = (tptr ==  0  && empty_n)  ? t_we0
                             : (iptr ==  0 ) ? i_we0 : 1'b0;
        assign buf_d0_0  = (tptr ==  0  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 0 ] = (tptr ==  0  && empty_n) ? t_ce1
                             : (iptr ==  0 ) ? i_ce1 : 1'b0;
        assign buf_a1_0  = (tptr ==  0  && empty_n) ?  t_address1 : i_address1;
        assign buf_ce0[ 1 ] = (tptr ==  1  && empty_n) ? t_ce0
                             : (iptr ==  1 ) ? i_ce0 : 1'b0;
        assign buf_a0_1  = (tptr ==  1  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 1 ] = (tptr ==  1  && empty_n)  ? t_we0
                             : (iptr ==  1 ) ? i_we0 : 1'b0;
        assign buf_d0_1  = (tptr ==  1  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 1 ] = (tptr ==  1  && empty_n) ? t_ce1
                             : (iptr ==  1 ) ? i_ce1 : 1'b0;
        assign buf_a1_1  = (tptr ==  1  && empty_n) ?  t_address1 : i_address1;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//------------------------Body---------------------------
assign i_q0      = (prev_iptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign t_q0      = reg_valid0 ? reg_q0 : (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign i_q1      = (prev_iptr == 1'b1 ? buf_q1_1 : buf_q1_0);
assign t_q1      = reg_valid1 ? reg_q1 : (prev_tptr == 1'b1 ? buf_q1_1 : buf_q1_0);

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// prev_iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_iptr <= 1'b0;
    else begin
        prev_iptr <= iptr;
    end
end

// prev_tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_tptr <= 1'b0;
    else begin
        prev_tptr <= tptr;
    end
end

// reg_q0 and reg_valid0
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q0     <= 1'b0;
        reg_valid0 <= 1'b0;
    end else if (!t_ce0 && !reg_valid0) begin
        reg_q0     <= (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
        reg_valid0 <= 1'b1;
    end else if (t_ce0) begin
        reg_valid0 <= 1'b0;
    end
end

// reg_q1 and reg_valid1
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q1     <= 1'b0;
        reg_valid1 <= 1'b0;
    end else if (!t_ce1 && !reg_valid1) begin
        reg_q1     <= (prev_tptr == 1'b1 ? buf_q1_1 : buf_q1_0);
        reg_valid1 <= 1'b1;
    end else if (t_ce1) begin
        reg_valid1 <= 1'b0;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_dataflow_in_loop_TOP_LOOP37454 (
        ap_clk,
        ap_rst,
        in_data_address0,
        in_data_ce0,
        in_data_d0,
        in_data_q0,
        in_data_we0,
        in_data_address1,
        in_data_ce1,
        in_data_d1,
        in_data_q1,
        in_data_we1,
        filter_data_address0,
        filter_data_ce0,
        filter_data_d0,
        filter_data_q0,
        filter_data_we0,
        filter_data_address1,
        filter_data_ce1,
        filter_data_d1,
        filter_data_q1,
        filter_data_we1,
        adjustments_address0,
        adjustments_ce0,
        adjustments_d0,
        adjustments_q0,
        adjustments_we0,
        adjustments_address1,
        adjustments_ce1,
        adjustments_d1,
        adjustments_q1,
        adjustments_we1,
        out_data_address0,
        out_data_ce0,
        out_data_d0,
        out_data_q0,
        out_data_we0,
        out_data_address1,
        out_data_ce1,
        out_data_d1,
        out_data_q1,
        out_data_we1,
        ap_start,
        in_data_empty_n,
        in_data_read,
        out_data_full_n,
        out_data_write,
        ap_done,
        ap_ready,
        ap_idle,
        ap_continue
);


input   ap_clk;
input   ap_rst;
output  [12:0] in_data_address0;
output   in_data_ce0;
output  [63:0] in_data_d0;
input  [63:0] in_data_q0;
output   in_data_we0;
output  [12:0] in_data_address1;
output   in_data_ce1;
output  [63:0] in_data_d1;
input  [63:0] in_data_q1;
output   in_data_we1;
output  [16:0] filter_data_address0;
output   filter_data_ce0;
output  [15:0] filter_data_d0;
input  [15:0] filter_data_q0;
output   filter_data_we0;
output  [16:0] filter_data_address1;
output   filter_data_ce1;
output  [15:0] filter_data_d1;
input  [15:0] filter_data_q1;
output   filter_data_we1;
output  [7:0] adjustments_address0;
output   adjustments_ce0;
output  [47:0] adjustments_d0;
input  [47:0] adjustments_q0;
output   adjustments_we0;
output  [7:0] adjustments_address1;
output   adjustments_ce1;
output  [47:0] adjustments_d1;
input  [47:0] adjustments_q1;
output   adjustments_we1;
output  [13:0] out_data_address0;
output   out_data_ce0;
output  [63:0] out_data_d0;
input  [63:0] out_data_q0;
output   out_data_we0;
output  [13:0] out_data_address1;
output   out_data_ce1;
output  [63:0] out_data_d1;
input  [63:0] out_data_q1;
output   out_data_we1;
input   ap_start;
input   in_data_empty_n;
output   in_data_read;
input   out_data_full_n;
output   out_data_write;
output   ap_done;
output   ap_ready;
output   ap_idle;
input   ap_continue;

wire   [15:0] ifmap_vec_i_q0;
wire   [15:0] ifmap_vec_t_q0;
wire   [15:0] weight_vecs_0_i_q0;
wire   [15:0] weight_vecs_0_t_q0;
wire   [15:0] products_0_i_q0;
wire   [15:0] products_0_i_q1;
wire   [15:0] products_0_t_q0;
wire   [15:0] products_0_t_q1;
wire   [15:0] accum1_out_0_i_q0;
wire   [15:0] accum1_out_0_t_q0;
wire    tdf8_get_next_ijk_U0_ap_start;
wire    tdf8_get_next_ijk_U0_ap_done;
wire    tdf8_get_next_ijk_U0_ap_continue;
wire    tdf8_get_next_ijk_U0_ap_idle;
wire    tdf8_get_next_ijk_U0_ap_ready;
wire    tdf8_get_next_ijk_U0_start_out;
wire    tdf8_get_next_ijk_U0_start_write;
wire   [7:0] tdf8_get_next_ijk_U0_input_indices_2_out_din;
wire    tdf8_get_next_ijk_U0_input_indices_2_out_write;
wire   [7:0] tdf8_get_next_ijk_U0_input_indices_2_out1_din;
wire    tdf8_get_next_ijk_U0_input_indices_2_out1_write;
wire   [3:0] tdf8_get_next_ijk_U0_output_indices_0_din;
wire    tdf8_get_next_ijk_U0_output_indices_0_write;
wire   [7:0] tdf8_get_next_ijk_U0_output_indices_1_din;
wire    tdf8_get_next_ijk_U0_output_indices_1_write;
wire    tdf8_get_next_ijk_U0_resetMaximum_din;
wire    tdf8_get_next_ijk_U0_resetMaximum_write;
wire    tdf8_get_next_ijk_U0_storeOutput_din;
wire    tdf8_get_next_ijk_U0_storeOutput_write;
wire   [15:0] tdf8_get_next_ijk_U0_ap_return_0;
wire   [15:0] tdf8_get_next_ijk_U0_ap_return_1;
wire    ap_channel_done_input_indices_1;
wire    input_indices_1_full_n;
reg    ap_sync_reg_channel_write_input_indices_1;
wire    ap_sync_channel_write_input_indices_1;
wire    ap_channel_done_input_indices_0;
wire    input_indices_0_full_n;
reg    ap_sync_reg_channel_write_input_indices_0;
wire    ap_sync_channel_write_input_indices_0;
wire    tdf8_readInputs57_U0_ap_start;
wire    tdf8_readInputs57_U0_ap_done;
wire    tdf8_readInputs57_U0_ap_continue;
wire    tdf8_readInputs57_U0_ap_idle;
wire    tdf8_readInputs57_U0_ap_ready;
wire   [12:0] tdf8_readInputs57_U0_in_data_address0;
wire    tdf8_readInputs57_U0_in_data_ce0;
wire   [8:0] tdf8_readInputs57_U0_ifmap_vec_address0;
wire    tdf8_readInputs57_U0_ifmap_vec_ce0;
wire    tdf8_readInputs57_U0_ifmap_vec_we0;
wire   [15:0] tdf8_readInputs57_U0_ifmap_vec_d0;
wire   [8:0] tdf8_readInputs57_U0_ifmap_vec_address1;
wire    tdf8_readInputs57_U0_ifmap_vec_ce1;
wire    tdf8_readInputs57_U0_ifmap_vec_we1;
wire   [15:0] tdf8_readInputs57_U0_ifmap_vec_d1;
wire    tdf8_readInputs57_U0_in_data_full_n;
wire    tdf8_readInputs57_U0_in_data_write;
wire    ap_channel_done_ifmap_vec;
wire    tdf8_readInputs57_U0_ifmap_vec_full_n;
wire    tdf8_readFilters56_U0_ap_start;
wire    tdf8_readFilters56_U0_ap_done;
wire    tdf8_readFilters56_U0_ap_continue;
wire    tdf8_readFilters56_U0_ap_idle;
wire    tdf8_readFilters56_U0_ap_ready;
wire   [16:0] tdf8_readFilters56_U0_filter_data_address0;
wire    tdf8_readFilters56_U0_filter_data_ce0;
wire    tdf8_readFilters56_U0_input_indices_23_read;
wire   [8:0] tdf8_readFilters56_U0_weight_vecs_0_address0;
wire    tdf8_readFilters56_U0_weight_vecs_0_ce0;
wire    tdf8_readFilters56_U0_weight_vecs_0_we0;
wire   [15:0] tdf8_readFilters56_U0_weight_vecs_0_d0;
wire    ap_channel_done_weight_vecs_0;
wire    tdf8_readFilters56_U0_weight_vecs_0_full_n;
wire    tdf8_dot_product_U0_ap_start;
wire    tdf8_dot_product_U0_ap_done;
wire    tdf8_dot_product_U0_ap_continue;
wire    tdf8_dot_product_U0_ap_idle;
wire    tdf8_dot_product_U0_ap_ready;
wire   [8:0] tdf8_dot_product_U0_ifmap_vec_address0;
wire    tdf8_dot_product_U0_ifmap_vec_ce0;
wire   [8:0] tdf8_dot_product_U0_weight_vecs_0_address0;
wire    tdf8_dot_product_U0_weight_vecs_0_ce0;
wire   [8:0] tdf8_dot_product_U0_products_0_address0;
wire    tdf8_dot_product_U0_products_0_ce0;
wire    tdf8_dot_product_U0_products_0_we0;
wire   [15:0] tdf8_dot_product_U0_products_0_d0;
wire    ap_channel_done_products_0;
wire    tdf8_dot_product_U0_products_0_full_n;
wire    tdf8_accum_1_U0_ap_start;
wire    tdf8_accum_1_U0_ap_done;
wire    tdf8_accum_1_U0_ap_continue;
wire    tdf8_accum_1_U0_ap_idle;
wire    tdf8_accum_1_U0_ap_ready;
wire   [8:0] tdf8_accum_1_U0_accum_in_0_address0;
wire    tdf8_accum_1_U0_accum_in_0_ce0;
wire   [8:0] tdf8_accum_1_U0_accum_in_0_address1;
wire    tdf8_accum_1_U0_accum_in_0_ce1;
wire   [2:0] tdf8_accum_1_U0_accum_out_address0;
wire    tdf8_accum_1_U0_accum_out_ce0;
wire    tdf8_accum_1_U0_accum_out_we0;
wire   [15:0] tdf8_accum_1_U0_accum_out_d0;
wire   [2:0] tdf8_accum_1_U0_accum_out_address1;
wire    tdf8_accum_1_U0_accum_out_ce1;
wire    tdf8_accum_1_U0_accum_out_we1;
wire   [15:0] tdf8_accum_1_U0_accum_out_d1;
wire    ap_channel_done_accum1_out_0;
wire    tdf8_accum_1_U0_accum_out_full_n;
wire    tdf8_accum_2_U0_ap_start;
wire    tdf8_accum_2_U0_ap_done;
wire    tdf8_accum_2_U0_ap_continue;
wire    tdf8_accum_2_U0_ap_idle;
wire    tdf8_accum_2_U0_ap_ready;
wire   [15:0] tdf8_accum_2_U0_accum_in_4;
wire    tdf8_accum_2_U0_accum_in_4_ap_vld;
wire   [2:0] tdf8_accum_2_U0_accum_in_address0;
wire    tdf8_accum_2_U0_accum_in_ce0;
wire    ap_channel_done_tmp_channel;
wire    tmp_channel_full_n;
wire    Block_entry_proc_proc424_U0_ap_start;
wire    Block_entry_proc_proc424_U0_ap_done;
wire    Block_entry_proc_proc424_U0_ap_continue;
wire    Block_entry_proc_proc424_U0_ap_idle;
wire    Block_entry_proc_proc424_U0_ap_ready;
wire   [15:0] Block_entry_proc_proc424_U0_ap_return;
wire    ap_channel_done_sums_0;
wire    sums_0_full_n;
wire    tdf8_adjust_U0_ap_start;
wire    tdf8_adjust_U0_ap_done;
wire    tdf8_adjust_U0_ap_continue;
wire    tdf8_adjust_U0_ap_idle;
wire    tdf8_adjust_U0_ap_ready;
wire   [7:0] tdf8_adjust_U0_adjustments_address0;
wire    tdf8_adjust_U0_adjustments_ce0;
wire    tdf8_adjust_U0_input_indices_23_read;
wire   [15:0] tdf8_adjust_U0_ap_return;
wire    ap_channel_done_outputs_0;
wire    outputs_0_full_n;
wire    tdf8_poolOutputs_U0_ap_start;
wire    tdf8_poolOutputs_U0_ap_done;
wire    tdf8_poolOutputs_U0_ap_continue;
wire    tdf8_poolOutputs_U0_ap_idle;
wire    tdf8_poolOutputs_U0_ap_ready;
wire    tdf8_poolOutputs_U0_output_indices_04_read;
wire    tdf8_poolOutputs_U0_output_indices_15_read;
wire    tdf8_poolOutputs_U0_resetMaximum6_read;
wire    tdf8_poolOutputs_U0_storeOutput7_read;
wire   [13:0] tdf8_poolOutputs_U0_out_data_address1;
wire    tdf8_poolOutputs_U0_out_data_ce1;
wire    tdf8_poolOutputs_U0_out_data_we1;
wire   [63:0] tdf8_poolOutputs_U0_out_data_d1;
wire    tdf8_poolOutputs_U0_out_data_full_n;
wire    tdf8_poolOutputs_U0_out_data_write;
wire    ap_sync_continue;
wire    ifmap_vec_i_full_n;
wire    ifmap_vec_t_empty_n;
wire    weight_vecs_0_i_full_n;
wire    weight_vecs_0_t_empty_n;
wire    products_0_i_full_n;
wire    products_0_t_empty_n;
wire   [15:0] products_0_t_d1;
wire    products_0_t_we1;
wire    accum1_out_0_i_full_n;
wire    accum1_out_0_t_empty_n;
wire    input_indices_23_c_full_n;
wire   [7:0] input_indices_23_c_dout;
wire    input_indices_23_c_empty_n;
wire    input_indices_23_c1_full_n;
wire   [7:0] input_indices_23_c1_dout;
wire    input_indices_23_c1_empty_n;
wire    output_indices_04_c_full_n;
wire   [3:0] output_indices_04_c_dout;
wire    output_indices_04_c_empty_n;
wire    output_indices_15_c_full_n;
wire   [7:0] output_indices_15_c_dout;
wire    output_indices_15_c_empty_n;
wire   [0:0] resetMaximum6_c_din;
wire    resetMaximum6_c_full_n;
wire   [0:0] resetMaximum6_c_dout;
wire    resetMaximum6_c_empty_n;
wire   [0:0] storeOutput7_c_din;
wire    storeOutput7_c_full_n;
wire   [0:0] storeOutput7_c_dout;
wire    storeOutput7_c_empty_n;
wire   [15:0] input_indices_0_dout;
wire    input_indices_0_empty_n;
wire   [15:0] input_indices_1_dout;
wire    input_indices_1_empty_n;
wire   [15:0] tmp_channel_dout;
wire    tmp_channel_empty_n;
wire   [15:0] sums_0_dout;
wire    sums_0_empty_n;
wire   [15:0] outputs_0_dout;
wire    outputs_0_empty_n;
wire    ap_sync_done;
wire    ap_sync_ready;
reg    ap_sync_reg_tdf8_get_next_ijk_U0_ap_ready;
wire    ap_sync_tdf8_get_next_ijk_U0_ap_ready;
reg    ap_sync_reg_tdf8_readInputs57_U0_ap_ready;
wire    ap_sync_tdf8_readInputs57_U0_ap_ready;
wire   [0:0] start_for_tdf8_readFilters56_U0_din;
wire    start_for_tdf8_readFilters56_U0_full_n;
wire   [0:0] start_for_tdf8_readFilters56_U0_dout;
wire    start_for_tdf8_readFilters56_U0_empty_n;
wire    tdf8_readInputs57_U0_start_full_n;
wire    tdf8_readInputs57_U0_start_write;
wire    tdf8_readFilters56_U0_start_full_n;
wire    tdf8_readFilters56_U0_start_write;
wire    tdf8_dot_product_U0_start_full_n;
wire    tdf8_dot_product_U0_start_write;
wire    tdf8_accum_1_U0_start_full_n;
wire    tdf8_accum_1_U0_start_write;
wire    tdf8_accum_2_U0_start_full_n;
wire    tdf8_accum_2_U0_start_write;
wire    Block_entry_proc_proc424_U0_start_full_n;
wire    Block_entry_proc_proc424_U0_start_write;
wire    tdf8_adjust_U0_start_full_n;
wire    tdf8_adjust_U0_start_write;
wire    tdf8_poolOutputs_U0_start_full_n;
wire    tdf8_poolOutputs_U0_start_write;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_sync_reg_channel_write_input_indices_1 = 1'b0;
#0 ap_sync_reg_channel_write_input_indices_0 = 1'b0;
#0 ap_sync_reg_tdf8_get_next_ijk_U0_ap_ready = 1'b0;
#0 ap_sync_reg_tdf8_readInputs57_U0_ap_ready = 1'b0;
end

td_fused_top_dataflow_in_loop_TOP_LOOP37454_ifmap_vec #(
    .DataWidth( 16 ),
    .AddressRange( 288 ),
    .AddressWidth( 9 ))
ifmap_vec_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf8_readInputs57_U0_ap_done),
    .i_full_n(ifmap_vec_i_full_n),
    .i_ce0(tdf8_readInputs57_U0_ifmap_vec_ce0),
    .i_we0(tdf8_readInputs57_U0_ifmap_vec_we0),
    .i_address0(tdf8_readInputs57_U0_ifmap_vec_address0),
    .i_d0(tdf8_readInputs57_U0_ifmap_vec_d0),
    .i_q0(ifmap_vec_i_q0),
    .i_ce1(tdf8_readInputs57_U0_ifmap_vec_ce1),
    .i_we1(tdf8_readInputs57_U0_ifmap_vec_we1),
    .i_address1(tdf8_readInputs57_U0_ifmap_vec_address1),
    .i_d1(tdf8_readInputs57_U0_ifmap_vec_d1),
    .t_ce(1'b1),
    .t_read(tdf8_dot_product_U0_ap_ready),
    .t_empty_n(ifmap_vec_t_empty_n),
    .t_ce0(tdf8_dot_product_U0_ifmap_vec_ce0),
    .t_we0(1'b0),
    .t_address0(tdf8_dot_product_U0_ifmap_vec_address0),
    .t_d0(16'd0),
    .t_q0(ifmap_vec_t_q0),
    .t_ce1(1'b0),
    .t_we1(1'b0),
    .t_address1(9'd0),
    .t_d1(16'd0)
);

td_fused_top_dataflow_in_loop_TOP_LOOP37454_weight_vecs_0 #(
    .DataWidth( 16 ),
    .AddressRange( 288 ),
    .AddressWidth( 9 ))
weight_vecs_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf8_readFilters56_U0_ap_done),
    .i_full_n(weight_vecs_0_i_full_n),
    .i_ce0(tdf8_readFilters56_U0_weight_vecs_0_ce0),
    .i_we0(tdf8_readFilters56_U0_weight_vecs_0_we0),
    .i_address0(tdf8_readFilters56_U0_weight_vecs_0_address0),
    .i_d0(tdf8_readFilters56_U0_weight_vecs_0_d0),
    .i_q0(weight_vecs_0_i_q0),
    .t_ce(1'b1),
    .t_read(tdf8_dot_product_U0_ap_ready),
    .t_empty_n(weight_vecs_0_t_empty_n),
    .t_ce0(tdf8_dot_product_U0_weight_vecs_0_ce0),
    .t_we0(1'b0),
    .t_address0(tdf8_dot_product_U0_weight_vecs_0_address0),
    .t_d0(16'd0),
    .t_q0(weight_vecs_0_t_q0)
);

td_fused_top_dataflow_in_loop_TOP_LOOP37454_products_0 #(
    .DataWidth( 16 ),
    .AddressRange( 288 ),
    .AddressWidth( 9 ))
products_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf8_dot_product_U0_ap_done),
    .i_full_n(products_0_i_full_n),
    .i_ce0(tdf8_dot_product_U0_products_0_ce0),
    .i_we0(tdf8_dot_product_U0_products_0_we0),
    .i_address0(tdf8_dot_product_U0_products_0_address0),
    .i_d0(tdf8_dot_product_U0_products_0_d0),
    .i_q0(products_0_i_q0),
    .i_ce1(1'b0),
    .i_address1(9'd0),
    .i_q1(products_0_i_q1),
    .t_ce(1'b1),
    .t_read(tdf8_accum_1_U0_ap_ready),
    .t_empty_n(products_0_t_empty_n),
    .t_ce0(tdf8_accum_1_U0_accum_in_0_ce0),
    .t_we0(1'b0),
    .t_address0(tdf8_accum_1_U0_accum_in_0_address0),
    .t_d0(16'd0),
    .t_q0(products_0_t_q0),
    .t_ce1(tdf8_accum_1_U0_accum_in_0_ce1),
    .t_address1(tdf8_accum_1_U0_accum_in_0_address1),
    .t_q1(products_0_t_q1)
);

td_fused_top_dataflow_in_loop_TOP_LOOP37454_accum1_out_0 #(
    .DataWidth( 16 ),
    .AddressRange( 8 ),
    .AddressWidth( 3 ))
accum1_out_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf8_accum_1_U0_ap_done),
    .i_full_n(accum1_out_0_i_full_n),
    .i_ce0(tdf8_accum_1_U0_accum_out_ce0),
    .i_we0(tdf8_accum_1_U0_accum_out_we0),
    .i_address0(tdf8_accum_1_U0_accum_out_address0),
    .i_d0(tdf8_accum_1_U0_accum_out_d0),
    .i_q0(accum1_out_0_i_q0),
    .i_ce1(tdf8_accum_1_U0_accum_out_ce1),
    .i_we1(tdf8_accum_1_U0_accum_out_we1),
    .i_address1(tdf8_accum_1_U0_accum_out_address1),
    .i_d1(tdf8_accum_1_U0_accum_out_d1),
    .t_ce(1'b1),
    .t_read(tdf8_accum_2_U0_ap_ready),
    .t_empty_n(accum1_out_0_t_empty_n),
    .t_ce0(tdf8_accum_2_U0_accum_in_ce0),
    .t_we0(1'b0),
    .t_address0(tdf8_accum_2_U0_accum_in_address0),
    .t_d0(16'd0),
    .t_q0(accum1_out_0_t_q0),
    .t_ce1(1'b0),
    .t_we1(1'b0),
    .t_address1(3'd0),
    .t_d1(16'd0)
);

td_fused_top_tdf8_get_next_ijk tdf8_get_next_ijk_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf8_get_next_ijk_U0_ap_start),
    .start_full_n(start_for_tdf8_readFilters56_U0_full_n),
    .ap_done(tdf8_get_next_ijk_U0_ap_done),
    .ap_continue(tdf8_get_next_ijk_U0_ap_continue),
    .ap_idle(tdf8_get_next_ijk_U0_ap_idle),
    .ap_ready(tdf8_get_next_ijk_U0_ap_ready),
    .start_out(tdf8_get_next_ijk_U0_start_out),
    .start_write(tdf8_get_next_ijk_U0_start_write),
    .input_indices_2_out_din(tdf8_get_next_ijk_U0_input_indices_2_out_din),
    .input_indices_2_out_full_n(input_indices_23_c_full_n),
    .input_indices_2_out_write(tdf8_get_next_ijk_U0_input_indices_2_out_write),
    .input_indices_2_out1_din(tdf8_get_next_ijk_U0_input_indices_2_out1_din),
    .input_indices_2_out1_full_n(input_indices_23_c1_full_n),
    .input_indices_2_out1_write(tdf8_get_next_ijk_U0_input_indices_2_out1_write),
    .output_indices_0_din(tdf8_get_next_ijk_U0_output_indices_0_din),
    .output_indices_0_full_n(output_indices_04_c_full_n),
    .output_indices_0_write(tdf8_get_next_ijk_U0_output_indices_0_write),
    .output_indices_1_din(tdf8_get_next_ijk_U0_output_indices_1_din),
    .output_indices_1_full_n(output_indices_15_c_full_n),
    .output_indices_1_write(tdf8_get_next_ijk_U0_output_indices_1_write),
    .resetMaximum_din(tdf8_get_next_ijk_U0_resetMaximum_din),
    .resetMaximum_full_n(resetMaximum6_c_full_n),
    .resetMaximum_write(tdf8_get_next_ijk_U0_resetMaximum_write),
    .storeOutput_din(tdf8_get_next_ijk_U0_storeOutput_din),
    .storeOutput_full_n(storeOutput7_c_full_n),
    .storeOutput_write(tdf8_get_next_ijk_U0_storeOutput_write),
    .ap_return_0(tdf8_get_next_ijk_U0_ap_return_0),
    .ap_return_1(tdf8_get_next_ijk_U0_ap_return_1)
);

td_fused_top_tdf8_readInputs57 tdf8_readInputs57_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf8_readInputs57_U0_ap_start),
    .ap_done(tdf8_readInputs57_U0_ap_done),
    .ap_continue(tdf8_readInputs57_U0_ap_continue),
    .ap_idle(tdf8_readInputs57_U0_ap_idle),
    .ap_ready(tdf8_readInputs57_U0_ap_ready),
    .in_data_address0(tdf8_readInputs57_U0_in_data_address0),
    .in_data_ce0(tdf8_readInputs57_U0_in_data_ce0),
    .in_data_q0(in_data_q0),
    .i_13(input_indices_0_dout),
    .j_13(input_indices_1_dout),
    .ifmap_vec_address0(tdf8_readInputs57_U0_ifmap_vec_address0),
    .ifmap_vec_ce0(tdf8_readInputs57_U0_ifmap_vec_ce0),
    .ifmap_vec_we0(tdf8_readInputs57_U0_ifmap_vec_we0),
    .ifmap_vec_d0(tdf8_readInputs57_U0_ifmap_vec_d0),
    .ifmap_vec_address1(tdf8_readInputs57_U0_ifmap_vec_address1),
    .ifmap_vec_ce1(tdf8_readInputs57_U0_ifmap_vec_ce1),
    .ifmap_vec_we1(tdf8_readInputs57_U0_ifmap_vec_we1),
    .ifmap_vec_d1(tdf8_readInputs57_U0_ifmap_vec_d1)
);

td_fused_top_tdf8_readFilters56 tdf8_readFilters56_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf8_readFilters56_U0_ap_start),
    .ap_done(tdf8_readFilters56_U0_ap_done),
    .ap_continue(tdf8_readFilters56_U0_ap_continue),
    .ap_idle(tdf8_readFilters56_U0_ap_idle),
    .ap_ready(tdf8_readFilters56_U0_ap_ready),
    .filter_data_address0(tdf8_readFilters56_U0_filter_data_address0),
    .filter_data_ce0(tdf8_readFilters56_U0_filter_data_ce0),
    .filter_data_q0(filter_data_q0),
    .input_indices_23_dout(input_indices_23_c_dout),
    .input_indices_23_empty_n(input_indices_23_c_empty_n),
    .input_indices_23_read(tdf8_readFilters56_U0_input_indices_23_read),
    .weight_vecs_0_address0(tdf8_readFilters56_U0_weight_vecs_0_address0),
    .weight_vecs_0_ce0(tdf8_readFilters56_U0_weight_vecs_0_ce0),
    .weight_vecs_0_we0(tdf8_readFilters56_U0_weight_vecs_0_we0),
    .weight_vecs_0_d0(tdf8_readFilters56_U0_weight_vecs_0_d0)
);

td_fused_top_tdf8_dot_product tdf8_dot_product_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf8_dot_product_U0_ap_start),
    .ap_done(tdf8_dot_product_U0_ap_done),
    .ap_continue(tdf8_dot_product_U0_ap_continue),
    .ap_idle(tdf8_dot_product_U0_ap_idle),
    .ap_ready(tdf8_dot_product_U0_ap_ready),
    .ifmap_vec_address0(tdf8_dot_product_U0_ifmap_vec_address0),
    .ifmap_vec_ce0(tdf8_dot_product_U0_ifmap_vec_ce0),
    .ifmap_vec_q0(ifmap_vec_t_q0),
    .weight_vecs_0_address0(tdf8_dot_product_U0_weight_vecs_0_address0),
    .weight_vecs_0_ce0(tdf8_dot_product_U0_weight_vecs_0_ce0),
    .weight_vecs_0_q0(weight_vecs_0_t_q0),
    .products_0_address0(tdf8_dot_product_U0_products_0_address0),
    .products_0_ce0(tdf8_dot_product_U0_products_0_ce0),
    .products_0_we0(tdf8_dot_product_U0_products_0_we0),
    .products_0_d0(tdf8_dot_product_U0_products_0_d0)
);

td_fused_top_tdf8_accum_1 tdf8_accum_1_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf8_accum_1_U0_ap_start),
    .ap_done(tdf8_accum_1_U0_ap_done),
    .ap_continue(tdf8_accum_1_U0_ap_continue),
    .ap_idle(tdf8_accum_1_U0_ap_idle),
    .ap_ready(tdf8_accum_1_U0_ap_ready),
    .accum_in_0_address0(tdf8_accum_1_U0_accum_in_0_address0),
    .accum_in_0_ce0(tdf8_accum_1_U0_accum_in_0_ce0),
    .accum_in_0_q0(products_0_t_q0),
    .accum_in_0_address1(tdf8_accum_1_U0_accum_in_0_address1),
    .accum_in_0_ce1(tdf8_accum_1_U0_accum_in_0_ce1),
    .accum_in_0_q1(products_0_t_q1),
    .accum_out_address0(tdf8_accum_1_U0_accum_out_address0),
    .accum_out_ce0(tdf8_accum_1_U0_accum_out_ce0),
    .accum_out_we0(tdf8_accum_1_U0_accum_out_we0),
    .accum_out_d0(tdf8_accum_1_U0_accum_out_d0),
    .accum_out_address1(tdf8_accum_1_U0_accum_out_address1),
    .accum_out_ce1(tdf8_accum_1_U0_accum_out_ce1),
    .accum_out_we1(tdf8_accum_1_U0_accum_out_we1),
    .accum_out_d1(tdf8_accum_1_U0_accum_out_d1)
);

td_fused_top_tdf8_accum_2 tdf8_accum_2_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf8_accum_2_U0_ap_start),
    .ap_done(tdf8_accum_2_U0_ap_done),
    .ap_continue(tdf8_accum_2_U0_ap_continue),
    .ap_idle(tdf8_accum_2_U0_ap_idle),
    .ap_ready(tdf8_accum_2_U0_ap_ready),
    .accum_in_4(tdf8_accum_2_U0_accum_in_4),
    .accum_in_4_ap_vld(tdf8_accum_2_U0_accum_in_4_ap_vld),
    .accum_in_address0(tdf8_accum_2_U0_accum_in_address0),
    .accum_in_ce0(tdf8_accum_2_U0_accum_in_ce0),
    .accum_in_q0(accum1_out_0_t_q0)
);

td_fused_top_Block_entry_proc_proc424 Block_entry_proc_proc424_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(Block_entry_proc_proc424_U0_ap_start),
    .ap_done(Block_entry_proc_proc424_U0_ap_done),
    .ap_continue(Block_entry_proc_proc424_U0_ap_continue),
    .ap_idle(Block_entry_proc_proc424_U0_ap_idle),
    .ap_ready(Block_entry_proc_proc424_U0_ap_ready),
    .tmp(tmp_channel_dout),
    .ap_return(Block_entry_proc_proc424_U0_ap_return)
);

td_fused_top_tdf8_adjust tdf8_adjust_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf8_adjust_U0_ap_start),
    .ap_done(tdf8_adjust_U0_ap_done),
    .ap_continue(tdf8_adjust_U0_ap_continue),
    .ap_idle(tdf8_adjust_U0_ap_idle),
    .ap_ready(tdf8_adjust_U0_ap_ready),
    .sums_read(sums_0_dout),
    .adjustments_address0(tdf8_adjust_U0_adjustments_address0),
    .adjustments_ce0(tdf8_adjust_U0_adjustments_ce0),
    .adjustments_q0(adjustments_q0),
    .input_indices_23_dout(input_indices_23_c1_dout),
    .input_indices_23_empty_n(input_indices_23_c1_empty_n),
    .input_indices_23_read(tdf8_adjust_U0_input_indices_23_read),
    .ap_return(tdf8_adjust_U0_ap_return)
);

td_fused_top_tdf8_poolOutputs tdf8_poolOutputs_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf8_poolOutputs_U0_ap_start),
    .ap_done(tdf8_poolOutputs_U0_ap_done),
    .ap_continue(tdf8_poolOutputs_U0_ap_continue),
    .ap_idle(tdf8_poolOutputs_U0_ap_idle),
    .ap_ready(tdf8_poolOutputs_U0_ap_ready),
    .output_indices_04_dout(output_indices_04_c_dout),
    .output_indices_04_empty_n(output_indices_04_c_empty_n),
    .output_indices_04_read(tdf8_poolOutputs_U0_output_indices_04_read),
    .output_indices_15_dout(output_indices_15_c_dout),
    .output_indices_15_empty_n(output_indices_15_c_empty_n),
    .output_indices_15_read(tdf8_poolOutputs_U0_output_indices_15_read),
    .resetMaximum6_dout(resetMaximum6_c_dout),
    .resetMaximum6_empty_n(resetMaximum6_c_empty_n),
    .resetMaximum6_read(tdf8_poolOutputs_U0_resetMaximum6_read),
    .storeOutput7_dout(storeOutput7_c_dout),
    .storeOutput7_empty_n(storeOutput7_c_empty_n),
    .storeOutput7_read(tdf8_poolOutputs_U0_storeOutput7_read),
    .p_read(outputs_0_dout),
    .out_data_address1(tdf8_poolOutputs_U0_out_data_address1),
    .out_data_ce1(tdf8_poolOutputs_U0_out_data_ce1),
    .out_data_we1(tdf8_poolOutputs_U0_out_data_we1),
    .out_data_d1(tdf8_poolOutputs_U0_out_data_d1)
);

td_fused_top_fifo_w8_d2_S_x input_indices_23_c_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(input_indices_23_c_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf8_readFilters56_U0_input_indices_23_read),
    .if_dout(input_indices_23_c_dout),
    .if_full_n(input_indices_23_c_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf8_get_next_ijk_U0_input_indices_2_out_write),
    .if_din(tdf8_get_next_ijk_U0_input_indices_2_out_din)
);

td_fused_top_fifo_w8_d7_S input_indices_23_c1_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(input_indices_23_c1_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf8_adjust_U0_input_indices_23_read),
    .if_dout(input_indices_23_c1_dout),
    .if_full_n(input_indices_23_c1_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf8_get_next_ijk_U0_input_indices_2_out1_write),
    .if_din(tdf8_get_next_ijk_U0_input_indices_2_out1_din)
);

td_fused_top_fifo_w4_d8_S_x output_indices_04_c_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(output_indices_04_c_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf8_poolOutputs_U0_output_indices_04_read),
    .if_dout(output_indices_04_c_dout),
    .if_full_n(output_indices_04_c_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf8_get_next_ijk_U0_output_indices_0_write),
    .if_din(tdf8_get_next_ijk_U0_output_indices_0_din)
);

td_fused_top_fifo_w8_d8_S output_indices_15_c_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(output_indices_15_c_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf8_poolOutputs_U0_output_indices_15_read),
    .if_dout(output_indices_15_c_dout),
    .if_full_n(output_indices_15_c_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf8_get_next_ijk_U0_output_indices_1_write),
    .if_din(tdf8_get_next_ijk_U0_output_indices_1_din)
);

td_fused_top_fifo_w1_d8_S_x0 resetMaximum6_c_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(resetMaximum6_c_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf8_poolOutputs_U0_resetMaximum6_read),
    .if_dout(resetMaximum6_c_dout),
    .if_full_n(resetMaximum6_c_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf8_get_next_ijk_U0_resetMaximum_write),
    .if_din(resetMaximum6_c_din)
);

td_fused_top_fifo_w1_d8_S_x0 storeOutput7_c_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(storeOutput7_c_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf8_poolOutputs_U0_storeOutput7_read),
    .if_dout(storeOutput7_c_dout),
    .if_full_n(storeOutput7_c_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf8_get_next_ijk_U0_storeOutput_write),
    .if_din(storeOutput7_c_din)
);

td_fused_top_fifo_w16_d2_S_x5 input_indices_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(input_indices_0_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf8_readInputs57_U0_ap_ready),
    .if_dout(input_indices_0_dout),
    .if_full_n(input_indices_0_full_n),
    .if_write_ce(1'b1),
    .if_write(ap_channel_done_input_indices_0),
    .if_din(tdf8_get_next_ijk_U0_ap_return_0)
);

td_fused_top_fifo_w16_d2_S_x5 input_indices_1_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(input_indices_1_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf8_readInputs57_U0_ap_ready),
    .if_dout(input_indices_1_dout),
    .if_full_n(input_indices_1_full_n),
    .if_write_ce(1'b1),
    .if_write(ap_channel_done_input_indices_1),
    .if_din(tdf8_get_next_ijk_U0_ap_return_1)
);

td_fused_top_fifo_w16_d2_S_x5 tmp_channel_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(tmp_channel_empty_n),
    .if_read_ce(1'b1),
    .if_read(Block_entry_proc_proc424_U0_ap_ready),
    .if_dout(tmp_channel_dout),
    .if_full_n(tmp_channel_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf8_accum_2_U0_ap_done),
    .if_din(tdf8_accum_2_U0_accum_in_4)
);

td_fused_top_fifo_w16_d2_S_x5 sums_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(sums_0_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf8_adjust_U0_ap_ready),
    .if_dout(sums_0_dout),
    .if_full_n(sums_0_full_n),
    .if_write_ce(1'b1),
    .if_write(Block_entry_proc_proc424_U0_ap_done),
    .if_din(Block_entry_proc_proc424_U0_ap_return)
);

td_fused_top_fifo_w16_d2_S_x5 outputs_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(outputs_0_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf8_poolOutputs_U0_ap_ready),
    .if_dout(outputs_0_dout),
    .if_full_n(outputs_0_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf8_adjust_U0_ap_done),
    .if_din(tdf8_adjust_U0_ap_return)
);

td_fused_top_start_for_tdf8_readFilters56_U0 start_for_tdf8_readFilters56_U0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(start_for_tdf8_readFilters56_U0_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf8_readFilters56_U0_ap_ready),
    .if_dout(start_for_tdf8_readFilters56_U0_dout),
    .if_full_n(start_for_tdf8_readFilters56_U0_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf8_get_next_ijk_U0_start_write),
    .if_din(start_for_tdf8_readFilters56_U0_din)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_sync_reg_channel_write_input_indices_0 <= 1'b0;
    end else begin
        if (((tdf8_get_next_ijk_U0_ap_done & tdf8_get_next_ijk_U0_ap_continue) == 1'b1)) begin
            ap_sync_reg_channel_write_input_indices_0 <= 1'b0;
        end else begin
            ap_sync_reg_channel_write_input_indices_0 <= ap_sync_channel_write_input_indices_0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_sync_reg_channel_write_input_indices_1 <= 1'b0;
    end else begin
        if (((tdf8_get_next_ijk_U0_ap_done & tdf8_get_next_ijk_U0_ap_continue) == 1'b1)) begin
            ap_sync_reg_channel_write_input_indices_1 <= 1'b0;
        end else begin
            ap_sync_reg_channel_write_input_indices_1 <= ap_sync_channel_write_input_indices_1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_sync_reg_tdf8_get_next_ijk_U0_ap_ready <= 1'b0;
    end else begin
        if (((ap_sync_ready & ap_start) == 1'b1)) begin
            ap_sync_reg_tdf8_get_next_ijk_U0_ap_ready <= 1'b0;
        end else begin
            ap_sync_reg_tdf8_get_next_ijk_U0_ap_ready <= ap_sync_tdf8_get_next_ijk_U0_ap_ready;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_sync_reg_tdf8_readInputs57_U0_ap_ready <= 1'b0;
    end else begin
        if (((ap_sync_ready & ap_start) == 1'b1)) begin
            ap_sync_reg_tdf8_readInputs57_U0_ap_ready <= 1'b0;
        end else begin
            ap_sync_reg_tdf8_readInputs57_U0_ap_ready <= ap_sync_tdf8_readInputs57_U0_ap_ready;
        end
    end
end

assign Block_entry_proc_proc424_U0_ap_continue = sums_0_full_n;

assign Block_entry_proc_proc424_U0_ap_start = tmp_channel_empty_n;

assign Block_entry_proc_proc424_U0_start_full_n = 1'b1;

assign Block_entry_proc_proc424_U0_start_write = 1'b0;

assign adjustments_address0 = tdf8_adjust_U0_adjustments_address0;

assign adjustments_address1 = 8'd0;

assign adjustments_ce0 = tdf8_adjust_U0_adjustments_ce0;

assign adjustments_ce1 = 1'b0;

assign adjustments_d0 = 48'd0;

assign adjustments_d1 = 48'd0;

assign adjustments_we0 = 1'b0;

assign adjustments_we1 = 1'b0;

assign ap_channel_done_accum1_out_0 = tdf8_accum_1_U0_ap_done;

assign ap_channel_done_ifmap_vec = tdf8_readInputs57_U0_ap_done;

assign ap_channel_done_input_indices_0 = (tdf8_get_next_ijk_U0_ap_done & (ap_sync_reg_channel_write_input_indices_0 ^ 1'b1));

assign ap_channel_done_input_indices_1 = (tdf8_get_next_ijk_U0_ap_done & (ap_sync_reg_channel_write_input_indices_1 ^ 1'b1));

assign ap_channel_done_outputs_0 = tdf8_adjust_U0_ap_done;

assign ap_channel_done_products_0 = tdf8_dot_product_U0_ap_done;

assign ap_channel_done_sums_0 = Block_entry_proc_proc424_U0_ap_done;

assign ap_channel_done_tmp_channel = tdf8_accum_2_U0_ap_done;

assign ap_channel_done_weight_vecs_0 = tdf8_readFilters56_U0_ap_done;

assign ap_done = tdf8_poolOutputs_U0_ap_done;

assign ap_idle = (tdf8_readInputs57_U0_ap_idle & tdf8_readFilters56_U0_ap_idle & tdf8_poolOutputs_U0_ap_idle & tdf8_get_next_ijk_U0_ap_idle & tdf8_dot_product_U0_ap_idle & tdf8_adjust_U0_ap_idle & tdf8_accum_2_U0_ap_idle & tdf8_accum_1_U0_ap_idle & (outputs_0_empty_n ^ 1'b1) & (sums_0_empty_n ^ 1'b1) & (tmp_channel_empty_n ^ 1'b1) & (input_indices_1_empty_n ^ 1'b1) & (input_indices_0_empty_n ^ 1'b1) & (products_0_t_empty_n ^ 1'b1) & (weight_vecs_0_t_empty_n ^ 1'b1) & (ifmap_vec_t_empty_n ^ 1'b1) & (1'b1 ^ accum1_out_0_t_empty_n) & Block_entry_proc_proc424_U0_ap_idle);

assign ap_ready = ap_sync_ready;

assign ap_sync_channel_write_input_indices_0 = ((input_indices_0_full_n & ap_channel_done_input_indices_0) | ap_sync_reg_channel_write_input_indices_0);

assign ap_sync_channel_write_input_indices_1 = ((input_indices_1_full_n & ap_channel_done_input_indices_1) | ap_sync_reg_channel_write_input_indices_1);

assign ap_sync_continue = ap_continue;

assign ap_sync_done = tdf8_poolOutputs_U0_ap_done;

assign ap_sync_ready = (ap_sync_tdf8_readInputs57_U0_ap_ready & ap_sync_tdf8_get_next_ijk_U0_ap_ready);

assign ap_sync_tdf8_get_next_ijk_U0_ap_ready = (tdf8_get_next_ijk_U0_ap_ready | ap_sync_reg_tdf8_get_next_ijk_U0_ap_ready);

assign ap_sync_tdf8_readInputs57_U0_ap_ready = (tdf8_readInputs57_U0_ap_ready | ap_sync_reg_tdf8_readInputs57_U0_ap_ready);

assign filter_data_address0 = tdf8_readFilters56_U0_filter_data_address0;

assign filter_data_address1 = 17'd0;

assign filter_data_ce0 = tdf8_readFilters56_U0_filter_data_ce0;

assign filter_data_ce1 = 1'b0;

assign filter_data_d0 = 16'd0;

assign filter_data_d1 = 16'd0;

assign filter_data_we0 = 1'b0;

assign filter_data_we1 = 1'b0;

assign in_data_address0 = tdf8_readInputs57_U0_in_data_address0;

assign in_data_address1 = 13'd0;

assign in_data_ce0 = tdf8_readInputs57_U0_in_data_ce0;

assign in_data_ce1 = 1'b0;

assign in_data_d0 = 64'd0;

assign in_data_d1 = 64'd0;

assign in_data_read = tdf8_readInputs57_U0_in_data_write;

assign in_data_we0 = 1'b0;

assign in_data_we1 = 1'b0;

assign out_data_address0 = 14'd0;

assign out_data_address1 = tdf8_poolOutputs_U0_out_data_address1;

assign out_data_ce0 = 1'b0;

assign out_data_ce1 = tdf8_poolOutputs_U0_out_data_ce1;

assign out_data_d0 = 64'd0;

assign out_data_d1 = tdf8_poolOutputs_U0_out_data_d1;

assign out_data_we0 = 1'b0;

assign out_data_we1 = tdf8_poolOutputs_U0_out_data_we1;

assign out_data_write = tdf8_poolOutputs_U0_out_data_write;

assign products_0_t_d1 = 16'd0;

assign products_0_t_we1 = 1'b0;

assign resetMaximum6_c_din = tdf8_get_next_ijk_U0_resetMaximum_din;

assign start_for_tdf8_readFilters56_U0_din = 1'b1;

assign storeOutput7_c_din = tdf8_get_next_ijk_U0_storeOutput_din;

assign tdf8_accum_1_U0_accum_out_full_n = accum1_out_0_i_full_n;

assign tdf8_accum_1_U0_ap_continue = accum1_out_0_i_full_n;

assign tdf8_accum_1_U0_ap_start = products_0_t_empty_n;

assign tdf8_accum_1_U0_start_full_n = 1'b1;

assign tdf8_accum_1_U0_start_write = 1'b0;

assign tdf8_accum_2_U0_ap_continue = tmp_channel_full_n;

assign tdf8_accum_2_U0_ap_start = accum1_out_0_t_empty_n;

assign tdf8_accum_2_U0_start_full_n = 1'b1;

assign tdf8_accum_2_U0_start_write = 1'b0;

assign tdf8_adjust_U0_ap_continue = outputs_0_full_n;

assign tdf8_adjust_U0_ap_start = sums_0_empty_n;

assign tdf8_adjust_U0_start_full_n = 1'b1;

assign tdf8_adjust_U0_start_write = 1'b0;

assign tdf8_dot_product_U0_ap_continue = products_0_i_full_n;

assign tdf8_dot_product_U0_ap_start = (weight_vecs_0_t_empty_n & ifmap_vec_t_empty_n);

assign tdf8_dot_product_U0_products_0_full_n = products_0_i_full_n;

assign tdf8_dot_product_U0_start_full_n = 1'b1;

assign tdf8_dot_product_U0_start_write = 1'b0;

assign tdf8_get_next_ijk_U0_ap_continue = (ap_sync_channel_write_input_indices_1 & ap_sync_channel_write_input_indices_0);

assign tdf8_get_next_ijk_U0_ap_start = ((ap_sync_reg_tdf8_get_next_ijk_U0_ap_ready ^ 1'b1) & ap_start);

assign tdf8_poolOutputs_U0_ap_continue = ap_continue;

assign tdf8_poolOutputs_U0_ap_start = outputs_0_empty_n;

assign tdf8_poolOutputs_U0_out_data_full_n = out_data_full_n;

assign tdf8_poolOutputs_U0_out_data_write = 1'b0;

assign tdf8_poolOutputs_U0_start_full_n = 1'b1;

assign tdf8_poolOutputs_U0_start_write = 1'b0;

assign tdf8_readFilters56_U0_ap_continue = weight_vecs_0_i_full_n;

assign tdf8_readFilters56_U0_ap_start = start_for_tdf8_readFilters56_U0_empty_n;

assign tdf8_readFilters56_U0_start_full_n = 1'b1;

assign tdf8_readFilters56_U0_start_write = 1'b0;

assign tdf8_readFilters56_U0_weight_vecs_0_full_n = weight_vecs_0_i_full_n;

assign tdf8_readInputs57_U0_ap_continue = ifmap_vec_i_full_n;

assign tdf8_readInputs57_U0_ap_start = (input_indices_1_empty_n & input_indices_0_empty_n & (ap_sync_reg_tdf8_readInputs57_U0_ap_ready ^ 1'b1) & ap_start);

assign tdf8_readInputs57_U0_ifmap_vec_full_n = ifmap_vec_i_full_n;

assign tdf8_readInputs57_U0_in_data_full_n = in_data_empty_n;

assign tdf8_readInputs57_U0_in_data_write = 1'b0;

assign tdf8_readInputs57_U0_start_full_n = 1'b1;

assign tdf8_readInputs57_U0_start_write = 1'b0;

endmodule //td_fused_top_dataflow_in_loop_TOP_LOOP37454
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37454_weight_vecs_0_memcore_ram (addr0, ce0, d0, we0, q0, addr1, ce1, d1, we1, q1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 10;
parameter MEM_SIZE = 576;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
output reg[DWIDTH-1:0] q1;
input clk;

reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];




always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1) 
            ram[addr1] <= d1; 
        q1 <= ram[addr1];
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37454_weight_vecs_0_memcore(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    q0,
    address1,
    ce1,
    we1,
    d1,
    q1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd576;
parameter AddressWidth = 32'd10;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;
output[DataWidth - 1:0] q1;



td_fused_top_dataflow_in_loop_TOP_LOOP37454_weight_vecs_0_memcore_ram td_fused_top_dataflow_in_loop_TOP_LOOP37454_weight_vecs_0_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 ),
    .q1( q1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_dataflow_in_loop_TOP_LOOP37454_weight_vecs_0
#(parameter
    DataWidth    = 16,
    AddressRange = 32,
    AddressWidth = 9,
    BufferCount  = 2,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire                    i_we0,
    input  wire [AddressWidth-1:0] i_address0,
    input  wire [DataWidth-1:0]    i_d0,
    output wire [DataWidth-1:0]    i_q0,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire                    t_we0,
    input  wire [AddressWidth-1:0] t_address0,
    input  wire [DataWidth-1:0]    t_d0,
    output wire [DataWidth-1:0]    t_q0
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
wire [AddressWidth+IndexWidth-1:0]   memcore_iaddr;
wire [AddressWidth+IndexWidth-1:0]   memcore_taddr;

//------------------------Instantiation------------------
assign memcore_iaddr = {i_address0, iptr};
assign memcore_taddr = {t_address0, tptr};
td_fused_top_dataflow_in_loop_TOP_LOOP37454_weight_vecs_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP37454_weight_vecs_0_memcore_U (
    .reset    ( reset ),
    .clk      ( clk ),
    .address0 ( memcore_iaddr ),
    .ce0      ( i_ce0 ),
    .we0      ( i_we0),
    .d0       ( i_d0 ),
    .q0       ( i_q0 ),
    .address1 ( memcore_taddr ),
    .ce1      ( t_ce0 ),
    .we1      ( t_we0),
    .d1       ( t_d0 ),
    .q1       ( t_q0 )

);

//------------------------Body---------------------------

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37548_accum1_out_0_memcore_ram (addr0, ce0, d0, we0, q0, addr1, ce1, d1, we1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 3;
parameter MEM_SIZE = 8;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
input clk;

reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];




always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1) 
            ram[addr1] <= d1; 
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37548_accum1_out_0_memcore(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    q0,
    address1,
    ce1,
    we1,
    d1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd8;
parameter AddressWidth = 32'd3;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;



td_fused_top_dataflow_in_loop_TOP_LOOP37548_accum1_out_0_memcore_ram td_fused_top_dataflow_in_loop_TOP_LOOP37548_accum1_out_0_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_dataflow_in_loop_TOP_LOOP37548_accum1_out_0
#(parameter
    DataWidth    = 16,
    AddressRange = 32,
    AddressWidth = 3,
    BufferCount  = 2,
    MemLatency   = 1,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire                    i_we0,
    input  wire [AddressWidth-1:0] i_address0,
    input  wire [DataWidth-1:0]    i_d0,
    output wire [DataWidth-1:0]    i_q0,
    input  wire                    i_ce1,
    input  wire                    i_we1,
    input  wire [AddressWidth-1:0] i_address1,
    input  wire [DataWidth-1:0]    i_d1,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire                    t_we0,
    input  wire [AddressWidth-1:0] t_address0,
    input  wire [DataWidth-1:0]    t_d0,
    output wire [DataWidth-1:0]    t_q0,
    input  wire                    t_ce1,
    input  wire                    t_we1,
    input  wire [AddressWidth-1:0] t_address1,
    input  wire [DataWidth-1:0]    t_d1
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth-1:0]   prev_iptr    = 1'b0; // previous initiator index
reg  [IndexWidth-1:0]   prev_tptr    = 1'b0; // previous target index
reg  [DataWidth-1:0]    reg_q0      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid0    = 1'b0; // buffer has valid data
reg  [DataWidth-1:0]    reg_q1      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid1    = 1'b0; // buffer has valid data
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
// buffer signals
wire [BufferCount-1:0] buf_ce0;
wire [BufferCount-1:0] buf_we0;
wire [AddressWidth-1:0] buf_a0_0, buf_a0_1;
wire [DataWidth-1:0] buf_d0_0, buf_d0_1;
wire [DataWidth-1:0] buf_q0_0, buf_q0_1;
wire [BufferCount-1:0] buf_ce1;
wire [BufferCount-1:0] buf_we1;
wire [AddressWidth-1:0] buf_a1_0, buf_a1_1;
wire [DataWidth-1:0] buf_d1_0, buf_d1_1;
//------------------------Instantiation------------------
//genvar i;
        td_fused_top_dataflow_in_loop_TOP_LOOP37548_accum1_out_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP37548_accum1_out_0_memcore_U_0 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_0 ),
            .ce0      ( buf_ce0[ 0 ] ),
            .we0      ( buf_we0[ 0 ] ),
            .d0       ( buf_d0_0 ),
            .q0       ( buf_q0_0 ),
            .address1 ( buf_a1_0 ),
            .ce1      ( buf_ce1[ 0 ] ),
            .we1      ( buf_we1[ 0 ] ),
            .d1       ( buf_d1_0 )
        );
        td_fused_top_dataflow_in_loop_TOP_LOOP37548_accum1_out_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP37548_accum1_out_0_memcore_U_1 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_1 ),
            .ce0      ( buf_ce0[ 1 ] ),
            .we0      ( buf_we0[ 1 ] ),
            .d0       ( buf_d0_1 ),
            .q0       ( buf_q0_1 ),
            .address1 ( buf_a1_1 ),
            .ce1      ( buf_ce1[ 1 ] ),
            .we1      ( buf_we1[ 1 ] ),
            .d1       ( buf_d1_1 )
        );

//++++++++++++++++++++++++buffer signals+++++++++++++++++
        assign buf_ce0[ 0 ] = (tptr ==  0  && empty_n) ? t_ce0
                             : (iptr ==  0 ) ? i_ce0 : 1'b0;
        assign buf_a0_0  = (tptr ==  0  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 0 ] = (tptr ==  0  && empty_n)  ? t_we0
                             : (iptr ==  0 ) ? i_we0 : 1'b0;
        assign buf_d0_0  = (tptr ==  0  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 0 ] = (tptr ==  0  && empty_n) ? t_ce1
                             : (iptr ==  0 ) ? i_ce1 : 1'b0;
        assign buf_a1_0  = (tptr ==  0  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 0 ] = (tptr ==  0  && empty_n)  ? t_we1
                             : (iptr ==  0 ) ? i_we1 : 1'b0;
        assign buf_d1_0  = (tptr ==  0  && empty_n) ? t_d1       : i_d1;
        assign buf_ce0[ 1 ] = (tptr ==  1  && empty_n) ? t_ce0
                             : (iptr ==  1 ) ? i_ce0 : 1'b0;
        assign buf_a0_1  = (tptr ==  1  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 1 ] = (tptr ==  1  && empty_n)  ? t_we0
                             : (iptr ==  1 ) ? i_we0 : 1'b0;
        assign buf_d0_1  = (tptr ==  1  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 1 ] = (tptr ==  1  && empty_n) ? t_ce1
                             : (iptr ==  1 ) ? i_ce1 : 1'b0;
        assign buf_a1_1  = (tptr ==  1  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 1 ] = (tptr ==  1  && empty_n)  ? t_we1
                             : (iptr ==  1 ) ? i_we1 : 1'b0;
        assign buf_d1_1  = (tptr ==  1  && empty_n) ? t_d1       : i_d1;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//------------------------Body---------------------------
assign i_q0      = (prev_iptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign t_q0      = reg_valid0 ? reg_q0 : (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// prev_iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_iptr <= 1'b0;
    else begin
        prev_iptr <= iptr;
    end
end

// prev_tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_tptr <= 1'b0;
    else begin
        prev_tptr <= tptr;
    end
end

// reg_q0 and reg_valid0
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q0     <= 1'b0;
        reg_valid0 <= 1'b0;
    end else if (!t_ce0 && !reg_valid0) begin
        reg_q0     <= (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
        reg_valid0 <= 1'b1;
    end else if (t_ce0) begin
        reg_valid0 <= 1'b0;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37548_ifmap_vec_memcore_ram (addr0, ce0, d0, we0, q0, addr1, ce1, d1, we1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 9;
parameter MEM_SIZE = 288;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
input clk;

reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];




always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1) 
            ram[addr1] <= d1; 
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37548_ifmap_vec_memcore(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    q0,
    address1,
    ce1,
    we1,
    d1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd288;
parameter AddressWidth = 32'd9;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;



td_fused_top_dataflow_in_loop_TOP_LOOP37548_ifmap_vec_memcore_ram td_fused_top_dataflow_in_loop_TOP_LOOP37548_ifmap_vec_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_dataflow_in_loop_TOP_LOOP37548_ifmap_vec
#(parameter
    DataWidth    = 16,
    AddressRange = 32,
    AddressWidth = 9,
    BufferCount  = 2,
    MemLatency   = 1,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire                    i_we0,
    input  wire [AddressWidth-1:0] i_address0,
    input  wire [DataWidth-1:0]    i_d0,
    output wire [DataWidth-1:0]    i_q0,
    input  wire                    i_ce1,
    input  wire                    i_we1,
    input  wire [AddressWidth-1:0] i_address1,
    input  wire [DataWidth-1:0]    i_d1,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire                    t_we0,
    input  wire [AddressWidth-1:0] t_address0,
    input  wire [DataWidth-1:0]    t_d0,
    output wire [DataWidth-1:0]    t_q0,
    input  wire                    t_ce1,
    input  wire                    t_we1,
    input  wire [AddressWidth-1:0] t_address1,
    input  wire [DataWidth-1:0]    t_d1
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth-1:0]   prev_iptr    = 1'b0; // previous initiator index
reg  [IndexWidth-1:0]   prev_tptr    = 1'b0; // previous target index
reg  [DataWidth-1:0]    reg_q0      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid0    = 1'b0; // buffer has valid data
reg  [DataWidth-1:0]    reg_q1      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid1    = 1'b0; // buffer has valid data
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
// buffer signals
wire [BufferCount-1:0] buf_ce0;
wire [BufferCount-1:0] buf_we0;
wire [AddressWidth-1:0] buf_a0_0, buf_a0_1;
wire [DataWidth-1:0] buf_d0_0, buf_d0_1;
wire [DataWidth-1:0] buf_q0_0, buf_q0_1;
wire [BufferCount-1:0] buf_ce1;
wire [BufferCount-1:0] buf_we1;
wire [AddressWidth-1:0] buf_a1_0, buf_a1_1;
wire [DataWidth-1:0] buf_d1_0, buf_d1_1;
//------------------------Instantiation------------------
//genvar i;
        td_fused_top_dataflow_in_loop_TOP_LOOP37548_ifmap_vec_memcore td_fused_top_dataflow_in_loop_TOP_LOOP37548_ifmap_vec_memcore_U_0 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_0 ),
            .ce0      ( buf_ce0[ 0 ] ),
            .we0      ( buf_we0[ 0 ] ),
            .d0       ( buf_d0_0 ),
            .q0       ( buf_q0_0 ),
            .address1 ( buf_a1_0 ),
            .ce1      ( buf_ce1[ 0 ] ),
            .we1      ( buf_we1[ 0 ] ),
            .d1       ( buf_d1_0 )
        );
        td_fused_top_dataflow_in_loop_TOP_LOOP37548_ifmap_vec_memcore td_fused_top_dataflow_in_loop_TOP_LOOP37548_ifmap_vec_memcore_U_1 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_1 ),
            .ce0      ( buf_ce0[ 1 ] ),
            .we0      ( buf_we0[ 1 ] ),
            .d0       ( buf_d0_1 ),
            .q0       ( buf_q0_1 ),
            .address1 ( buf_a1_1 ),
            .ce1      ( buf_ce1[ 1 ] ),
            .we1      ( buf_we1[ 1 ] ),
            .d1       ( buf_d1_1 )
        );

//++++++++++++++++++++++++buffer signals+++++++++++++++++
        assign buf_ce0[ 0 ] = (tptr ==  0  && empty_n) ? t_ce0
                             : (iptr ==  0 ) ? i_ce0 : 1'b0;
        assign buf_a0_0  = (tptr ==  0  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 0 ] = (tptr ==  0  && empty_n)  ? t_we0
                             : (iptr ==  0 ) ? i_we0 : 1'b0;
        assign buf_d0_0  = (tptr ==  0  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 0 ] = (tptr ==  0  && empty_n) ? t_ce1
                             : (iptr ==  0 ) ? i_ce1 : 1'b0;
        assign buf_a1_0  = (tptr ==  0  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 0 ] = (tptr ==  0  && empty_n)  ? t_we1
                             : (iptr ==  0 ) ? i_we1 : 1'b0;
        assign buf_d1_0  = (tptr ==  0  && empty_n) ? t_d1       : i_d1;
        assign buf_ce0[ 1 ] = (tptr ==  1  && empty_n) ? t_ce0
                             : (iptr ==  1 ) ? i_ce0 : 1'b0;
        assign buf_a0_1  = (tptr ==  1  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 1 ] = (tptr ==  1  && empty_n)  ? t_we0
                             : (iptr ==  1 ) ? i_we0 : 1'b0;
        assign buf_d0_1  = (tptr ==  1  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 1 ] = (tptr ==  1  && empty_n) ? t_ce1
                             : (iptr ==  1 ) ? i_ce1 : 1'b0;
        assign buf_a1_1  = (tptr ==  1  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 1 ] = (tptr ==  1  && empty_n)  ? t_we1
                             : (iptr ==  1 ) ? i_we1 : 1'b0;
        assign buf_d1_1  = (tptr ==  1  && empty_n) ? t_d1       : i_d1;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//------------------------Body---------------------------
assign i_q0      = (prev_iptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign t_q0      = reg_valid0 ? reg_q0 : (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// prev_iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_iptr <= 1'b0;
    else begin
        prev_iptr <= iptr;
    end
end

// prev_tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_tptr <= 1'b0;
    else begin
        prev_tptr <= tptr;
    end
end

// reg_q0 and reg_valid0
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q0     <= 1'b0;
        reg_valid0 <= 1'b0;
    end else if (!t_ce0 && !reg_valid0) begin
        reg_q0     <= (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
        reg_valid0 <= 1'b1;
    end else if (t_ce0) begin
        reg_valid0 <= 1'b0;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37548_l2_products_memcore_ram (addr0, ce0, d0, we0, q0, addr1, ce1, d1, we1, q1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
output reg[DWIDTH-1:0] q1;
input clk;

 reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];




always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1) 
            ram[addr1] <= d1; 
        q1 <= ram[addr1];
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37548_l2_products_memcore(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    q0,
    address1,
    ce1,
    we1,
    d1,
    q1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;
output[DataWidth - 1:0] q1;



td_fused_top_dataflow_in_loop_TOP_LOOP37548_l2_products_memcore_ram td_fused_top_dataflow_in_loop_TOP_LOOP37548_l2_products_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 ),
    .q1( q1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_dataflow_in_loop_TOP_LOOP37548_l2_products
#(parameter
    DataWidth    = 16,
    AddressRange = 32,
    AddressWidth = 5,
    BufferCount  = 2,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire                    i_we0,
    input  wire [AddressWidth-1:0] i_address0,
    input  wire [DataWidth-1:0]    i_d0,
    output wire [DataWidth-1:0]    i_q0,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire                    t_we0,
    input  wire [AddressWidth-1:0] t_address0,
    input  wire [DataWidth-1:0]    t_d0,
    output wire [DataWidth-1:0]    t_q0
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
wire [AddressWidth+IndexWidth-1:0]   memcore_iaddr;
wire [AddressWidth+IndexWidth-1:0]   memcore_taddr;

//------------------------Instantiation------------------
assign memcore_iaddr = {i_address0, iptr};
assign memcore_taddr = {t_address0, tptr};
td_fused_top_dataflow_in_loop_TOP_LOOP37548_l2_products_memcore td_fused_top_dataflow_in_loop_TOP_LOOP37548_l2_products_memcore_U (
    .reset    ( reset ),
    .clk      ( clk ),
    .address0 ( memcore_iaddr ),
    .ce0      ( i_ce0 ),
    .we0      ( i_we0),
    .d0       ( i_d0 ),
    .q0       ( i_q0 ),
    .address1 ( memcore_taddr ),
    .ce1      ( t_ce0 ),
    .we1      ( t_we0),
    .d1       ( t_d0 ),
    .q1       ( t_q0 )

);

//------------------------Body---------------------------

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37548_products_0_memcore_ram (addr0, ce0, d0, we0, q0, addr1, ce1, q1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 9;
parameter MEM_SIZE = 288;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
output reg[DWIDTH-1:0] q1;
input clk;

reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];




always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        q1 <= ram[addr1];
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37548_products_0_memcore(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    q0,
    address1,
    ce1,
    q1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd288;
parameter AddressWidth = 32'd9;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
output[DataWidth - 1:0] q1;



td_fused_top_dataflow_in_loop_TOP_LOOP37548_products_0_memcore_ram td_fused_top_dataflow_in_loop_TOP_LOOP37548_products_0_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .q1( q1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_dataflow_in_loop_TOP_LOOP37548_products_0
#(parameter
    DataWidth    = 16,
    AddressRange = 32,
    AddressWidth = 9,
    BufferCount  = 2,
    MemLatency   = 1,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire                    i_we0,
    input  wire [AddressWidth-1:0] i_address0,
    input  wire [DataWidth-1:0]    i_d0,
    output wire [DataWidth-1:0]    i_q0,
    input  wire                    i_ce1,
    input  wire [AddressWidth-1:0] i_address1,
    output wire [DataWidth-1:0]    i_q1,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire                    t_we0,
    input  wire [AddressWidth-1:0] t_address0,
    input  wire [DataWidth-1:0]    t_d0,
    output wire [DataWidth-1:0]    t_q0,
    input  wire                    t_ce1,
    input  wire [AddressWidth-1:0] t_address1,
    output wire [DataWidth-1:0]    t_q1
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth-1:0]   prev_iptr    = 1'b0; // previous initiator index
reg  [IndexWidth-1:0]   prev_tptr    = 1'b0; // previous target index
reg  [DataWidth-1:0]    reg_q0      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid0    = 1'b0; // buffer has valid data
reg  [DataWidth-1:0]    reg_q1      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid1    = 1'b0; // buffer has valid data
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
// buffer signals
wire [BufferCount-1:0] buf_ce0;
wire [BufferCount-1:0] buf_we0;
wire [AddressWidth-1:0] buf_a0_0, buf_a0_1;
wire [DataWidth-1:0] buf_d0_0, buf_d0_1;
wire [DataWidth-1:0] buf_q0_0, buf_q0_1;
wire [BufferCount-1:0] buf_ce1;
wire [AddressWidth-1:0] buf_a1_0, buf_a1_1;
wire [DataWidth-1:0] buf_q1_0, buf_q1_1;
//------------------------Instantiation------------------
//genvar i;
        td_fused_top_dataflow_in_loop_TOP_LOOP37548_products_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP37548_products_0_memcore_U_0 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_0 ),
            .ce0      ( buf_ce0[ 0 ] ),
            .we0      ( buf_we0[ 0 ] ),
            .d0       ( buf_d0_0 ),
            .q0       ( buf_q0_0 ),
            .address1 ( buf_a1_0 ),
            .ce1      ( buf_ce1[ 0 ] ),
            .q1       ( buf_q1_0 )
        );
        td_fused_top_dataflow_in_loop_TOP_LOOP37548_products_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP37548_products_0_memcore_U_1 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_1 ),
            .ce0      ( buf_ce0[ 1 ] ),
            .we0      ( buf_we0[ 1 ] ),
            .d0       ( buf_d0_1 ),
            .q0       ( buf_q0_1 ),
            .address1 ( buf_a1_1 ),
            .ce1      ( buf_ce1[ 1 ] ),
            .q1       ( buf_q1_1 )
        );

//++++++++++++++++++++++++buffer signals+++++++++++++++++
        assign buf_ce0[ 0 ] = (tptr ==  0  && empty_n) ? t_ce0
                             : (iptr ==  0 ) ? i_ce0 : 1'b0;
        assign buf_a0_0  = (tptr ==  0  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 0 ] = (tptr ==  0  && empty_n)  ? t_we0
                             : (iptr ==  0 ) ? i_we0 : 1'b0;
        assign buf_d0_0  = (tptr ==  0  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 0 ] = (tptr ==  0  && empty_n) ? t_ce1
                             : (iptr ==  0 ) ? i_ce1 : 1'b0;
        assign buf_a1_0  = (tptr ==  0  && empty_n) ?  t_address1 : i_address1;
        assign buf_ce0[ 1 ] = (tptr ==  1  && empty_n) ? t_ce0
                             : (iptr ==  1 ) ? i_ce0 : 1'b0;
        assign buf_a0_1  = (tptr ==  1  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 1 ] = (tptr ==  1  && empty_n)  ? t_we0
                             : (iptr ==  1 ) ? i_we0 : 1'b0;
        assign buf_d0_1  = (tptr ==  1  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 1 ] = (tptr ==  1  && empty_n) ? t_ce1
                             : (iptr ==  1 ) ? i_ce1 : 1'b0;
        assign buf_a1_1  = (tptr ==  1  && empty_n) ?  t_address1 : i_address1;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//------------------------Body---------------------------
assign i_q0      = (prev_iptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign t_q0      = reg_valid0 ? reg_q0 : (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign i_q1      = (prev_iptr == 1'b1 ? buf_q1_1 : buf_q1_0);
assign t_q1      = reg_valid1 ? reg_q1 : (prev_tptr == 1'b1 ? buf_q1_1 : buf_q1_0);

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// prev_iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_iptr <= 1'b0;
    else begin
        prev_iptr <= iptr;
    end
end

// prev_tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_tptr <= 1'b0;
    else begin
        prev_tptr <= tptr;
    end
end

// reg_q0 and reg_valid0
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q0     <= 1'b0;
        reg_valid0 <= 1'b0;
    end else if (!t_ce0 && !reg_valid0) begin
        reg_q0     <= (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
        reg_valid0 <= 1'b1;
    end else if (t_ce0) begin
        reg_valid0 <= 1'b0;
    end
end

// reg_q1 and reg_valid1
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q1     <= 1'b0;
        reg_valid1 <= 1'b0;
    end else if (!t_ce1 && !reg_valid1) begin
        reg_q1     <= (prev_tptr == 1'b1 ? buf_q1_1 : buf_q1_0);
        reg_valid1 <= 1'b1;
    end else if (t_ce1) begin
        reg_valid1 <= 1'b0;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_dataflow_in_loop_TOP_LOOP37548 (
        ap_clk,
        ap_rst,
        in_data_address0,
        in_data_ce0,
        in_data_d0,
        in_data_q0,
        in_data_we0,
        in_data_address1,
        in_data_ce1,
        in_data_d1,
        in_data_q1,
        in_data_we1,
        l1_filter_data_address0,
        l1_filter_data_ce0,
        l1_filter_data_d0,
        l1_filter_data_q0,
        l1_filter_data_we0,
        l1_filter_data_address1,
        l1_filter_data_ce1,
        l1_filter_data_d1,
        l1_filter_data_q1,
        l1_filter_data_we1,
        l1_adjustments_address0,
        l1_adjustments_ce0,
        l1_adjustments_d0,
        l1_adjustments_q0,
        l1_adjustments_we0,
        l1_adjustments_address1,
        l1_adjustments_ce1,
        l1_adjustments_d1,
        l1_adjustments_q1,
        l1_adjustments_we1,
        l2_filter_data_address0,
        l2_filter_data_ce0,
        l2_filter_data_d0,
        l2_filter_data_q0,
        l2_filter_data_we0,
        l2_filter_data_address1,
        l2_filter_data_ce1,
        l2_filter_data_d1,
        l2_filter_data_q1,
        l2_filter_data_we1,
        out_data_address0,
        out_data_ce0,
        out_data_d0,
        out_data_q0,
        out_data_we0,
        out_data_address1,
        out_data_ce1,
        out_data_d1,
        out_data_q1,
        out_data_we1,
        l2_adjustments_address0,
        l2_adjustments_ce0,
        l2_adjustments_d0,
        l2_adjustments_q0,
        l2_adjustments_we0,
        l2_adjustments_address1,
        l2_adjustments_ce1,
        l2_adjustments_d1,
        l2_adjustments_q1,
        l2_adjustments_we1,
        ap_start,
        in_data_empty_n,
        in_data_read,
        out_data_full_n,
        out_data_write,
        ap_done,
        ap_ready,
        ap_idle,
        ap_continue
);


input   ap_clk;
input   ap_rst;
output  [12:0] in_data_address0;
output   in_data_ce0;
output  [63:0] in_data_d0;
input  [63:0] in_data_q0;
output   in_data_we0;
output  [12:0] in_data_address1;
output   in_data_ce1;
output  [63:0] in_data_d1;
input  [63:0] in_data_q1;
output   in_data_we1;
output  [16:0] l1_filter_data_address0;
output   l1_filter_data_ce0;
output  [15:0] l1_filter_data_d0;
input  [15:0] l1_filter_data_q0;
output   l1_filter_data_we0;
output  [16:0] l1_filter_data_address1;
output   l1_filter_data_ce1;
output  [15:0] l1_filter_data_d1;
input  [15:0] l1_filter_data_q1;
output   l1_filter_data_we1;
output  [7:0] l1_adjustments_address0;
output   l1_adjustments_ce0;
output  [47:0] l1_adjustments_d0;
input  [47:0] l1_adjustments_q0;
output   l1_adjustments_we0;
output  [7:0] l1_adjustments_address1;
output   l1_adjustments_ce1;
output  [47:0] l1_adjustments_d1;
input  [47:0] l1_adjustments_q1;
output   l1_adjustments_we1;
output  [12:0] l2_filter_data_address0;
output   l2_filter_data_ce0;
output  [15:0] l2_filter_data_d0;
input  [15:0] l2_filter_data_q0;
output   l2_filter_data_we0;
output  [12:0] l2_filter_data_address1;
output   l2_filter_data_ce1;
output  [15:0] l2_filter_data_d1;
input  [15:0] l2_filter_data_q1;
output   l2_filter_data_we1;
output  [12:0] out_data_address0;
output   out_data_ce0;
output  [63:0] out_data_d0;
input  [63:0] out_data_q0;
output   out_data_we0;
output  [12:0] out_data_address1;
output   out_data_ce1;
output  [63:0] out_data_d1;
input  [63:0] out_data_q1;
output   out_data_we1;
output  [4:0] l2_adjustments_address0;
output   l2_adjustments_ce0;
output  [47:0] l2_adjustments_d0;
input  [47:0] l2_adjustments_q0;
output   l2_adjustments_we0;
output  [4:0] l2_adjustments_address1;
output   l2_adjustments_ce1;
output  [47:0] l2_adjustments_d1;
input  [47:0] l2_adjustments_q1;
output   l2_adjustments_we1;
input   ap_start;
input   in_data_empty_n;
output   in_data_read;
input   out_data_full_n;
output   out_data_write;
output   ap_done;
output   ap_ready;
output   ap_idle;
input   ap_continue;

wire   [15:0] ifmap_vec_i_q0;
wire   [15:0] ifmap_vec_t_q0;
wire   [15:0] weight_vecs_0_i_q0;
wire   [15:0] weight_vecs_0_t_q0;
wire   [15:0] products_0_i_q0;
wire   [15:0] products_0_i_q1;
wire   [15:0] products_0_t_q0;
wire   [15:0] products_0_t_q1;
wire   [15:0] accum1_out_0_i_q0;
wire   [15:0] accum1_out_0_t_q0;
wire   [15:0] l2_products_i_q0;
wire   [15:0] l2_products_t_q0;
wire    tdf7_get_next_ijk_U0_ap_start;
wire    tdf7_get_next_ijk_U0_ap_done;
wire    tdf7_get_next_ijk_U0_ap_continue;
wire    tdf7_get_next_ijk_U0_ap_idle;
wire    tdf7_get_next_ijk_U0_ap_ready;
wire    tdf7_get_next_ijk_U0_start_out;
wire    tdf7_get_next_ijk_U0_start_write;
wire   [15:0] tdf7_get_next_ijk_U0_indices_0_din;
wire    tdf7_get_next_ijk_U0_indices_0_write;
wire   [15:0] tdf7_get_next_ijk_U0_indices_1_din;
wire    tdf7_get_next_ijk_U0_indices_1_write;
wire   [7:0] tdf7_get_next_ijk_U0_indices_2_out_din;
wire    tdf7_get_next_ijk_U0_indices_2_out_write;
wire   [12:0] tdf7_get_next_ijk_U0_indices_2_out1_din;
wire    tdf7_get_next_ijk_U0_indices_2_out1_write;
wire    tdf7_get_next_ijk_U0_write_r_din;
wire    tdf7_get_next_ijk_U0_write_r_write;
wire    tdf7_readInputs53_U0_ap_start;
wire    tdf7_readInputs53_U0_ap_done;
wire    tdf7_readInputs53_U0_ap_continue;
wire    tdf7_readInputs53_U0_ap_idle;
wire    tdf7_readInputs53_U0_ap_ready;
wire   [12:0] tdf7_readInputs53_U0_in_data_address0;
wire    tdf7_readInputs53_U0_in_data_ce0;
wire    tdf7_readInputs53_U0_indices_01_read;
wire    tdf7_readInputs53_U0_indices_12_read;
wire   [8:0] tdf7_readInputs53_U0_ifmap_vec_address0;
wire    tdf7_readInputs53_U0_ifmap_vec_ce0;
wire    tdf7_readInputs53_U0_ifmap_vec_we0;
wire   [15:0] tdf7_readInputs53_U0_ifmap_vec_d0;
wire   [8:0] tdf7_readInputs53_U0_ifmap_vec_address1;
wire    tdf7_readInputs53_U0_ifmap_vec_ce1;
wire    tdf7_readInputs53_U0_ifmap_vec_we1;
wire   [15:0] tdf7_readInputs53_U0_ifmap_vec_d1;
wire   [4:0] tdf7_readInputs53_U0_indices_01_out_din;
wire    tdf7_readInputs53_U0_indices_01_out_write;
wire   [9:0] tdf7_readInputs53_U0_indices_12_out_din;
wire    tdf7_readInputs53_U0_indices_12_out_write;
wire    tdf7_readInputs53_U0_in_data_full_n;
wire    tdf7_readInputs53_U0_in_data_write;
wire    ap_channel_done_ifmap_vec;
wire    tdf7_readInputs53_U0_ifmap_vec_full_n;
wire    tdf7_readFilters52_U0_ap_start;
wire    tdf7_readFilters52_U0_ap_done;
wire    tdf7_readFilters52_U0_ap_continue;
wire    tdf7_readFilters52_U0_ap_idle;
wire    tdf7_readFilters52_U0_ap_ready;
wire   [16:0] tdf7_readFilters52_U0_filter_data_address0;
wire    tdf7_readFilters52_U0_filter_data_ce0;
wire    tdf7_readFilters52_U0_indices_23_read;
wire   [8:0] tdf7_readFilters52_U0_weight_vecs_0_address0;
wire    tdf7_readFilters52_U0_weight_vecs_0_ce0;
wire    tdf7_readFilters52_U0_weight_vecs_0_we0;
wire   [15:0] tdf7_readFilters52_U0_weight_vecs_0_d0;
wire    ap_channel_done_weight_vecs_0;
wire    tdf7_readFilters52_U0_weight_vecs_0_full_n;
wire    tdf7_dot_product_U0_ap_start;
wire    tdf7_dot_product_U0_ap_done;
wire    tdf7_dot_product_U0_ap_continue;
wire    tdf7_dot_product_U0_ap_idle;
wire    tdf7_dot_product_U0_ap_ready;
wire   [8:0] tdf7_dot_product_U0_ifmap_vec_address0;
wire    tdf7_dot_product_U0_ifmap_vec_ce0;
wire   [8:0] tdf7_dot_product_U0_weight_vecs_0_address0;
wire    tdf7_dot_product_U0_weight_vecs_0_ce0;
wire   [8:0] tdf7_dot_product_U0_products_0_address0;
wire    tdf7_dot_product_U0_products_0_ce0;
wire    tdf7_dot_product_U0_products_0_we0;
wire   [15:0] tdf7_dot_product_U0_products_0_d0;
wire    ap_channel_done_products_0;
wire    tdf7_dot_product_U0_products_0_full_n;
wire    tdf7_accum_1_U0_ap_start;
wire    tdf7_accum_1_U0_ap_done;
wire    tdf7_accum_1_U0_ap_continue;
wire    tdf7_accum_1_U0_ap_idle;
wire    tdf7_accum_1_U0_ap_ready;
wire   [8:0] tdf7_accum_1_U0_accum_in_0_address0;
wire    tdf7_accum_1_U0_accum_in_0_ce0;
wire   [8:0] tdf7_accum_1_U0_accum_in_0_address1;
wire    tdf7_accum_1_U0_accum_in_0_ce1;
wire   [2:0] tdf7_accum_1_U0_accum_out_address0;
wire    tdf7_accum_1_U0_accum_out_ce0;
wire    tdf7_accum_1_U0_accum_out_we0;
wire   [15:0] tdf7_accum_1_U0_accum_out_d0;
wire   [2:0] tdf7_accum_1_U0_accum_out_address1;
wire    tdf7_accum_1_U0_accum_out_ce1;
wire    tdf7_accum_1_U0_accum_out_we1;
wire   [15:0] tdf7_accum_1_U0_accum_out_d1;
wire    ap_channel_done_accum1_out_0;
wire    tdf7_accum_1_U0_accum_out_full_n;
wire    tdf7_accum_2_U0_ap_start;
wire    tdf7_accum_2_U0_ap_done;
wire    tdf7_accum_2_U0_ap_continue;
wire    tdf7_accum_2_U0_ap_idle;
wire    tdf7_accum_2_U0_ap_ready;
wire   [15:0] tdf7_accum_2_U0_accum_in_6;
wire    tdf7_accum_2_U0_accum_in_6_ap_vld;
wire   [2:0] tdf7_accum_2_U0_accum_in_address0;
wire    tdf7_accum_2_U0_accum_in_ce0;
wire    ap_channel_done_tmp_channel;
wire    tmp_channel_full_n;
wire    Block_entry_proc_proc419_U0_ap_start;
wire    Block_entry_proc_proc419_U0_ap_done;
wire    Block_entry_proc_proc419_U0_ap_continue;
wire    Block_entry_proc_proc419_U0_ap_idle;
wire    Block_entry_proc_proc419_U0_ap_ready;
wire   [15:0] Block_entry_proc_proc419_U0_ap_return;
wire    ap_channel_done_sums_0;
wire    sums_0_full_n;
wire    tdf7_adjust_U0_ap_start;
wire    tdf7_adjust_U0_ap_done;
wire    tdf7_adjust_U0_ap_continue;
wire    tdf7_adjust_U0_ap_idle;
wire    tdf7_adjust_U0_ap_ready;
wire   [7:0] tdf7_adjust_U0_adjustments_address0;
wire    tdf7_adjust_U0_adjustments_ce0;
wire    tdf7_adjust_U0_indices_23_read;
wire   [12:0] tdf7_adjust_U0_indices_23_out_din;
wire    tdf7_adjust_U0_indices_23_out_write;
wire   [15:0] tdf7_adjust_U0_ap_return;
wire    ap_channel_done_intermediate_fmaps_0;
wire    intermediate_fmaps_0_full_n;
wire    tdf7_l2_multiply50_U0_ap_start;
wire    tdf7_l2_multiply50_U0_ap_done;
wire    tdf7_l2_multiply50_U0_ap_continue;
wire    tdf7_l2_multiply50_U0_ap_idle;
wire    tdf7_l2_multiply50_U0_ap_ready;
wire   [12:0] tdf7_l2_multiply50_U0_l2_filter_data_address0;
wire    tdf7_l2_multiply50_U0_l2_filter_data_ce0;
wire   [4:0] tdf7_l2_multiply50_U0_l2_products_address0;
wire    tdf7_l2_multiply50_U0_l2_products_ce0;
wire    tdf7_l2_multiply50_U0_l2_products_we0;
wire   [15:0] tdf7_l2_multiply50_U0_l2_products_d0;
wire    tdf7_l2_multiply50_U0_indices_23_read;
wire    ap_channel_done_l2_products;
wire    tdf7_l2_multiply50_U0_l2_products_full_n;
wire    tdf7_l2_writeOutputs_149_U0_ap_start;
wire    tdf7_l2_writeOutputs_149_U0_ap_done;
wire    tdf7_l2_writeOutputs_149_U0_ap_continue;
wire    tdf7_l2_writeOutputs_149_U0_ap_idle;
wire    tdf7_l2_writeOutputs_149_U0_ap_ready;
wire    tdf7_l2_writeOutputs_149_U0_indices_01_read;
wire    tdf7_l2_writeOutputs_149_U0_indices_12_read;
wire    tdf7_l2_writeOutputs_149_U0_write4_read;
wire   [4:0] tdf7_l2_writeOutputs_149_U0_l2_partial_sums_address0;
wire    tdf7_l2_writeOutputs_149_U0_l2_partial_sums_ce0;
wire   [12:0] tdf7_l2_writeOutputs_149_U0_out_data_address1;
wire    tdf7_l2_writeOutputs_149_U0_out_data_ce1;
wire    tdf7_l2_writeOutputs_149_U0_out_data_we1;
wire   [63:0] tdf7_l2_writeOutputs_149_U0_out_data_d1;
wire   [4:0] tdf7_l2_writeOutputs_149_U0_l2_adjustments_address0;
wire    tdf7_l2_writeOutputs_149_U0_l2_adjustments_ce0;
wire    tdf7_l2_writeOutputs_149_U0_out_data_full_n;
wire    tdf7_l2_writeOutputs_149_U0_out_data_write;
wire    ap_sync_continue;
wire    ifmap_vec_i_full_n;
wire    ifmap_vec_t_empty_n;
wire    weight_vecs_0_i_full_n;
wire    weight_vecs_0_t_empty_n;
wire    products_0_i_full_n;
wire    products_0_t_empty_n;
wire   [15:0] products_0_t_d1;
wire    products_0_t_we1;
wire    accum1_out_0_i_full_n;
wire    accum1_out_0_t_empty_n;
wire    l2_products_i_full_n;
wire    l2_products_t_empty_n;
wire    indices_01_c_full_n;
wire   [15:0] indices_01_c_dout;
wire    indices_01_c_empty_n;
wire    indices_12_c_full_n;
wire   [15:0] indices_12_c_dout;
wire    indices_12_c_empty_n;
wire    indices_23_c_full_n;
wire   [7:0] indices_23_c_dout;
wire    indices_23_c_empty_n;
wire    indices_23_c1_full_n;
wire   [12:0] indices_23_c1_dout;
wire    indices_23_c1_empty_n;
wire   [0:0] write4_c_din;
wire    write4_c_full_n;
wire   [0:0] write4_c_dout;
wire    write4_c_empty_n;
wire    indices_01_c2_full_n;
wire   [4:0] indices_01_c2_dout;
wire    indices_01_c2_empty_n;
wire    indices_12_c3_full_n;
wire   [9:0] indices_12_c3_dout;
wire    indices_12_c3_empty_n;
wire   [15:0] tmp_channel_dout;
wire    tmp_channel_empty_n;
wire   [15:0] sums_0_dout;
wire    sums_0_empty_n;
wire    indices_23_c4_full_n;
wire   [12:0] indices_23_c4_dout;
wire    indices_23_c4_empty_n;
wire   [15:0] intermediate_fmaps_0_dout;
wire    intermediate_fmaps_0_empty_n;
wire    ap_sync_done;
wire    ap_sync_ready;
reg    ap_sync_reg_tdf7_get_next_ijk_U0_ap_ready;
wire    ap_sync_tdf7_get_next_ijk_U0_ap_ready;
reg    ap_sync_reg_tdf7_readInputs53_U0_ap_ready;
wire    ap_sync_tdf7_readInputs53_U0_ap_ready;
wire   [0:0] start_for_tdf7_readFilters52_U0_din;
wire    start_for_tdf7_readFilters52_U0_full_n;
wire   [0:0] start_for_tdf7_readFilters52_U0_dout;
wire    start_for_tdf7_readFilters52_U0_empty_n;
wire    tdf7_readInputs53_U0_start_full_n;
wire    tdf7_readInputs53_U0_start_write;
wire    tdf7_readFilters52_U0_start_full_n;
wire    tdf7_readFilters52_U0_start_write;
wire    tdf7_dot_product_U0_start_full_n;
wire    tdf7_dot_product_U0_start_write;
wire    tdf7_accum_1_U0_start_full_n;
wire    tdf7_accum_1_U0_start_write;
wire    tdf7_accum_2_U0_start_full_n;
wire    tdf7_accum_2_U0_start_write;
wire    Block_entry_proc_proc419_U0_start_full_n;
wire    Block_entry_proc_proc419_U0_start_write;
wire    tdf7_adjust_U0_start_full_n;
wire    tdf7_adjust_U0_start_write;
wire    tdf7_l2_multiply50_U0_start_full_n;
wire    tdf7_l2_multiply50_U0_start_write;
wire    tdf7_l2_writeOutputs_149_U0_start_full_n;
wire    tdf7_l2_writeOutputs_149_U0_start_write;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_sync_reg_tdf7_get_next_ijk_U0_ap_ready = 1'b0;
#0 ap_sync_reg_tdf7_readInputs53_U0_ap_ready = 1'b0;
end

td_fused_top_dataflow_in_loop_TOP_LOOP37548_ifmap_vec #(
    .DataWidth( 16 ),
    .AddressRange( 288 ),
    .AddressWidth( 9 ))
ifmap_vec_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf7_readInputs53_U0_ap_done),
    .i_full_n(ifmap_vec_i_full_n),
    .i_ce0(tdf7_readInputs53_U0_ifmap_vec_ce0),
    .i_we0(tdf7_readInputs53_U0_ifmap_vec_we0),
    .i_address0(tdf7_readInputs53_U0_ifmap_vec_address0),
    .i_d0(tdf7_readInputs53_U0_ifmap_vec_d0),
    .i_q0(ifmap_vec_i_q0),
    .i_ce1(tdf7_readInputs53_U0_ifmap_vec_ce1),
    .i_we1(tdf7_readInputs53_U0_ifmap_vec_we1),
    .i_address1(tdf7_readInputs53_U0_ifmap_vec_address1),
    .i_d1(tdf7_readInputs53_U0_ifmap_vec_d1),
    .t_ce(1'b1),
    .t_read(tdf7_dot_product_U0_ap_ready),
    .t_empty_n(ifmap_vec_t_empty_n),
    .t_ce0(tdf7_dot_product_U0_ifmap_vec_ce0),
    .t_we0(1'b0),
    .t_address0(tdf7_dot_product_U0_ifmap_vec_address0),
    .t_d0(16'd0),
    .t_q0(ifmap_vec_t_q0),
    .t_ce1(1'b0),
    .t_we1(1'b0),
    .t_address1(9'd0),
    .t_d1(16'd0)
);

td_fused_top_dataflow_in_loop_TOP_LOOP37548_weight_vecs_0 #(
    .DataWidth( 16 ),
    .AddressRange( 288 ),
    .AddressWidth( 9 ))
weight_vecs_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf7_readFilters52_U0_ap_done),
    .i_full_n(weight_vecs_0_i_full_n),
    .i_ce0(tdf7_readFilters52_U0_weight_vecs_0_ce0),
    .i_we0(tdf7_readFilters52_U0_weight_vecs_0_we0),
    .i_address0(tdf7_readFilters52_U0_weight_vecs_0_address0),
    .i_d0(tdf7_readFilters52_U0_weight_vecs_0_d0),
    .i_q0(weight_vecs_0_i_q0),
    .t_ce(1'b1),
    .t_read(tdf7_dot_product_U0_ap_ready),
    .t_empty_n(weight_vecs_0_t_empty_n),
    .t_ce0(tdf7_dot_product_U0_weight_vecs_0_ce0),
    .t_we0(1'b0),
    .t_address0(tdf7_dot_product_U0_weight_vecs_0_address0),
    .t_d0(16'd0),
    .t_q0(weight_vecs_0_t_q0)
);

td_fused_top_dataflow_in_loop_TOP_LOOP37548_products_0 #(
    .DataWidth( 16 ),
    .AddressRange( 288 ),
    .AddressWidth( 9 ))
products_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf7_dot_product_U0_ap_done),
    .i_full_n(products_0_i_full_n),
    .i_ce0(tdf7_dot_product_U0_products_0_ce0),
    .i_we0(tdf7_dot_product_U0_products_0_we0),
    .i_address0(tdf7_dot_product_U0_products_0_address0),
    .i_d0(tdf7_dot_product_U0_products_0_d0),
    .i_q0(products_0_i_q0),
    .i_ce1(1'b0),
    .i_address1(9'd0),
    .i_q1(products_0_i_q1),
    .t_ce(1'b1),
    .t_read(tdf7_accum_1_U0_ap_ready),
    .t_empty_n(products_0_t_empty_n),
    .t_ce0(tdf7_accum_1_U0_accum_in_0_ce0),
    .t_we0(1'b0),
    .t_address0(tdf7_accum_1_U0_accum_in_0_address0),
    .t_d0(16'd0),
    .t_q0(products_0_t_q0),
    .t_ce1(tdf7_accum_1_U0_accum_in_0_ce1),
    .t_address1(tdf7_accum_1_U0_accum_in_0_address1),
    .t_q1(products_0_t_q1)
);

td_fused_top_dataflow_in_loop_TOP_LOOP37548_accum1_out_0 #(
    .DataWidth( 16 ),
    .AddressRange( 8 ),
    .AddressWidth( 3 ))
accum1_out_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf7_accum_1_U0_ap_done),
    .i_full_n(accum1_out_0_i_full_n),
    .i_ce0(tdf7_accum_1_U0_accum_out_ce0),
    .i_we0(tdf7_accum_1_U0_accum_out_we0),
    .i_address0(tdf7_accum_1_U0_accum_out_address0),
    .i_d0(tdf7_accum_1_U0_accum_out_d0),
    .i_q0(accum1_out_0_i_q0),
    .i_ce1(tdf7_accum_1_U0_accum_out_ce1),
    .i_we1(tdf7_accum_1_U0_accum_out_we1),
    .i_address1(tdf7_accum_1_U0_accum_out_address1),
    .i_d1(tdf7_accum_1_U0_accum_out_d1),
    .t_ce(1'b1),
    .t_read(tdf7_accum_2_U0_ap_ready),
    .t_empty_n(accum1_out_0_t_empty_n),
    .t_ce0(tdf7_accum_2_U0_accum_in_ce0),
    .t_we0(1'b0),
    .t_address0(tdf7_accum_2_U0_accum_in_address0),
    .t_d0(16'd0),
    .t_q0(accum1_out_0_t_q0),
    .t_ce1(1'b0),
    .t_we1(1'b0),
    .t_address1(3'd0),
    .t_d1(16'd0)
);

td_fused_top_dataflow_in_loop_TOP_LOOP37548_l2_products #(
    .DataWidth( 16 ),
    .AddressRange( 32 ),
    .AddressWidth( 5 ))
l2_products_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf7_l2_multiply50_U0_ap_done),
    .i_full_n(l2_products_i_full_n),
    .i_ce0(tdf7_l2_multiply50_U0_l2_products_ce0),
    .i_we0(tdf7_l2_multiply50_U0_l2_products_we0),
    .i_address0(tdf7_l2_multiply50_U0_l2_products_address0),
    .i_d0(tdf7_l2_multiply50_U0_l2_products_d0),
    .i_q0(l2_products_i_q0),
    .t_ce(1'b1),
    .t_read(tdf7_l2_writeOutputs_149_U0_ap_ready),
    .t_empty_n(l2_products_t_empty_n),
    .t_ce0(tdf7_l2_writeOutputs_149_U0_l2_partial_sums_ce0),
    .t_we0(1'b0),
    .t_address0(tdf7_l2_writeOutputs_149_U0_l2_partial_sums_address0),
    .t_d0(16'd0),
    .t_q0(l2_products_t_q0)
);

td_fused_top_tdf7_get_next_ijk tdf7_get_next_ijk_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf7_get_next_ijk_U0_ap_start),
    .start_full_n(start_for_tdf7_readFilters52_U0_full_n),
    .ap_done(tdf7_get_next_ijk_U0_ap_done),
    .ap_continue(tdf7_get_next_ijk_U0_ap_continue),
    .ap_idle(tdf7_get_next_ijk_U0_ap_idle),
    .ap_ready(tdf7_get_next_ijk_U0_ap_ready),
    .start_out(tdf7_get_next_ijk_U0_start_out),
    .start_write(tdf7_get_next_ijk_U0_start_write),
    .indices_0_din(tdf7_get_next_ijk_U0_indices_0_din),
    .indices_0_full_n(indices_01_c_full_n),
    .indices_0_write(tdf7_get_next_ijk_U0_indices_0_write),
    .indices_1_din(tdf7_get_next_ijk_U0_indices_1_din),
    .indices_1_full_n(indices_12_c_full_n),
    .indices_1_write(tdf7_get_next_ijk_U0_indices_1_write),
    .indices_2_out_din(tdf7_get_next_ijk_U0_indices_2_out_din),
    .indices_2_out_full_n(indices_23_c_full_n),
    .indices_2_out_write(tdf7_get_next_ijk_U0_indices_2_out_write),
    .indices_2_out1_din(tdf7_get_next_ijk_U0_indices_2_out1_din),
    .indices_2_out1_full_n(indices_23_c1_full_n),
    .indices_2_out1_write(tdf7_get_next_ijk_U0_indices_2_out1_write),
    .write_r_din(tdf7_get_next_ijk_U0_write_r_din),
    .write_r_full_n(write4_c_full_n),
    .write_r_write(tdf7_get_next_ijk_U0_write_r_write)
);

td_fused_top_tdf7_readInputs53 tdf7_readInputs53_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf7_readInputs53_U0_ap_start),
    .ap_done(tdf7_readInputs53_U0_ap_done),
    .ap_continue(tdf7_readInputs53_U0_ap_continue),
    .ap_idle(tdf7_readInputs53_U0_ap_idle),
    .ap_ready(tdf7_readInputs53_U0_ap_ready),
    .in_data_address0(tdf7_readInputs53_U0_in_data_address0),
    .in_data_ce0(tdf7_readInputs53_U0_in_data_ce0),
    .in_data_q0(in_data_q0),
    .indices_01_dout(indices_01_c_dout),
    .indices_01_empty_n(indices_01_c_empty_n),
    .indices_01_read(tdf7_readInputs53_U0_indices_01_read),
    .indices_12_dout(indices_12_c_dout),
    .indices_12_empty_n(indices_12_c_empty_n),
    .indices_12_read(tdf7_readInputs53_U0_indices_12_read),
    .ifmap_vec_address0(tdf7_readInputs53_U0_ifmap_vec_address0),
    .ifmap_vec_ce0(tdf7_readInputs53_U0_ifmap_vec_ce0),
    .ifmap_vec_we0(tdf7_readInputs53_U0_ifmap_vec_we0),
    .ifmap_vec_d0(tdf7_readInputs53_U0_ifmap_vec_d0),
    .ifmap_vec_address1(tdf7_readInputs53_U0_ifmap_vec_address1),
    .ifmap_vec_ce1(tdf7_readInputs53_U0_ifmap_vec_ce1),
    .ifmap_vec_we1(tdf7_readInputs53_U0_ifmap_vec_we1),
    .ifmap_vec_d1(tdf7_readInputs53_U0_ifmap_vec_d1),
    .indices_01_out_din(tdf7_readInputs53_U0_indices_01_out_din),
    .indices_01_out_full_n(indices_01_c2_full_n),
    .indices_01_out_write(tdf7_readInputs53_U0_indices_01_out_write),
    .indices_12_out_din(tdf7_readInputs53_U0_indices_12_out_din),
    .indices_12_out_full_n(indices_12_c3_full_n),
    .indices_12_out_write(tdf7_readInputs53_U0_indices_12_out_write)
);

td_fused_top_tdf7_readFilters52 tdf7_readFilters52_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf7_readFilters52_U0_ap_start),
    .ap_done(tdf7_readFilters52_U0_ap_done),
    .ap_continue(tdf7_readFilters52_U0_ap_continue),
    .ap_idle(tdf7_readFilters52_U0_ap_idle),
    .ap_ready(tdf7_readFilters52_U0_ap_ready),
    .filter_data_address0(tdf7_readFilters52_U0_filter_data_address0),
    .filter_data_ce0(tdf7_readFilters52_U0_filter_data_ce0),
    .filter_data_q0(l1_filter_data_q0),
    .indices_23_dout(indices_23_c_dout),
    .indices_23_empty_n(indices_23_c_empty_n),
    .indices_23_read(tdf7_readFilters52_U0_indices_23_read),
    .weight_vecs_0_address0(tdf7_readFilters52_U0_weight_vecs_0_address0),
    .weight_vecs_0_ce0(tdf7_readFilters52_U0_weight_vecs_0_ce0),
    .weight_vecs_0_we0(tdf7_readFilters52_U0_weight_vecs_0_we0),
    .weight_vecs_0_d0(tdf7_readFilters52_U0_weight_vecs_0_d0)
);

td_fused_top_tdf7_dot_product tdf7_dot_product_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf7_dot_product_U0_ap_start),
    .ap_done(tdf7_dot_product_U0_ap_done),
    .ap_continue(tdf7_dot_product_U0_ap_continue),
    .ap_idle(tdf7_dot_product_U0_ap_idle),
    .ap_ready(tdf7_dot_product_U0_ap_ready),
    .ifmap_vec_address0(tdf7_dot_product_U0_ifmap_vec_address0),
    .ifmap_vec_ce0(tdf7_dot_product_U0_ifmap_vec_ce0),
    .ifmap_vec_q0(ifmap_vec_t_q0),
    .weight_vecs_0_address0(tdf7_dot_product_U0_weight_vecs_0_address0),
    .weight_vecs_0_ce0(tdf7_dot_product_U0_weight_vecs_0_ce0),
    .weight_vecs_0_q0(weight_vecs_0_t_q0),
    .products_0_address0(tdf7_dot_product_U0_products_0_address0),
    .products_0_ce0(tdf7_dot_product_U0_products_0_ce0),
    .products_0_we0(tdf7_dot_product_U0_products_0_we0),
    .products_0_d0(tdf7_dot_product_U0_products_0_d0)
);

td_fused_top_tdf7_accum_1 tdf7_accum_1_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf7_accum_1_U0_ap_start),
    .ap_done(tdf7_accum_1_U0_ap_done),
    .ap_continue(tdf7_accum_1_U0_ap_continue),
    .ap_idle(tdf7_accum_1_U0_ap_idle),
    .ap_ready(tdf7_accum_1_U0_ap_ready),
    .accum_in_0_address0(tdf7_accum_1_U0_accum_in_0_address0),
    .accum_in_0_ce0(tdf7_accum_1_U0_accum_in_0_ce0),
    .accum_in_0_q0(products_0_t_q0),
    .accum_in_0_address1(tdf7_accum_1_U0_accum_in_0_address1),
    .accum_in_0_ce1(tdf7_accum_1_U0_accum_in_0_ce1),
    .accum_in_0_q1(products_0_t_q1),
    .accum_out_address0(tdf7_accum_1_U0_accum_out_address0),
    .accum_out_ce0(tdf7_accum_1_U0_accum_out_ce0),
    .accum_out_we0(tdf7_accum_1_U0_accum_out_we0),
    .accum_out_d0(tdf7_accum_1_U0_accum_out_d0),
    .accum_out_address1(tdf7_accum_1_U0_accum_out_address1),
    .accum_out_ce1(tdf7_accum_1_U0_accum_out_ce1),
    .accum_out_we1(tdf7_accum_1_U0_accum_out_we1),
    .accum_out_d1(tdf7_accum_1_U0_accum_out_d1)
);

td_fused_top_tdf7_accum_2 tdf7_accum_2_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf7_accum_2_U0_ap_start),
    .ap_done(tdf7_accum_2_U0_ap_done),
    .ap_continue(tdf7_accum_2_U0_ap_continue),
    .ap_idle(tdf7_accum_2_U0_ap_idle),
    .ap_ready(tdf7_accum_2_U0_ap_ready),
    .accum_in_6(tdf7_accum_2_U0_accum_in_6),
    .accum_in_6_ap_vld(tdf7_accum_2_U0_accum_in_6_ap_vld),
    .accum_in_address0(tdf7_accum_2_U0_accum_in_address0),
    .accum_in_ce0(tdf7_accum_2_U0_accum_in_ce0),
    .accum_in_q0(accum1_out_0_t_q0)
);

td_fused_top_Block_entry_proc_proc419 Block_entry_proc_proc419_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(Block_entry_proc_proc419_U0_ap_start),
    .ap_done(Block_entry_proc_proc419_U0_ap_done),
    .ap_continue(Block_entry_proc_proc419_U0_ap_continue),
    .ap_idle(Block_entry_proc_proc419_U0_ap_idle),
    .ap_ready(Block_entry_proc_proc419_U0_ap_ready),
    .tmp(tmp_channel_dout),
    .ap_return(Block_entry_proc_proc419_U0_ap_return)
);

td_fused_top_tdf7_adjust tdf7_adjust_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf7_adjust_U0_ap_start),
    .ap_done(tdf7_adjust_U0_ap_done),
    .ap_continue(tdf7_adjust_U0_ap_continue),
    .ap_idle(tdf7_adjust_U0_ap_idle),
    .ap_ready(tdf7_adjust_U0_ap_ready),
    .sums_read(sums_0_dout),
    .adjustments_address0(tdf7_adjust_U0_adjustments_address0),
    .adjustments_ce0(tdf7_adjust_U0_adjustments_ce0),
    .adjustments_q0(l1_adjustments_q0),
    .indices_23_dout(indices_23_c1_dout),
    .indices_23_empty_n(indices_23_c1_empty_n),
    .indices_23_read(tdf7_adjust_U0_indices_23_read),
    .indices_23_out_din(tdf7_adjust_U0_indices_23_out_din),
    .indices_23_out_full_n(indices_23_c4_full_n),
    .indices_23_out_write(tdf7_adjust_U0_indices_23_out_write),
    .ap_return(tdf7_adjust_U0_ap_return)
);

td_fused_top_tdf7_l2_multiply50 tdf7_l2_multiply50_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf7_l2_multiply50_U0_ap_start),
    .ap_done(tdf7_l2_multiply50_U0_ap_done),
    .ap_continue(tdf7_l2_multiply50_U0_ap_continue),
    .ap_idle(tdf7_l2_multiply50_U0_ap_idle),
    .ap_ready(tdf7_l2_multiply50_U0_ap_ready),
    .intermediate_fmaps_read(intermediate_fmaps_0_dout),
    .l2_filter_data_address0(tdf7_l2_multiply50_U0_l2_filter_data_address0),
    .l2_filter_data_ce0(tdf7_l2_multiply50_U0_l2_filter_data_ce0),
    .l2_filter_data_q0(l2_filter_data_q0),
    .l2_products_address0(tdf7_l2_multiply50_U0_l2_products_address0),
    .l2_products_ce0(tdf7_l2_multiply50_U0_l2_products_ce0),
    .l2_products_we0(tdf7_l2_multiply50_U0_l2_products_we0),
    .l2_products_d0(tdf7_l2_multiply50_U0_l2_products_d0),
    .indices_23_dout(indices_23_c4_dout),
    .indices_23_empty_n(indices_23_c4_empty_n),
    .indices_23_read(tdf7_l2_multiply50_U0_indices_23_read)
);

td_fused_top_tdf7_l2_writeOutputs_149 tdf7_l2_writeOutputs_149_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf7_l2_writeOutputs_149_U0_ap_start),
    .ap_done(tdf7_l2_writeOutputs_149_U0_ap_done),
    .ap_continue(tdf7_l2_writeOutputs_149_U0_ap_continue),
    .ap_idle(tdf7_l2_writeOutputs_149_U0_ap_idle),
    .ap_ready(tdf7_l2_writeOutputs_149_U0_ap_ready),
    .indices_01_dout(indices_01_c2_dout),
    .indices_01_empty_n(indices_01_c2_empty_n),
    .indices_01_read(tdf7_l2_writeOutputs_149_U0_indices_01_read),
    .indices_12_dout(indices_12_c3_dout),
    .indices_12_empty_n(indices_12_c3_empty_n),
    .indices_12_read(tdf7_l2_writeOutputs_149_U0_indices_12_read),
    .write4_dout(write4_c_dout),
    .write4_empty_n(write4_c_empty_n),
    .write4_read(tdf7_l2_writeOutputs_149_U0_write4_read),
    .l2_partial_sums_address0(tdf7_l2_writeOutputs_149_U0_l2_partial_sums_address0),
    .l2_partial_sums_ce0(tdf7_l2_writeOutputs_149_U0_l2_partial_sums_ce0),
    .l2_partial_sums_q0(l2_products_t_q0),
    .out_data_address1(tdf7_l2_writeOutputs_149_U0_out_data_address1),
    .out_data_ce1(tdf7_l2_writeOutputs_149_U0_out_data_ce1),
    .out_data_we1(tdf7_l2_writeOutputs_149_U0_out_data_we1),
    .out_data_d1(tdf7_l2_writeOutputs_149_U0_out_data_d1),
    .l2_adjustments_address0(tdf7_l2_writeOutputs_149_U0_l2_adjustments_address0),
    .l2_adjustments_ce0(tdf7_l2_writeOutputs_149_U0_l2_adjustments_ce0),
    .l2_adjustments_q0(l2_adjustments_q0)
);

td_fused_top_fifo_w16_d2_S_x4 indices_01_c_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(indices_01_c_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf7_readInputs53_U0_indices_01_read),
    .if_dout(indices_01_c_dout),
    .if_full_n(indices_01_c_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf7_get_next_ijk_U0_indices_0_write),
    .if_din(tdf7_get_next_ijk_U0_indices_0_din)
);

td_fused_top_fifo_w16_d2_S_x4 indices_12_c_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(indices_12_c_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf7_readInputs53_U0_indices_12_read),
    .if_dout(indices_12_c_dout),
    .if_full_n(indices_12_c_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf7_get_next_ijk_U0_indices_1_write),
    .if_din(tdf7_get_next_ijk_U0_indices_1_din)
);

td_fused_top_fifo_w8_d2_S indices_23_c_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(indices_23_c_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf7_readFilters52_U0_indices_23_read),
    .if_dout(indices_23_c_dout),
    .if_full_n(indices_23_c_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf7_get_next_ijk_U0_indices_2_out_write),
    .if_din(tdf7_get_next_ijk_U0_indices_2_out_din)
);

td_fused_top_fifo_w13_d7_S indices_23_c1_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(indices_23_c1_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf7_adjust_U0_indices_23_read),
    .if_dout(indices_23_c1_dout),
    .if_full_n(indices_23_c1_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf7_get_next_ijk_U0_indices_2_out1_write),
    .if_din(tdf7_get_next_ijk_U0_indices_2_out1_din)
);

td_fused_top_fifo_w1_d9_S_x0 write4_c_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(write4_c_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf7_l2_writeOutputs_149_U0_write4_read),
    .if_dout(write4_c_dout),
    .if_full_n(write4_c_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf7_get_next_ijk_U0_write_r_write),
    .if_din(write4_c_din)
);

td_fused_top_fifo_w5_d8_S_x indices_01_c2_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(indices_01_c2_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf7_l2_writeOutputs_149_U0_indices_01_read),
    .if_dout(indices_01_c2_dout),
    .if_full_n(indices_01_c2_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf7_readInputs53_U0_indices_01_out_write),
    .if_din(tdf7_readInputs53_U0_indices_01_out_din)
);

td_fused_top_fifo_w10_d8_S_x indices_12_c3_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(indices_12_c3_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf7_l2_writeOutputs_149_U0_indices_12_read),
    .if_dout(indices_12_c3_dout),
    .if_full_n(indices_12_c3_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf7_readInputs53_U0_indices_12_out_write),
    .if_din(tdf7_readInputs53_U0_indices_12_out_din)
);

td_fused_top_fifo_w16_d2_S_x4 tmp_channel_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(tmp_channel_empty_n),
    .if_read_ce(1'b1),
    .if_read(Block_entry_proc_proc419_U0_ap_ready),
    .if_dout(tmp_channel_dout),
    .if_full_n(tmp_channel_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf7_accum_2_U0_ap_done),
    .if_din(tdf7_accum_2_U0_accum_in_6)
);

td_fused_top_fifo_w16_d2_S_x4 sums_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(sums_0_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf7_adjust_U0_ap_ready),
    .if_dout(sums_0_dout),
    .if_full_n(sums_0_full_n),
    .if_write_ce(1'b1),
    .if_write(Block_entry_proc_proc419_U0_ap_done),
    .if_din(Block_entry_proc_proc419_U0_ap_return)
);

td_fused_top_fifo_w13_d2_S indices_23_c4_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(indices_23_c4_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf7_l2_multiply50_U0_indices_23_read),
    .if_dout(indices_23_c4_dout),
    .if_full_n(indices_23_c4_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf7_adjust_U0_indices_23_out_write),
    .if_din(tdf7_adjust_U0_indices_23_out_din)
);

td_fused_top_fifo_w16_d2_S_x4 intermediate_fmaps_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(intermediate_fmaps_0_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf7_l2_multiply50_U0_ap_ready),
    .if_dout(intermediate_fmaps_0_dout),
    .if_full_n(intermediate_fmaps_0_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf7_adjust_U0_ap_done),
    .if_din(tdf7_adjust_U0_ap_return)
);

td_fused_top_start_for_tdf7_readFilters52_U0 start_for_tdf7_readFilters52_U0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(start_for_tdf7_readFilters52_U0_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf7_readFilters52_U0_ap_ready),
    .if_dout(start_for_tdf7_readFilters52_U0_dout),
    .if_full_n(start_for_tdf7_readFilters52_U0_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf7_get_next_ijk_U0_start_write),
    .if_din(start_for_tdf7_readFilters52_U0_din)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_sync_reg_tdf7_get_next_ijk_U0_ap_ready <= 1'b0;
    end else begin
        if (((ap_sync_ready & ap_start) == 1'b1)) begin
            ap_sync_reg_tdf7_get_next_ijk_U0_ap_ready <= 1'b0;
        end else begin
            ap_sync_reg_tdf7_get_next_ijk_U0_ap_ready <= ap_sync_tdf7_get_next_ijk_U0_ap_ready;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_sync_reg_tdf7_readInputs53_U0_ap_ready <= 1'b0;
    end else begin
        if (((ap_sync_ready & ap_start) == 1'b1)) begin
            ap_sync_reg_tdf7_readInputs53_U0_ap_ready <= 1'b0;
        end else begin
            ap_sync_reg_tdf7_readInputs53_U0_ap_ready <= ap_sync_tdf7_readInputs53_U0_ap_ready;
        end
    end
end

assign Block_entry_proc_proc419_U0_ap_continue = sums_0_full_n;

assign Block_entry_proc_proc419_U0_ap_start = tmp_channel_empty_n;

assign Block_entry_proc_proc419_U0_start_full_n = 1'b1;

assign Block_entry_proc_proc419_U0_start_write = 1'b0;

assign ap_channel_done_accum1_out_0 = tdf7_accum_1_U0_ap_done;

assign ap_channel_done_ifmap_vec = tdf7_readInputs53_U0_ap_done;

assign ap_channel_done_intermediate_fmaps_0 = tdf7_adjust_U0_ap_done;

assign ap_channel_done_l2_products = tdf7_l2_multiply50_U0_ap_done;

assign ap_channel_done_products_0 = tdf7_dot_product_U0_ap_done;

assign ap_channel_done_sums_0 = Block_entry_proc_proc419_U0_ap_done;

assign ap_channel_done_tmp_channel = tdf7_accum_2_U0_ap_done;

assign ap_channel_done_weight_vecs_0 = tdf7_readFilters52_U0_ap_done;

assign ap_done = tdf7_l2_writeOutputs_149_U0_ap_done;

assign ap_idle = (tdf7_readInputs53_U0_ap_idle & tdf7_readFilters52_U0_ap_idle & tdf7_l2_writeOutputs_149_U0_ap_idle & tdf7_l2_multiply50_U0_ap_idle & tdf7_get_next_ijk_U0_ap_idle & tdf7_dot_product_U0_ap_idle & tdf7_adjust_U0_ap_idle & tdf7_accum_2_U0_ap_idle & tdf7_accum_1_U0_ap_idle & (intermediate_fmaps_0_empty_n ^ 1'b1) & (sums_0_empty_n ^ 1'b1) & (tmp_channel_empty_n ^ 1'b1) & (l2_products_t_empty_n ^ 1'b1) & (products_0_t_empty_n ^ 1'b1) & (weight_vecs_0_t_empty_n ^ 1'b1) & (ifmap_vec_t_empty_n ^ 1'b1) & (1'b1 ^ accum1_out_0_t_empty_n) & Block_entry_proc_proc419_U0_ap_idle);

assign ap_ready = ap_sync_ready;

assign ap_sync_continue = ap_continue;

assign ap_sync_done = tdf7_l2_writeOutputs_149_U0_ap_done;

assign ap_sync_ready = (ap_sync_tdf7_readInputs53_U0_ap_ready & ap_sync_tdf7_get_next_ijk_U0_ap_ready);

assign ap_sync_tdf7_get_next_ijk_U0_ap_ready = (tdf7_get_next_ijk_U0_ap_ready | ap_sync_reg_tdf7_get_next_ijk_U0_ap_ready);

assign ap_sync_tdf7_readInputs53_U0_ap_ready = (tdf7_readInputs53_U0_ap_ready | ap_sync_reg_tdf7_readInputs53_U0_ap_ready);

assign in_data_address0 = tdf7_readInputs53_U0_in_data_address0;

assign in_data_address1 = 13'd0;

assign in_data_ce0 = tdf7_readInputs53_U0_in_data_ce0;

assign in_data_ce1 = 1'b0;

assign in_data_d0 = 64'd0;

assign in_data_d1 = 64'd0;

assign in_data_read = tdf7_readInputs53_U0_in_data_write;

assign in_data_we0 = 1'b0;

assign in_data_we1 = 1'b0;

assign l1_adjustments_address0 = tdf7_adjust_U0_adjustments_address0;

assign l1_adjustments_address1 = 8'd0;

assign l1_adjustments_ce0 = tdf7_adjust_U0_adjustments_ce0;

assign l1_adjustments_ce1 = 1'b0;

assign l1_adjustments_d0 = 48'd0;

assign l1_adjustments_d1 = 48'd0;

assign l1_adjustments_we0 = 1'b0;

assign l1_adjustments_we1 = 1'b0;

assign l1_filter_data_address0 = tdf7_readFilters52_U0_filter_data_address0;

assign l1_filter_data_address1 = 17'd0;

assign l1_filter_data_ce0 = tdf7_readFilters52_U0_filter_data_ce0;

assign l1_filter_data_ce1 = 1'b0;

assign l1_filter_data_d0 = 16'd0;

assign l1_filter_data_d1 = 16'd0;

assign l1_filter_data_we0 = 1'b0;

assign l1_filter_data_we1 = 1'b0;

assign l2_adjustments_address0 = tdf7_l2_writeOutputs_149_U0_l2_adjustments_address0;

assign l2_adjustments_address1 = 5'd0;

assign l2_adjustments_ce0 = tdf7_l2_writeOutputs_149_U0_l2_adjustments_ce0;

assign l2_adjustments_ce1 = 1'b0;

assign l2_adjustments_d0 = 48'd0;

assign l2_adjustments_d1 = 48'd0;

assign l2_adjustments_we0 = 1'b0;

assign l2_adjustments_we1 = 1'b0;

assign l2_filter_data_address0 = tdf7_l2_multiply50_U0_l2_filter_data_address0;

assign l2_filter_data_address1 = 13'd0;

assign l2_filter_data_ce0 = tdf7_l2_multiply50_U0_l2_filter_data_ce0;

assign l2_filter_data_ce1 = 1'b0;

assign l2_filter_data_d0 = 16'd0;

assign l2_filter_data_d1 = 16'd0;

assign l2_filter_data_we0 = 1'b0;

assign l2_filter_data_we1 = 1'b0;

assign out_data_address0 = 13'd0;

assign out_data_address1 = tdf7_l2_writeOutputs_149_U0_out_data_address1;

assign out_data_ce0 = 1'b0;

assign out_data_ce1 = tdf7_l2_writeOutputs_149_U0_out_data_ce1;

assign out_data_d0 = 64'd0;

assign out_data_d1 = tdf7_l2_writeOutputs_149_U0_out_data_d1;

assign out_data_we0 = 1'b0;

assign out_data_we1 = tdf7_l2_writeOutputs_149_U0_out_data_we1;

assign out_data_write = tdf7_l2_writeOutputs_149_U0_out_data_write;

assign products_0_t_d1 = 16'd0;

assign products_0_t_we1 = 1'b0;

assign start_for_tdf7_readFilters52_U0_din = 1'b1;

assign tdf7_accum_1_U0_accum_out_full_n = accum1_out_0_i_full_n;

assign tdf7_accum_1_U0_ap_continue = accum1_out_0_i_full_n;

assign tdf7_accum_1_U0_ap_start = products_0_t_empty_n;

assign tdf7_accum_1_U0_start_full_n = 1'b1;

assign tdf7_accum_1_U0_start_write = 1'b0;

assign tdf7_accum_2_U0_ap_continue = tmp_channel_full_n;

assign tdf7_accum_2_U0_ap_start = accum1_out_0_t_empty_n;

assign tdf7_accum_2_U0_start_full_n = 1'b1;

assign tdf7_accum_2_U0_start_write = 1'b0;

assign tdf7_adjust_U0_ap_continue = intermediate_fmaps_0_full_n;

assign tdf7_adjust_U0_ap_start = sums_0_empty_n;

assign tdf7_adjust_U0_start_full_n = 1'b1;

assign tdf7_adjust_U0_start_write = 1'b0;

assign tdf7_dot_product_U0_ap_continue = products_0_i_full_n;

assign tdf7_dot_product_U0_ap_start = (weight_vecs_0_t_empty_n & ifmap_vec_t_empty_n);

assign tdf7_dot_product_U0_products_0_full_n = products_0_i_full_n;

assign tdf7_dot_product_U0_start_full_n = 1'b1;

assign tdf7_dot_product_U0_start_write = 1'b0;

assign tdf7_get_next_ijk_U0_ap_continue = 1'b1;

assign tdf7_get_next_ijk_U0_ap_start = ((ap_sync_reg_tdf7_get_next_ijk_U0_ap_ready ^ 1'b1) & ap_start);

assign tdf7_l2_multiply50_U0_ap_continue = l2_products_i_full_n;

assign tdf7_l2_multiply50_U0_ap_start = intermediate_fmaps_0_empty_n;

assign tdf7_l2_multiply50_U0_l2_products_full_n = l2_products_i_full_n;

assign tdf7_l2_multiply50_U0_start_full_n = 1'b1;

assign tdf7_l2_multiply50_U0_start_write = 1'b0;

assign tdf7_l2_writeOutputs_149_U0_ap_continue = ap_continue;

assign tdf7_l2_writeOutputs_149_U0_ap_start = l2_products_t_empty_n;

assign tdf7_l2_writeOutputs_149_U0_out_data_full_n = out_data_full_n;

assign tdf7_l2_writeOutputs_149_U0_out_data_write = 1'b0;

assign tdf7_l2_writeOutputs_149_U0_start_full_n = 1'b1;

assign tdf7_l2_writeOutputs_149_U0_start_write = 1'b0;

assign tdf7_readFilters52_U0_ap_continue = weight_vecs_0_i_full_n;

assign tdf7_readFilters52_U0_ap_start = start_for_tdf7_readFilters52_U0_empty_n;

assign tdf7_readFilters52_U0_start_full_n = 1'b1;

assign tdf7_readFilters52_U0_start_write = 1'b0;

assign tdf7_readFilters52_U0_weight_vecs_0_full_n = weight_vecs_0_i_full_n;

assign tdf7_readInputs53_U0_ap_continue = ifmap_vec_i_full_n;

assign tdf7_readInputs53_U0_ap_start = ((ap_sync_reg_tdf7_readInputs53_U0_ap_ready ^ 1'b1) & ap_start);

assign tdf7_readInputs53_U0_ifmap_vec_full_n = ifmap_vec_i_full_n;

assign tdf7_readInputs53_U0_in_data_full_n = in_data_empty_n;

assign tdf7_readInputs53_U0_in_data_write = 1'b0;

assign tdf7_readInputs53_U0_start_full_n = 1'b1;

assign tdf7_readInputs53_U0_start_write = 1'b0;

assign write4_c_din = tdf7_get_next_ijk_U0_write_r_din;

endmodule //td_fused_top_dataflow_in_loop_TOP_LOOP37548
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37548_weight_vecs_0_memcore_ram (addr0, ce0, d0, we0, q0, addr1, ce1, d1, we1, q1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 10;
parameter MEM_SIZE = 576;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
output reg[DWIDTH-1:0] q1;
input clk;

reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];




always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1) 
            ram[addr1] <= d1; 
        q1 <= ram[addr1];
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37548_weight_vecs_0_memcore(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    q0,
    address1,
    ce1,
    we1,
    d1,
    q1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd576;
parameter AddressWidth = 32'd10;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;
output[DataWidth - 1:0] q1;



td_fused_top_dataflow_in_loop_TOP_LOOP37548_weight_vecs_0_memcore_ram td_fused_top_dataflow_in_loop_TOP_LOOP37548_weight_vecs_0_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 ),
    .q1( q1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_dataflow_in_loop_TOP_LOOP37548_weight_vecs_0
#(parameter
    DataWidth    = 16,
    AddressRange = 32,
    AddressWidth = 9,
    BufferCount  = 2,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire                    i_we0,
    input  wire [AddressWidth-1:0] i_address0,
    input  wire [DataWidth-1:0]    i_d0,
    output wire [DataWidth-1:0]    i_q0,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire                    t_we0,
    input  wire [AddressWidth-1:0] t_address0,
    input  wire [DataWidth-1:0]    t_d0,
    output wire [DataWidth-1:0]    t_q0
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
wire [AddressWidth+IndexWidth-1:0]   memcore_iaddr;
wire [AddressWidth+IndexWidth-1:0]   memcore_taddr;

//------------------------Instantiation------------------
assign memcore_iaddr = {i_address0, iptr};
assign memcore_taddr = {t_address0, tptr};
td_fused_top_dataflow_in_loop_TOP_LOOP37548_weight_vecs_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP37548_weight_vecs_0_memcore_U (
    .reset    ( reset ),
    .clk      ( clk ),
    .address0 ( memcore_iaddr ),
    .ce0      ( i_ce0 ),
    .we0      ( i_we0),
    .d0       ( i_d0 ),
    .q0       ( i_q0 ),
    .address1 ( memcore_taddr ),
    .ce1      ( t_ce0 ),
    .we1      ( t_we0),
    .d1       ( t_d0 ),
    .q1       ( t_q0 )

);

//------------------------Body---------------------------

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37644_accum1_out_0_memcore_ram (addr0, ce0, d0, we0, q0, addr1, ce1, d1, we1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 3;
parameter MEM_SIZE = 8;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
input clk;

reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];




always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1) 
            ram[addr1] <= d1; 
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37644_accum1_out_0_memcore(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    q0,
    address1,
    ce1,
    we1,
    d1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd8;
parameter AddressWidth = 32'd3;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;



td_fused_top_dataflow_in_loop_TOP_LOOP37644_accum1_out_0_memcore_ram td_fused_top_dataflow_in_loop_TOP_LOOP37644_accum1_out_0_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_dataflow_in_loop_TOP_LOOP37644_accum1_out_0
#(parameter
    DataWidth    = 16,
    AddressRange = 32,
    AddressWidth = 3,
    BufferCount  = 2,
    MemLatency   = 1,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire                    i_we0,
    input  wire [AddressWidth-1:0] i_address0,
    input  wire [DataWidth-1:0]    i_d0,
    output wire [DataWidth-1:0]    i_q0,
    input  wire                    i_ce1,
    input  wire                    i_we1,
    input  wire [AddressWidth-1:0] i_address1,
    input  wire [DataWidth-1:0]    i_d1,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire                    t_we0,
    input  wire [AddressWidth-1:0] t_address0,
    input  wire [DataWidth-1:0]    t_d0,
    output wire [DataWidth-1:0]    t_q0,
    input  wire                    t_ce1,
    input  wire                    t_we1,
    input  wire [AddressWidth-1:0] t_address1,
    input  wire [DataWidth-1:0]    t_d1
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth-1:0]   prev_iptr    = 1'b0; // previous initiator index
reg  [IndexWidth-1:0]   prev_tptr    = 1'b0; // previous target index
reg  [DataWidth-1:0]    reg_q0      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid0    = 1'b0; // buffer has valid data
reg  [DataWidth-1:0]    reg_q1      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid1    = 1'b0; // buffer has valid data
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
// buffer signals
wire [BufferCount-1:0] buf_ce0;
wire [BufferCount-1:0] buf_we0;
wire [AddressWidth-1:0] buf_a0_0, buf_a0_1;
wire [DataWidth-1:0] buf_d0_0, buf_d0_1;
wire [DataWidth-1:0] buf_q0_0, buf_q0_1;
wire [BufferCount-1:0] buf_ce1;
wire [BufferCount-1:0] buf_we1;
wire [AddressWidth-1:0] buf_a1_0, buf_a1_1;
wire [DataWidth-1:0] buf_d1_0, buf_d1_1;
//------------------------Instantiation------------------
//genvar i;
        td_fused_top_dataflow_in_loop_TOP_LOOP37644_accum1_out_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP37644_accum1_out_0_memcore_U_0 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_0 ),
            .ce0      ( buf_ce0[ 0 ] ),
            .we0      ( buf_we0[ 0 ] ),
            .d0       ( buf_d0_0 ),
            .q0       ( buf_q0_0 ),
            .address1 ( buf_a1_0 ),
            .ce1      ( buf_ce1[ 0 ] ),
            .we1      ( buf_we1[ 0 ] ),
            .d1       ( buf_d1_0 )
        );
        td_fused_top_dataflow_in_loop_TOP_LOOP37644_accum1_out_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP37644_accum1_out_0_memcore_U_1 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_1 ),
            .ce0      ( buf_ce0[ 1 ] ),
            .we0      ( buf_we0[ 1 ] ),
            .d0       ( buf_d0_1 ),
            .q0       ( buf_q0_1 ),
            .address1 ( buf_a1_1 ),
            .ce1      ( buf_ce1[ 1 ] ),
            .we1      ( buf_we1[ 1 ] ),
            .d1       ( buf_d1_1 )
        );

//++++++++++++++++++++++++buffer signals+++++++++++++++++
        assign buf_ce0[ 0 ] = (tptr ==  0  && empty_n) ? t_ce0
                             : (iptr ==  0 ) ? i_ce0 : 1'b0;
        assign buf_a0_0  = (tptr ==  0  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 0 ] = (tptr ==  0  && empty_n)  ? t_we0
                             : (iptr ==  0 ) ? i_we0 : 1'b0;
        assign buf_d0_0  = (tptr ==  0  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 0 ] = (tptr ==  0  && empty_n) ? t_ce1
                             : (iptr ==  0 ) ? i_ce1 : 1'b0;
        assign buf_a1_0  = (tptr ==  0  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 0 ] = (tptr ==  0  && empty_n)  ? t_we1
                             : (iptr ==  0 ) ? i_we1 : 1'b0;
        assign buf_d1_0  = (tptr ==  0  && empty_n) ? t_d1       : i_d1;
        assign buf_ce0[ 1 ] = (tptr ==  1  && empty_n) ? t_ce0
                             : (iptr ==  1 ) ? i_ce0 : 1'b0;
        assign buf_a0_1  = (tptr ==  1  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 1 ] = (tptr ==  1  && empty_n)  ? t_we0
                             : (iptr ==  1 ) ? i_we0 : 1'b0;
        assign buf_d0_1  = (tptr ==  1  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 1 ] = (tptr ==  1  && empty_n) ? t_ce1
                             : (iptr ==  1 ) ? i_ce1 : 1'b0;
        assign buf_a1_1  = (tptr ==  1  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 1 ] = (tptr ==  1  && empty_n)  ? t_we1
                             : (iptr ==  1 ) ? i_we1 : 1'b0;
        assign buf_d1_1  = (tptr ==  1  && empty_n) ? t_d1       : i_d1;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//------------------------Body---------------------------
assign i_q0      = (prev_iptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign t_q0      = reg_valid0 ? reg_q0 : (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// prev_iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_iptr <= 1'b0;
    else begin
        prev_iptr <= iptr;
    end
end

// prev_tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_tptr <= 1'b0;
    else begin
        prev_tptr <= tptr;
    end
end

// reg_q0 and reg_valid0
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q0     <= 1'b0;
        reg_valid0 <= 1'b0;
    end else if (!t_ce0 && !reg_valid0) begin
        reg_q0     <= (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
        reg_valid0 <= 1'b1;
    end else if (t_ce0) begin
        reg_valid0 <= 1'b0;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37644_ifmap_vec_0_0_memcore_ram (addr0, ce0, d0, we0, q0, addr1, ce1, d1, we1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
input clk;

reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];




always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1) 
            ram[addr1] <= d1; 
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37644_ifmap_vec_0_0_memcore(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    q0,
    address1,
    ce1,
    we1,
    d1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;



td_fused_top_dataflow_in_loop_TOP_LOOP37644_ifmap_vec_0_0_memcore_ram td_fused_top_dataflow_in_loop_TOP_LOOP37644_ifmap_vec_0_0_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_dataflow_in_loop_TOP_LOOP37644_ifmap_vec_0_0
#(parameter
    DataWidth    = 16,
    AddressRange = 32,
    AddressWidth = 7,
    BufferCount  = 2,
    MemLatency   = 1,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire                    i_we0,
    input  wire [AddressWidth-1:0] i_address0,
    input  wire [DataWidth-1:0]    i_d0,
    output wire [DataWidth-1:0]    i_q0,
    input  wire                    i_ce1,
    input  wire                    i_we1,
    input  wire [AddressWidth-1:0] i_address1,
    input  wire [DataWidth-1:0]    i_d1,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire                    t_we0,
    input  wire [AddressWidth-1:0] t_address0,
    input  wire [DataWidth-1:0]    t_d0,
    output wire [DataWidth-1:0]    t_q0,
    input  wire                    t_ce1,
    input  wire                    t_we1,
    input  wire [AddressWidth-1:0] t_address1,
    input  wire [DataWidth-1:0]    t_d1
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth-1:0]   prev_iptr    = 1'b0; // previous initiator index
reg  [IndexWidth-1:0]   prev_tptr    = 1'b0; // previous target index
reg  [DataWidth-1:0]    reg_q0      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid0    = 1'b0; // buffer has valid data
reg  [DataWidth-1:0]    reg_q1      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid1    = 1'b0; // buffer has valid data
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
// buffer signals
wire [BufferCount-1:0] buf_ce0;
wire [BufferCount-1:0] buf_we0;
wire [AddressWidth-1:0] buf_a0_0, buf_a0_1;
wire [DataWidth-1:0] buf_d0_0, buf_d0_1;
wire [DataWidth-1:0] buf_q0_0, buf_q0_1;
wire [BufferCount-1:0] buf_ce1;
wire [BufferCount-1:0] buf_we1;
wire [AddressWidth-1:0] buf_a1_0, buf_a1_1;
wire [DataWidth-1:0] buf_d1_0, buf_d1_1;
//------------------------Instantiation------------------
//genvar i;
        td_fused_top_dataflow_in_loop_TOP_LOOP37644_ifmap_vec_0_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP37644_ifmap_vec_0_0_memcore_U_0 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_0 ),
            .ce0      ( buf_ce0[ 0 ] ),
            .we0      ( buf_we0[ 0 ] ),
            .d0       ( buf_d0_0 ),
            .q0       ( buf_q0_0 ),
            .address1 ( buf_a1_0 ),
            .ce1      ( buf_ce1[ 0 ] ),
            .we1      ( buf_we1[ 0 ] ),
            .d1       ( buf_d1_0 )
        );
        td_fused_top_dataflow_in_loop_TOP_LOOP37644_ifmap_vec_0_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP37644_ifmap_vec_0_0_memcore_U_1 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_1 ),
            .ce0      ( buf_ce0[ 1 ] ),
            .we0      ( buf_we0[ 1 ] ),
            .d0       ( buf_d0_1 ),
            .q0       ( buf_q0_1 ),
            .address1 ( buf_a1_1 ),
            .ce1      ( buf_ce1[ 1 ] ),
            .we1      ( buf_we1[ 1 ] ),
            .d1       ( buf_d1_1 )
        );

//++++++++++++++++++++++++buffer signals+++++++++++++++++
        assign buf_ce0[ 0 ] = (tptr ==  0  && empty_n) ? t_ce0
                             : (iptr ==  0 ) ? i_ce0 : 1'b0;
        assign buf_a0_0  = (tptr ==  0  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 0 ] = (tptr ==  0  && empty_n)  ? t_we0
                             : (iptr ==  0 ) ? i_we0 : 1'b0;
        assign buf_d0_0  = (tptr ==  0  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 0 ] = (tptr ==  0  && empty_n) ? t_ce1
                             : (iptr ==  0 ) ? i_ce1 : 1'b0;
        assign buf_a1_0  = (tptr ==  0  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 0 ] = (tptr ==  0  && empty_n)  ? t_we1
                             : (iptr ==  0 ) ? i_we1 : 1'b0;
        assign buf_d1_0  = (tptr ==  0  && empty_n) ? t_d1       : i_d1;
        assign buf_ce0[ 1 ] = (tptr ==  1  && empty_n) ? t_ce0
                             : (iptr ==  1 ) ? i_ce0 : 1'b0;
        assign buf_a0_1  = (tptr ==  1  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 1 ] = (tptr ==  1  && empty_n)  ? t_we0
                             : (iptr ==  1 ) ? i_we0 : 1'b0;
        assign buf_d0_1  = (tptr ==  1  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 1 ] = (tptr ==  1  && empty_n) ? t_ce1
                             : (iptr ==  1 ) ? i_ce1 : 1'b0;
        assign buf_a1_1  = (tptr ==  1  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 1 ] = (tptr ==  1  && empty_n)  ? t_we1
                             : (iptr ==  1 ) ? i_we1 : 1'b0;
        assign buf_d1_1  = (tptr ==  1  && empty_n) ? t_d1       : i_d1;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//------------------------Body---------------------------
assign i_q0      = (prev_iptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign t_q0      = reg_valid0 ? reg_q0 : (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// prev_iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_iptr <= 1'b0;
    else begin
        prev_iptr <= iptr;
    end
end

// prev_tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_tptr <= 1'b0;
    else begin
        prev_tptr <= tptr;
    end
end

// reg_q0 and reg_valid0
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q0     <= 1'b0;
        reg_valid0 <= 1'b0;
    end else if (!t_ce0 && !reg_valid0) begin
        reg_q0     <= (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
        reg_valid0 <= 1'b1;
    end else if (t_ce0) begin
        reg_valid0 <= 1'b0;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37644_products_0_memcore_ram (addr0, ce0, d0, we0, q0, addr1, ce1, q1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
output reg[DWIDTH-1:0] q1;
input clk;

reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];




always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        q1 <= ram[addr1];
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37644_products_0_memcore(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    q0,
    address1,
    ce1,
    q1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
output[DataWidth - 1:0] q1;



td_fused_top_dataflow_in_loop_TOP_LOOP37644_products_0_memcore_ram td_fused_top_dataflow_in_loop_TOP_LOOP37644_products_0_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .q1( q1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_dataflow_in_loop_TOP_LOOP37644_products_0
#(parameter
    DataWidth    = 16,
    AddressRange = 32,
    AddressWidth = 7,
    BufferCount  = 2,
    MemLatency   = 1,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire                    i_we0,
    input  wire [AddressWidth-1:0] i_address0,
    input  wire [DataWidth-1:0]    i_d0,
    output wire [DataWidth-1:0]    i_q0,
    input  wire                    i_ce1,
    input  wire [AddressWidth-1:0] i_address1,
    output wire [DataWidth-1:0]    i_q1,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire                    t_we0,
    input  wire [AddressWidth-1:0] t_address0,
    input  wire [DataWidth-1:0]    t_d0,
    output wire [DataWidth-1:0]    t_q0,
    input  wire                    t_ce1,
    input  wire [AddressWidth-1:0] t_address1,
    output wire [DataWidth-1:0]    t_q1
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth-1:0]   prev_iptr    = 1'b0; // previous initiator index
reg  [IndexWidth-1:0]   prev_tptr    = 1'b0; // previous target index
reg  [DataWidth-1:0]    reg_q0      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid0    = 1'b0; // buffer has valid data
reg  [DataWidth-1:0]    reg_q1      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid1    = 1'b0; // buffer has valid data
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
// buffer signals
wire [BufferCount-1:0] buf_ce0;
wire [BufferCount-1:0] buf_we0;
wire [AddressWidth-1:0] buf_a0_0, buf_a0_1;
wire [DataWidth-1:0] buf_d0_0, buf_d0_1;
wire [DataWidth-1:0] buf_q0_0, buf_q0_1;
wire [BufferCount-1:0] buf_ce1;
wire [AddressWidth-1:0] buf_a1_0, buf_a1_1;
wire [DataWidth-1:0] buf_q1_0, buf_q1_1;
//------------------------Instantiation------------------
//genvar i;
        td_fused_top_dataflow_in_loop_TOP_LOOP37644_products_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP37644_products_0_memcore_U_0 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_0 ),
            .ce0      ( buf_ce0[ 0 ] ),
            .we0      ( buf_we0[ 0 ] ),
            .d0       ( buf_d0_0 ),
            .q0       ( buf_q0_0 ),
            .address1 ( buf_a1_0 ),
            .ce1      ( buf_ce1[ 0 ] ),
            .q1       ( buf_q1_0 )
        );
        td_fused_top_dataflow_in_loop_TOP_LOOP37644_products_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP37644_products_0_memcore_U_1 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_1 ),
            .ce0      ( buf_ce0[ 1 ] ),
            .we0      ( buf_we0[ 1 ] ),
            .d0       ( buf_d0_1 ),
            .q0       ( buf_q0_1 ),
            .address1 ( buf_a1_1 ),
            .ce1      ( buf_ce1[ 1 ] ),
            .q1       ( buf_q1_1 )
        );

//++++++++++++++++++++++++buffer signals+++++++++++++++++
        assign buf_ce0[ 0 ] = (tptr ==  0  && empty_n) ? t_ce0
                             : (iptr ==  0 ) ? i_ce0 : 1'b0;
        assign buf_a0_0  = (tptr ==  0  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 0 ] = (tptr ==  0  && empty_n)  ? t_we0
                             : (iptr ==  0 ) ? i_we0 : 1'b0;
        assign buf_d0_0  = (tptr ==  0  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 0 ] = (tptr ==  0  && empty_n) ? t_ce1
                             : (iptr ==  0 ) ? i_ce1 : 1'b0;
        assign buf_a1_0  = (tptr ==  0  && empty_n) ?  t_address1 : i_address1;
        assign buf_ce0[ 1 ] = (tptr ==  1  && empty_n) ? t_ce0
                             : (iptr ==  1 ) ? i_ce0 : 1'b0;
        assign buf_a0_1  = (tptr ==  1  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 1 ] = (tptr ==  1  && empty_n)  ? t_we0
                             : (iptr ==  1 ) ? i_we0 : 1'b0;
        assign buf_d0_1  = (tptr ==  1  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 1 ] = (tptr ==  1  && empty_n) ? t_ce1
                             : (iptr ==  1 ) ? i_ce1 : 1'b0;
        assign buf_a1_1  = (tptr ==  1  && empty_n) ?  t_address1 : i_address1;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//------------------------Body---------------------------
assign i_q0      = (prev_iptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign t_q0      = reg_valid0 ? reg_q0 : (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign i_q1      = (prev_iptr == 1'b1 ? buf_q1_1 : buf_q1_0);
assign t_q1      = reg_valid1 ? reg_q1 : (prev_tptr == 1'b1 ? buf_q1_1 : buf_q1_0);

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// prev_iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_iptr <= 1'b0;
    else begin
        prev_iptr <= iptr;
    end
end

// prev_tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_tptr <= 1'b0;
    else begin
        prev_tptr <= tptr;
    end
end

// reg_q0 and reg_valid0
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q0     <= 1'b0;
        reg_valid0 <= 1'b0;
    end else if (!t_ce0 && !reg_valid0) begin
        reg_q0     <= (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
        reg_valid0 <= 1'b1;
    end else if (t_ce0) begin
        reg_valid0 <= 1'b0;
    end
end

// reg_q1 and reg_valid1
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q1     <= 1'b0;
        reg_valid1 <= 1'b0;
    end else if (!t_ce1 && !reg_valid1) begin
        reg_q1     <= (prev_tptr == 1'b1 ? buf_q1_1 : buf_q1_0);
        reg_valid1 <= 1'b1;
    end else if (t_ce1) begin
        reg_valid1 <= 1'b0;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_dataflow_in_loop_TOP_LOOP37644 (
        ap_clk,
        ap_rst,
        in_data_address0,
        in_data_ce0,
        in_data_d0,
        in_data_q0,
        in_data_we0,
        in_data_address1,
        in_data_ce1,
        in_data_d1,
        in_data_q1,
        in_data_we1,
        filter_data_address0,
        filter_data_ce0,
        filter_data_d0,
        filter_data_q0,
        filter_data_we0,
        filter_data_address1,
        filter_data_ce1,
        filter_data_d1,
        filter_data_q1,
        filter_data_we1,
        adjustments_address0,
        adjustments_ce0,
        adjustments_d0,
        adjustments_q0,
        adjustments_we0,
        adjustments_address1,
        adjustments_ce1,
        adjustments_d1,
        adjustments_q1,
        adjustments_we1,
        out_data_address0,
        out_data_ce0,
        out_data_d0,
        out_data_q0,
        out_data_we0,
        out_data_address1,
        out_data_ce1,
        out_data_d1,
        out_data_q1,
        out_data_we1,
        ap_start,
        in_data_empty_n,
        in_data_read,
        out_data_full_n,
        out_data_write,
        ap_done,
        ap_ready,
        ap_idle,
        ap_continue
);


input   ap_clk;
input   ap_rst;
output  [14:0] in_data_address0;
output   in_data_ce0;
output  [63:0] in_data_d0;
input  [63:0] in_data_q0;
output   in_data_we0;
output  [14:0] in_data_address1;
output   in_data_ce1;
output  [63:0] in_data_d1;
input  [63:0] in_data_q1;
output   in_data_we1;
output  [11:0] filter_data_address0;
output   filter_data_ce0;
output  [15:0] filter_data_d0;
input  [15:0] filter_data_q0;
output   filter_data_we0;
output  [11:0] filter_data_address1;
output   filter_data_ce1;
output  [15:0] filter_data_d1;
input  [15:0] filter_data_q1;
output   filter_data_we1;
output  [4:0] adjustments_address0;
output   adjustments_ce0;
output  [47:0] adjustments_d0;
input  [47:0] adjustments_q0;
output   adjustments_we0;
output  [4:0] adjustments_address1;
output   adjustments_ce1;
output  [47:0] adjustments_d1;
input  [47:0] adjustments_q1;
output   adjustments_we1;
output  [12:0] out_data_address0;
output   out_data_ce0;
output  [63:0] out_data_d0;
input  [63:0] out_data_q0;
output   out_data_we0;
output  [12:0] out_data_address1;
output   out_data_ce1;
output  [63:0] out_data_d1;
input  [63:0] out_data_q1;
output   out_data_we1;
input   ap_start;
input   in_data_empty_n;
output   in_data_read;
input   out_data_full_n;
output   out_data_write;
output   ap_done;
output   ap_ready;
output   ap_idle;
input   ap_continue;

wire   [15:0] ifmap_vec_0_0_i_q0;
wire   [15:0] ifmap_vec_0_0_t_q0;
wire   [15:0] weight_vecs_0_0_0_i_q0;
wire   [15:0] weight_vecs_0_0_0_t_q0;
wire   [15:0] products_0_i_q0;
wire   [15:0] products_0_i_q1;
wire   [15:0] products_0_t_q0;
wire   [15:0] products_0_t_q1;
wire   [15:0] accum1_out_0_i_q0;
wire   [15:0] accum1_out_0_t_q0;
wire    tdf6_get_next_ijk_U0_ap_start;
wire    tdf6_get_next_ijk_U0_ap_done;
wire    tdf6_get_next_ijk_U0_ap_continue;
wire    tdf6_get_next_ijk_U0_ap_idle;
wire    tdf6_get_next_ijk_U0_ap_ready;
wire    tdf6_get_next_ijk_U0_start_out;
wire    tdf6_get_next_ijk_U0_start_write;
wire   [15:0] tdf6_get_next_ijk_U0_indices_0_din;
wire    tdf6_get_next_ijk_U0_indices_0_write;
wire   [15:0] tdf6_get_next_ijk_U0_indices_1_din;
wire    tdf6_get_next_ijk_U0_indices_1_write;
wire   [4:0] tdf6_get_next_ijk_U0_indices_2_out_din;
wire    tdf6_get_next_ijk_U0_indices_2_out_write;
wire   [4:0] tdf6_get_next_ijk_U0_indices_2_out1_din;
wire    tdf6_get_next_ijk_U0_indices_2_out1_write;
wire    tdf6_readInputs_U0_ap_start;
wire    tdf6_readInputs_U0_ap_done;
wire    tdf6_readInputs_U0_ap_continue;
wire    tdf6_readInputs_U0_ap_idle;
wire    tdf6_readInputs_U0_ap_ready;
wire   [14:0] tdf6_readInputs_U0_in_data_address0;
wire    tdf6_readInputs_U0_in_data_ce0;
wire    tdf6_readInputs_U0_indices_01_read;
wire    tdf6_readInputs_U0_indices_12_read;
wire   [6:0] tdf6_readInputs_U0_ifmap_vec_0_0_address0;
wire    tdf6_readInputs_U0_ifmap_vec_0_0_ce0;
wire    tdf6_readInputs_U0_ifmap_vec_0_0_we0;
wire   [15:0] tdf6_readInputs_U0_ifmap_vec_0_0_d0;
wire   [6:0] tdf6_readInputs_U0_ifmap_vec_0_0_address1;
wire    tdf6_readInputs_U0_ifmap_vec_0_0_ce1;
wire    tdf6_readInputs_U0_ifmap_vec_0_0_we1;
wire   [15:0] tdf6_readInputs_U0_ifmap_vec_0_0_d1;
wire   [4:0] tdf6_readInputs_U0_indices_01_out_din;
wire    tdf6_readInputs_U0_indices_01_out_write;
wire   [9:0] tdf6_readInputs_U0_indices_12_out_din;
wire    tdf6_readInputs_U0_indices_12_out_write;
wire    tdf6_readInputs_U0_in_data_full_n;
wire    tdf6_readInputs_U0_in_data_write;
wire    ap_channel_done_ifmap_vec_0_0;
wire    tdf6_readInputs_U0_ifmap_vec_0_0_full_n;
wire    tdf6_readFilters46_U0_ap_start;
wire    tdf6_readFilters46_U0_ap_done;
wire    tdf6_readFilters46_U0_ap_continue;
wire    tdf6_readFilters46_U0_ap_idle;
wire    tdf6_readFilters46_U0_ap_ready;
wire   [11:0] tdf6_readFilters46_U0_filter_data_address0;
wire    tdf6_readFilters46_U0_filter_data_ce0;
wire    tdf6_readFilters46_U0_indices_23_read;
wire   [6:0] tdf6_readFilters46_U0_weight_vecs_0_0_0_address0;
wire    tdf6_readFilters46_U0_weight_vecs_0_0_0_ce0;
wire    tdf6_readFilters46_U0_weight_vecs_0_0_0_we0;
wire   [15:0] tdf6_readFilters46_U0_weight_vecs_0_0_0_d0;
wire    ap_channel_done_weight_vecs_0_0_0;
wire    tdf6_readFilters46_U0_weight_vecs_0_0_0_full_n;
wire    tdf6_dot_product_U0_ap_start;
wire    tdf6_dot_product_U0_ap_done;
wire    tdf6_dot_product_U0_ap_continue;
wire    tdf6_dot_product_U0_ap_idle;
wire    tdf6_dot_product_U0_ap_ready;
wire   [6:0] tdf6_dot_product_U0_ifmap_vec_0_0_address0;
wire    tdf6_dot_product_U0_ifmap_vec_0_0_ce0;
wire   [6:0] tdf6_dot_product_U0_weight_vecs_0_0_0_address0;
wire    tdf6_dot_product_U0_weight_vecs_0_0_0_ce0;
wire   [6:0] tdf6_dot_product_U0_products_0_address0;
wire    tdf6_dot_product_U0_products_0_ce0;
wire    tdf6_dot_product_U0_products_0_we0;
wire   [15:0] tdf6_dot_product_U0_products_0_d0;
wire    ap_channel_done_products_0;
wire    tdf6_dot_product_U0_products_0_full_n;
wire    tdf6_accum_1_U0_ap_start;
wire    tdf6_accum_1_U0_ap_done;
wire    tdf6_accum_1_U0_ap_continue;
wire    tdf6_accum_1_U0_ap_idle;
wire    tdf6_accum_1_U0_ap_ready;
wire   [6:0] tdf6_accum_1_U0_accum_in_0_address0;
wire    tdf6_accum_1_U0_accum_in_0_ce0;
wire   [6:0] tdf6_accum_1_U0_accum_in_0_address1;
wire    tdf6_accum_1_U0_accum_in_0_ce1;
wire   [2:0] tdf6_accum_1_U0_accum_out_address0;
wire    tdf6_accum_1_U0_accum_out_ce0;
wire    tdf6_accum_1_U0_accum_out_we0;
wire   [15:0] tdf6_accum_1_U0_accum_out_d0;
wire   [2:0] tdf6_accum_1_U0_accum_out_address1;
wire    tdf6_accum_1_U0_accum_out_ce1;
wire    tdf6_accum_1_U0_accum_out_we1;
wire   [15:0] tdf6_accum_1_U0_accum_out_d1;
wire    ap_channel_done_accum1_out_0;
wire    tdf6_accum_1_U0_accum_out_full_n;
wire    tdf6_accum_2_U0_ap_start;
wire    tdf6_accum_2_U0_ap_done;
wire    tdf6_accum_2_U0_ap_continue;
wire    tdf6_accum_2_U0_ap_idle;
wire    tdf6_accum_2_U0_ap_ready;
wire   [15:0] tdf6_accum_2_U0_accum_in_8;
wire    tdf6_accum_2_U0_accum_in_8_ap_vld;
wire   [2:0] tdf6_accum_2_U0_accum_in_address0;
wire    tdf6_accum_2_U0_accum_in_ce0;
wire    ap_channel_done_tmp_channel;
wire    tmp_channel_full_n;
wire    Block_entry_proc_proc413_U0_ap_start;
wire    Block_entry_proc_proc413_U0_ap_done;
wire    Block_entry_proc_proc413_U0_ap_continue;
wire    Block_entry_proc_proc413_U0_ap_idle;
wire    Block_entry_proc_proc413_U0_ap_ready;
wire   [15:0] Block_entry_proc_proc413_U0_ap_return;
wire    ap_channel_done_sums_0;
wire    sums_0_full_n;
wire    tdf6_adjust_U0_ap_start;
wire    tdf6_adjust_U0_ap_done;
wire    tdf6_adjust_U0_ap_continue;
wire    tdf6_adjust_U0_ap_idle;
wire    tdf6_adjust_U0_ap_ready;
wire   [4:0] tdf6_adjust_U0_adjustments_address0;
wire    tdf6_adjust_U0_adjustments_ce0;
wire    tdf6_adjust_U0_indices_23_read;
wire   [15:0] tdf6_adjust_U0_ap_return;
wire    ap_channel_done_outputs_0;
wire    outputs_0_full_n;
wire    tdf6_writeOutputs_unaligned_U0_ap_start;
wire    tdf6_writeOutputs_unaligned_U0_ap_done;
wire    tdf6_writeOutputs_unaligned_U0_ap_continue;
wire    tdf6_writeOutputs_unaligned_U0_ap_idle;
wire    tdf6_writeOutputs_unaligned_U0_ap_ready;
wire    tdf6_writeOutputs_unaligned_U0_indices_01_read;
wire    tdf6_writeOutputs_unaligned_U0_indices_12_read;
wire   [12:0] tdf6_writeOutputs_unaligned_U0_out_data_address1;
wire    tdf6_writeOutputs_unaligned_U0_out_data_ce1;
wire    tdf6_writeOutputs_unaligned_U0_out_data_we1;
wire   [63:0] tdf6_writeOutputs_unaligned_U0_out_data_d1;
wire    tdf6_writeOutputs_unaligned_U0_out_data_full_n;
wire    tdf6_writeOutputs_unaligned_U0_out_data_write;
wire    ap_sync_continue;
wire    ifmap_vec_0_0_i_full_n;
wire    ifmap_vec_0_0_t_empty_n;
wire    weight_vecs_0_0_0_i_full_n;
wire    weight_vecs_0_0_0_t_empty_n;
wire    products_0_i_full_n;
wire    products_0_t_empty_n;
wire   [15:0] products_0_t_d1;
wire    products_0_t_we1;
wire    accum1_out_0_i_full_n;
wire    accum1_out_0_t_empty_n;
wire    indices_01_c_full_n;
wire   [15:0] indices_01_c_dout;
wire    indices_01_c_empty_n;
wire    indices_12_c_full_n;
wire   [15:0] indices_12_c_dout;
wire    indices_12_c_empty_n;
wire    indices_23_c_full_n;
wire   [4:0] indices_23_c_dout;
wire    indices_23_c_empty_n;
wire    indices_23_c1_full_n;
wire   [4:0] indices_23_c1_dout;
wire    indices_23_c1_empty_n;
wire    indices_01_c2_full_n;
wire   [4:0] indices_01_c2_dout;
wire    indices_01_c2_empty_n;
wire    indices_12_c3_full_n;
wire   [9:0] indices_12_c3_dout;
wire    indices_12_c3_empty_n;
wire   [15:0] tmp_channel_dout;
wire    tmp_channel_empty_n;
wire   [15:0] sums_0_dout;
wire    sums_0_empty_n;
wire   [15:0] outputs_0_dout;
wire    outputs_0_empty_n;
wire    ap_sync_done;
wire    ap_sync_ready;
reg    ap_sync_reg_tdf6_get_next_ijk_U0_ap_ready;
wire    ap_sync_tdf6_get_next_ijk_U0_ap_ready;
reg    ap_sync_reg_tdf6_readInputs_U0_ap_ready;
wire    ap_sync_tdf6_readInputs_U0_ap_ready;
wire   [0:0] start_for_tdf6_readFilters46_U0_din;
wire    start_for_tdf6_readFilters46_U0_full_n;
wire   [0:0] start_for_tdf6_readFilters46_U0_dout;
wire    start_for_tdf6_readFilters46_U0_empty_n;
wire    tdf6_readInputs_U0_start_full_n;
wire    tdf6_readInputs_U0_start_write;
wire    tdf6_readFilters46_U0_start_full_n;
wire    tdf6_readFilters46_U0_start_write;
wire    tdf6_dot_product_U0_start_full_n;
wire    tdf6_dot_product_U0_start_write;
wire    tdf6_accum_1_U0_start_full_n;
wire    tdf6_accum_1_U0_start_write;
wire    tdf6_accum_2_U0_start_full_n;
wire    tdf6_accum_2_U0_start_write;
wire    Block_entry_proc_proc413_U0_start_full_n;
wire    Block_entry_proc_proc413_U0_start_write;
wire    tdf6_adjust_U0_start_full_n;
wire    tdf6_adjust_U0_start_write;
wire    tdf6_writeOutputs_unaligned_U0_start_full_n;
wire    tdf6_writeOutputs_unaligned_U0_start_write;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_sync_reg_tdf6_get_next_ijk_U0_ap_ready = 1'b0;
#0 ap_sync_reg_tdf6_readInputs_U0_ap_ready = 1'b0;
end

td_fused_top_dataflow_in_loop_TOP_LOOP37644_ifmap_vec_0_0 #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
ifmap_vec_0_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf6_readInputs_U0_ap_done),
    .i_full_n(ifmap_vec_0_0_i_full_n),
    .i_ce0(tdf6_readInputs_U0_ifmap_vec_0_0_ce0),
    .i_we0(tdf6_readInputs_U0_ifmap_vec_0_0_we0),
    .i_address0(tdf6_readInputs_U0_ifmap_vec_0_0_address0),
    .i_d0(tdf6_readInputs_U0_ifmap_vec_0_0_d0),
    .i_q0(ifmap_vec_0_0_i_q0),
    .i_ce1(tdf6_readInputs_U0_ifmap_vec_0_0_ce1),
    .i_we1(tdf6_readInputs_U0_ifmap_vec_0_0_we1),
    .i_address1(tdf6_readInputs_U0_ifmap_vec_0_0_address1),
    .i_d1(tdf6_readInputs_U0_ifmap_vec_0_0_d1),
    .t_ce(1'b1),
    .t_read(tdf6_dot_product_U0_ap_ready),
    .t_empty_n(ifmap_vec_0_0_t_empty_n),
    .t_ce0(tdf6_dot_product_U0_ifmap_vec_0_0_ce0),
    .t_we0(1'b0),
    .t_address0(tdf6_dot_product_U0_ifmap_vec_0_0_address0),
    .t_d0(16'd0),
    .t_q0(ifmap_vec_0_0_t_q0),
    .t_ce1(1'b0),
    .t_we1(1'b0),
    .t_address1(7'd0),
    .t_d1(16'd0)
);

td_fused_top_dataflow_in_loop_TOP_LOOP37644_weight_vecs_0_0_0 #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
weight_vecs_0_0_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf6_readFilters46_U0_ap_done),
    .i_full_n(weight_vecs_0_0_0_i_full_n),
    .i_ce0(tdf6_readFilters46_U0_weight_vecs_0_0_0_ce0),
    .i_we0(tdf6_readFilters46_U0_weight_vecs_0_0_0_we0),
    .i_address0(tdf6_readFilters46_U0_weight_vecs_0_0_0_address0),
    .i_d0(tdf6_readFilters46_U0_weight_vecs_0_0_0_d0),
    .i_q0(weight_vecs_0_0_0_i_q0),
    .t_ce(1'b1),
    .t_read(tdf6_dot_product_U0_ap_ready),
    .t_empty_n(weight_vecs_0_0_0_t_empty_n),
    .t_ce0(tdf6_dot_product_U0_weight_vecs_0_0_0_ce0),
    .t_we0(1'b0),
    .t_address0(tdf6_dot_product_U0_weight_vecs_0_0_0_address0),
    .t_d0(16'd0),
    .t_q0(weight_vecs_0_0_0_t_q0)
);

td_fused_top_dataflow_in_loop_TOP_LOOP37644_products_0 #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
products_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf6_dot_product_U0_ap_done),
    .i_full_n(products_0_i_full_n),
    .i_ce0(tdf6_dot_product_U0_products_0_ce0),
    .i_we0(tdf6_dot_product_U0_products_0_we0),
    .i_address0(tdf6_dot_product_U0_products_0_address0),
    .i_d0(tdf6_dot_product_U0_products_0_d0),
    .i_q0(products_0_i_q0),
    .i_ce1(1'b0),
    .i_address1(7'd0),
    .i_q1(products_0_i_q1),
    .t_ce(1'b1),
    .t_read(tdf6_accum_1_U0_ap_ready),
    .t_empty_n(products_0_t_empty_n),
    .t_ce0(tdf6_accum_1_U0_accum_in_0_ce0),
    .t_we0(1'b0),
    .t_address0(tdf6_accum_1_U0_accum_in_0_address0),
    .t_d0(16'd0),
    .t_q0(products_0_t_q0),
    .t_ce1(tdf6_accum_1_U0_accum_in_0_ce1),
    .t_address1(tdf6_accum_1_U0_accum_in_0_address1),
    .t_q1(products_0_t_q1)
);

td_fused_top_dataflow_in_loop_TOP_LOOP37644_accum1_out_0 #(
    .DataWidth( 16 ),
    .AddressRange( 8 ),
    .AddressWidth( 3 ))
accum1_out_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf6_accum_1_U0_ap_done),
    .i_full_n(accum1_out_0_i_full_n),
    .i_ce0(tdf6_accum_1_U0_accum_out_ce0),
    .i_we0(tdf6_accum_1_U0_accum_out_we0),
    .i_address0(tdf6_accum_1_U0_accum_out_address0),
    .i_d0(tdf6_accum_1_U0_accum_out_d0),
    .i_q0(accum1_out_0_i_q0),
    .i_ce1(tdf6_accum_1_U0_accum_out_ce1),
    .i_we1(tdf6_accum_1_U0_accum_out_we1),
    .i_address1(tdf6_accum_1_U0_accum_out_address1),
    .i_d1(tdf6_accum_1_U0_accum_out_d1),
    .t_ce(1'b1),
    .t_read(tdf6_accum_2_U0_ap_ready),
    .t_empty_n(accum1_out_0_t_empty_n),
    .t_ce0(tdf6_accum_2_U0_accum_in_ce0),
    .t_we0(1'b0),
    .t_address0(tdf6_accum_2_U0_accum_in_address0),
    .t_d0(16'd0),
    .t_q0(accum1_out_0_t_q0),
    .t_ce1(1'b0),
    .t_we1(1'b0),
    .t_address1(3'd0),
    .t_d1(16'd0)
);

td_fused_top_tdf6_get_next_ijk tdf6_get_next_ijk_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf6_get_next_ijk_U0_ap_start),
    .start_full_n(start_for_tdf6_readFilters46_U0_full_n),
    .ap_done(tdf6_get_next_ijk_U0_ap_done),
    .ap_continue(tdf6_get_next_ijk_U0_ap_continue),
    .ap_idle(tdf6_get_next_ijk_U0_ap_idle),
    .ap_ready(tdf6_get_next_ijk_U0_ap_ready),
    .start_out(tdf6_get_next_ijk_U0_start_out),
    .start_write(tdf6_get_next_ijk_U0_start_write),
    .indices_0_din(tdf6_get_next_ijk_U0_indices_0_din),
    .indices_0_full_n(indices_01_c_full_n),
    .indices_0_write(tdf6_get_next_ijk_U0_indices_0_write),
    .indices_1_din(tdf6_get_next_ijk_U0_indices_1_din),
    .indices_1_full_n(indices_12_c_full_n),
    .indices_1_write(tdf6_get_next_ijk_U0_indices_1_write),
    .indices_2_out_din(tdf6_get_next_ijk_U0_indices_2_out_din),
    .indices_2_out_full_n(indices_23_c_full_n),
    .indices_2_out_write(tdf6_get_next_ijk_U0_indices_2_out_write),
    .indices_2_out1_din(tdf6_get_next_ijk_U0_indices_2_out1_din),
    .indices_2_out1_full_n(indices_23_c1_full_n),
    .indices_2_out1_write(tdf6_get_next_ijk_U0_indices_2_out1_write)
);

td_fused_top_tdf6_readInputs tdf6_readInputs_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf6_readInputs_U0_ap_start),
    .ap_done(tdf6_readInputs_U0_ap_done),
    .ap_continue(tdf6_readInputs_U0_ap_continue),
    .ap_idle(tdf6_readInputs_U0_ap_idle),
    .ap_ready(tdf6_readInputs_U0_ap_ready),
    .in_data_address0(tdf6_readInputs_U0_in_data_address0),
    .in_data_ce0(tdf6_readInputs_U0_in_data_ce0),
    .in_data_q0(in_data_q0),
    .indices_01_dout(indices_01_c_dout),
    .indices_01_empty_n(indices_01_c_empty_n),
    .indices_01_read(tdf6_readInputs_U0_indices_01_read),
    .indices_12_dout(indices_12_c_dout),
    .indices_12_empty_n(indices_12_c_empty_n),
    .indices_12_read(tdf6_readInputs_U0_indices_12_read),
    .ifmap_vec_0_0_address0(tdf6_readInputs_U0_ifmap_vec_0_0_address0),
    .ifmap_vec_0_0_ce0(tdf6_readInputs_U0_ifmap_vec_0_0_ce0),
    .ifmap_vec_0_0_we0(tdf6_readInputs_U0_ifmap_vec_0_0_we0),
    .ifmap_vec_0_0_d0(tdf6_readInputs_U0_ifmap_vec_0_0_d0),
    .ifmap_vec_0_0_address1(tdf6_readInputs_U0_ifmap_vec_0_0_address1),
    .ifmap_vec_0_0_ce1(tdf6_readInputs_U0_ifmap_vec_0_0_ce1),
    .ifmap_vec_0_0_we1(tdf6_readInputs_U0_ifmap_vec_0_0_we1),
    .ifmap_vec_0_0_d1(tdf6_readInputs_U0_ifmap_vec_0_0_d1),
    .indices_01_out_din(tdf6_readInputs_U0_indices_01_out_din),
    .indices_01_out_full_n(indices_01_c2_full_n),
    .indices_01_out_write(tdf6_readInputs_U0_indices_01_out_write),
    .indices_12_out_din(tdf6_readInputs_U0_indices_12_out_din),
    .indices_12_out_full_n(indices_12_c3_full_n),
    .indices_12_out_write(tdf6_readInputs_U0_indices_12_out_write)
);

td_fused_top_tdf6_readFilters46 tdf6_readFilters46_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf6_readFilters46_U0_ap_start),
    .ap_done(tdf6_readFilters46_U0_ap_done),
    .ap_continue(tdf6_readFilters46_U0_ap_continue),
    .ap_idle(tdf6_readFilters46_U0_ap_idle),
    .ap_ready(tdf6_readFilters46_U0_ap_ready),
    .filter_data_address0(tdf6_readFilters46_U0_filter_data_address0),
    .filter_data_ce0(tdf6_readFilters46_U0_filter_data_ce0),
    .filter_data_q0(filter_data_q0),
    .indices_23_dout(indices_23_c_dout),
    .indices_23_empty_n(indices_23_c_empty_n),
    .indices_23_read(tdf6_readFilters46_U0_indices_23_read),
    .weight_vecs_0_0_0_address0(tdf6_readFilters46_U0_weight_vecs_0_0_0_address0),
    .weight_vecs_0_0_0_ce0(tdf6_readFilters46_U0_weight_vecs_0_0_0_ce0),
    .weight_vecs_0_0_0_we0(tdf6_readFilters46_U0_weight_vecs_0_0_0_we0),
    .weight_vecs_0_0_0_d0(tdf6_readFilters46_U0_weight_vecs_0_0_0_d0)
);

td_fused_top_tdf6_dot_product tdf6_dot_product_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf6_dot_product_U0_ap_start),
    .ap_done(tdf6_dot_product_U0_ap_done),
    .ap_continue(tdf6_dot_product_U0_ap_continue),
    .ap_idle(tdf6_dot_product_U0_ap_idle),
    .ap_ready(tdf6_dot_product_U0_ap_ready),
    .ifmap_vec_0_0_address0(tdf6_dot_product_U0_ifmap_vec_0_0_address0),
    .ifmap_vec_0_0_ce0(tdf6_dot_product_U0_ifmap_vec_0_0_ce0),
    .ifmap_vec_0_0_q0(ifmap_vec_0_0_t_q0),
    .weight_vecs_0_0_0_address0(tdf6_dot_product_U0_weight_vecs_0_0_0_address0),
    .weight_vecs_0_0_0_ce0(tdf6_dot_product_U0_weight_vecs_0_0_0_ce0),
    .weight_vecs_0_0_0_q0(weight_vecs_0_0_0_t_q0),
    .products_0_address0(tdf6_dot_product_U0_products_0_address0),
    .products_0_ce0(tdf6_dot_product_U0_products_0_ce0),
    .products_0_we0(tdf6_dot_product_U0_products_0_we0),
    .products_0_d0(tdf6_dot_product_U0_products_0_d0)
);

td_fused_top_tdf6_accum_1 tdf6_accum_1_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf6_accum_1_U0_ap_start),
    .ap_done(tdf6_accum_1_U0_ap_done),
    .ap_continue(tdf6_accum_1_U0_ap_continue),
    .ap_idle(tdf6_accum_1_U0_ap_idle),
    .ap_ready(tdf6_accum_1_U0_ap_ready),
    .accum_in_0_address0(tdf6_accum_1_U0_accum_in_0_address0),
    .accum_in_0_ce0(tdf6_accum_1_U0_accum_in_0_ce0),
    .accum_in_0_q0(products_0_t_q0),
    .accum_in_0_address1(tdf6_accum_1_U0_accum_in_0_address1),
    .accum_in_0_ce1(tdf6_accum_1_U0_accum_in_0_ce1),
    .accum_in_0_q1(products_0_t_q1),
    .accum_out_address0(tdf6_accum_1_U0_accum_out_address0),
    .accum_out_ce0(tdf6_accum_1_U0_accum_out_ce0),
    .accum_out_we0(tdf6_accum_1_U0_accum_out_we0),
    .accum_out_d0(tdf6_accum_1_U0_accum_out_d0),
    .accum_out_address1(tdf6_accum_1_U0_accum_out_address1),
    .accum_out_ce1(tdf6_accum_1_U0_accum_out_ce1),
    .accum_out_we1(tdf6_accum_1_U0_accum_out_we1),
    .accum_out_d1(tdf6_accum_1_U0_accum_out_d1)
);

td_fused_top_tdf6_accum_2 tdf6_accum_2_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf6_accum_2_U0_ap_start),
    .ap_done(tdf6_accum_2_U0_ap_done),
    .ap_continue(tdf6_accum_2_U0_ap_continue),
    .ap_idle(tdf6_accum_2_U0_ap_idle),
    .ap_ready(tdf6_accum_2_U0_ap_ready),
    .accum_in_8(tdf6_accum_2_U0_accum_in_8),
    .accum_in_8_ap_vld(tdf6_accum_2_U0_accum_in_8_ap_vld),
    .accum_in_address0(tdf6_accum_2_U0_accum_in_address0),
    .accum_in_ce0(tdf6_accum_2_U0_accum_in_ce0),
    .accum_in_q0(accum1_out_0_t_q0)
);

td_fused_top_Block_entry_proc_proc413 Block_entry_proc_proc413_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(Block_entry_proc_proc413_U0_ap_start),
    .ap_done(Block_entry_proc_proc413_U0_ap_done),
    .ap_continue(Block_entry_proc_proc413_U0_ap_continue),
    .ap_idle(Block_entry_proc_proc413_U0_ap_idle),
    .ap_ready(Block_entry_proc_proc413_U0_ap_ready),
    .tmp(tmp_channel_dout),
    .ap_return(Block_entry_proc_proc413_U0_ap_return)
);

td_fused_top_tdf6_adjust tdf6_adjust_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf6_adjust_U0_ap_start),
    .ap_done(tdf6_adjust_U0_ap_done),
    .ap_continue(tdf6_adjust_U0_ap_continue),
    .ap_idle(tdf6_adjust_U0_ap_idle),
    .ap_ready(tdf6_adjust_U0_ap_ready),
    .sums_read(sums_0_dout),
    .adjustments_address0(tdf6_adjust_U0_adjustments_address0),
    .adjustments_ce0(tdf6_adjust_U0_adjustments_ce0),
    .adjustments_q0(adjustments_q0),
    .indices_23_dout(indices_23_c1_dout),
    .indices_23_empty_n(indices_23_c1_empty_n),
    .indices_23_read(tdf6_adjust_U0_indices_23_read),
    .ap_return(tdf6_adjust_U0_ap_return)
);

td_fused_top_tdf6_writeOutputs_unaligned tdf6_writeOutputs_unaligned_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf6_writeOutputs_unaligned_U0_ap_start),
    .ap_done(tdf6_writeOutputs_unaligned_U0_ap_done),
    .ap_continue(tdf6_writeOutputs_unaligned_U0_ap_continue),
    .ap_idle(tdf6_writeOutputs_unaligned_U0_ap_idle),
    .ap_ready(tdf6_writeOutputs_unaligned_U0_ap_ready),
    .indices_01_dout(indices_01_c2_dout),
    .indices_01_empty_n(indices_01_c2_empty_n),
    .indices_01_read(tdf6_writeOutputs_unaligned_U0_indices_01_read),
    .indices_12_dout(indices_12_c3_dout),
    .indices_12_empty_n(indices_12_c3_empty_n),
    .indices_12_read(tdf6_writeOutputs_unaligned_U0_indices_12_read),
    .p_read(outputs_0_dout),
    .out_data_address1(tdf6_writeOutputs_unaligned_U0_out_data_address1),
    .out_data_ce1(tdf6_writeOutputs_unaligned_U0_out_data_ce1),
    .out_data_we1(tdf6_writeOutputs_unaligned_U0_out_data_we1),
    .out_data_d1(tdf6_writeOutputs_unaligned_U0_out_data_d1)
);

td_fused_top_fifo_w16_d2_S_x3 indices_01_c_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(indices_01_c_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf6_readInputs_U0_indices_01_read),
    .if_dout(indices_01_c_dout),
    .if_full_n(indices_01_c_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf6_get_next_ijk_U0_indices_0_write),
    .if_din(tdf6_get_next_ijk_U0_indices_0_din)
);

td_fused_top_fifo_w16_d2_S_x3 indices_12_c_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(indices_12_c_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf6_readInputs_U0_indices_12_read),
    .if_dout(indices_12_c_dout),
    .if_full_n(indices_12_c_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf6_get_next_ijk_U0_indices_1_write),
    .if_din(tdf6_get_next_ijk_U0_indices_1_din)
);

td_fused_top_fifo_w5_d2_S_x indices_23_c_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(indices_23_c_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf6_readFilters46_U0_indices_23_read),
    .if_dout(indices_23_c_dout),
    .if_full_n(indices_23_c_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf6_get_next_ijk_U0_indices_2_out_write),
    .if_din(tdf6_get_next_ijk_U0_indices_2_out_din)
);

td_fused_top_fifo_w5_d7_S_x indices_23_c1_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(indices_23_c1_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf6_adjust_U0_indices_23_read),
    .if_dout(indices_23_c1_dout),
    .if_full_n(indices_23_c1_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf6_get_next_ijk_U0_indices_2_out1_write),
    .if_din(tdf6_get_next_ijk_U0_indices_2_out1_din)
);

td_fused_top_fifo_w5_d7_S_x indices_01_c2_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(indices_01_c2_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf6_writeOutputs_unaligned_U0_indices_01_read),
    .if_dout(indices_01_c2_dout),
    .if_full_n(indices_01_c2_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf6_readInputs_U0_indices_01_out_write),
    .if_din(tdf6_readInputs_U0_indices_01_out_din)
);

td_fused_top_fifo_w10_d7_S indices_12_c3_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(indices_12_c3_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf6_writeOutputs_unaligned_U0_indices_12_read),
    .if_dout(indices_12_c3_dout),
    .if_full_n(indices_12_c3_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf6_readInputs_U0_indices_12_out_write),
    .if_din(tdf6_readInputs_U0_indices_12_out_din)
);

td_fused_top_fifo_w16_d2_S_x3 tmp_channel_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(tmp_channel_empty_n),
    .if_read_ce(1'b1),
    .if_read(Block_entry_proc_proc413_U0_ap_ready),
    .if_dout(tmp_channel_dout),
    .if_full_n(tmp_channel_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf6_accum_2_U0_ap_done),
    .if_din(tdf6_accum_2_U0_accum_in_8)
);

td_fused_top_fifo_w16_d2_S_x3 sums_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(sums_0_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf6_adjust_U0_ap_ready),
    .if_dout(sums_0_dout),
    .if_full_n(sums_0_full_n),
    .if_write_ce(1'b1),
    .if_write(Block_entry_proc_proc413_U0_ap_done),
    .if_din(Block_entry_proc_proc413_U0_ap_return)
);

td_fused_top_fifo_w16_d2_S_x3 outputs_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(outputs_0_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf6_writeOutputs_unaligned_U0_ap_ready),
    .if_dout(outputs_0_dout),
    .if_full_n(outputs_0_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf6_adjust_U0_ap_done),
    .if_din(tdf6_adjust_U0_ap_return)
);

td_fused_top_start_for_tdf6_readFilters46_U0 start_for_tdf6_readFilters46_U0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(start_for_tdf6_readFilters46_U0_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf6_readFilters46_U0_ap_ready),
    .if_dout(start_for_tdf6_readFilters46_U0_dout),
    .if_full_n(start_for_tdf6_readFilters46_U0_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf6_get_next_ijk_U0_start_write),
    .if_din(start_for_tdf6_readFilters46_U0_din)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_sync_reg_tdf6_get_next_ijk_U0_ap_ready <= 1'b0;
    end else begin
        if (((ap_sync_ready & ap_start) == 1'b1)) begin
            ap_sync_reg_tdf6_get_next_ijk_U0_ap_ready <= 1'b0;
        end else begin
            ap_sync_reg_tdf6_get_next_ijk_U0_ap_ready <= ap_sync_tdf6_get_next_ijk_U0_ap_ready;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_sync_reg_tdf6_readInputs_U0_ap_ready <= 1'b0;
    end else begin
        if (((ap_sync_ready & ap_start) == 1'b1)) begin
            ap_sync_reg_tdf6_readInputs_U0_ap_ready <= 1'b0;
        end else begin
            ap_sync_reg_tdf6_readInputs_U0_ap_ready <= ap_sync_tdf6_readInputs_U0_ap_ready;
        end
    end
end

assign Block_entry_proc_proc413_U0_ap_continue = sums_0_full_n;

assign Block_entry_proc_proc413_U0_ap_start = tmp_channel_empty_n;

assign Block_entry_proc_proc413_U0_start_full_n = 1'b1;

assign Block_entry_proc_proc413_U0_start_write = 1'b0;

assign adjustments_address0 = tdf6_adjust_U0_adjustments_address0;

assign adjustments_address1 = 5'd0;

assign adjustments_ce0 = tdf6_adjust_U0_adjustments_ce0;

assign adjustments_ce1 = 1'b0;

assign adjustments_d0 = 48'd0;

assign adjustments_d1 = 48'd0;

assign adjustments_we0 = 1'b0;

assign adjustments_we1 = 1'b0;

assign ap_channel_done_accum1_out_0 = tdf6_accum_1_U0_ap_done;

assign ap_channel_done_ifmap_vec_0_0 = tdf6_readInputs_U0_ap_done;

assign ap_channel_done_outputs_0 = tdf6_adjust_U0_ap_done;

assign ap_channel_done_products_0 = tdf6_dot_product_U0_ap_done;

assign ap_channel_done_sums_0 = Block_entry_proc_proc413_U0_ap_done;

assign ap_channel_done_tmp_channel = tdf6_accum_2_U0_ap_done;

assign ap_channel_done_weight_vecs_0_0_0 = tdf6_readFilters46_U0_ap_done;

assign ap_done = tdf6_writeOutputs_unaligned_U0_ap_done;

assign ap_idle = (tdf6_writeOutputs_unaligned_U0_ap_idle & tdf6_readInputs_U0_ap_idle & tdf6_readFilters46_U0_ap_idle & tdf6_get_next_ijk_U0_ap_idle & tdf6_dot_product_U0_ap_idle & tdf6_adjust_U0_ap_idle & tdf6_accum_2_U0_ap_idle & tdf6_accum_1_U0_ap_idle & (outputs_0_empty_n ^ 1'b1) & (sums_0_empty_n ^ 1'b1) & (tmp_channel_empty_n ^ 1'b1) & (products_0_t_empty_n ^ 1'b1) & (weight_vecs_0_0_0_t_empty_n ^ 1'b1) & (ifmap_vec_0_0_t_empty_n ^ 1'b1) & (1'b1 ^ accum1_out_0_t_empty_n) & Block_entry_proc_proc413_U0_ap_idle);

assign ap_ready = ap_sync_ready;

assign ap_sync_continue = ap_continue;

assign ap_sync_done = tdf6_writeOutputs_unaligned_U0_ap_done;

assign ap_sync_ready = (ap_sync_tdf6_readInputs_U0_ap_ready & ap_sync_tdf6_get_next_ijk_U0_ap_ready);

assign ap_sync_tdf6_get_next_ijk_U0_ap_ready = (tdf6_get_next_ijk_U0_ap_ready | ap_sync_reg_tdf6_get_next_ijk_U0_ap_ready);

assign ap_sync_tdf6_readInputs_U0_ap_ready = (tdf6_readInputs_U0_ap_ready | ap_sync_reg_tdf6_readInputs_U0_ap_ready);

assign filter_data_address0 = tdf6_readFilters46_U0_filter_data_address0;

assign filter_data_address1 = 12'd0;

assign filter_data_ce0 = tdf6_readFilters46_U0_filter_data_ce0;

assign filter_data_ce1 = 1'b0;

assign filter_data_d0 = 16'd0;

assign filter_data_d1 = 16'd0;

assign filter_data_we0 = 1'b0;

assign filter_data_we1 = 1'b0;

assign in_data_address0 = tdf6_readInputs_U0_in_data_address0;

assign in_data_address1 = 15'd0;

assign in_data_ce0 = tdf6_readInputs_U0_in_data_ce0;

assign in_data_ce1 = 1'b0;

assign in_data_d0 = 64'd0;

assign in_data_d1 = 64'd0;

assign in_data_read = tdf6_readInputs_U0_in_data_write;

assign in_data_we0 = 1'b0;

assign in_data_we1 = 1'b0;

assign out_data_address0 = 13'd0;

assign out_data_address1 = tdf6_writeOutputs_unaligned_U0_out_data_address1;

assign out_data_ce0 = 1'b0;

assign out_data_ce1 = tdf6_writeOutputs_unaligned_U0_out_data_ce1;

assign out_data_d0 = 64'd0;

assign out_data_d1 = tdf6_writeOutputs_unaligned_U0_out_data_d1;

assign out_data_we0 = 1'b0;

assign out_data_we1 = tdf6_writeOutputs_unaligned_U0_out_data_we1;

assign out_data_write = tdf6_writeOutputs_unaligned_U0_out_data_write;

assign products_0_t_d1 = 16'd0;

assign products_0_t_we1 = 1'b0;

assign start_for_tdf6_readFilters46_U0_din = 1'b1;

assign tdf6_accum_1_U0_accum_out_full_n = accum1_out_0_i_full_n;

assign tdf6_accum_1_U0_ap_continue = accum1_out_0_i_full_n;

assign tdf6_accum_1_U0_ap_start = products_0_t_empty_n;

assign tdf6_accum_1_U0_start_full_n = 1'b1;

assign tdf6_accum_1_U0_start_write = 1'b0;

assign tdf6_accum_2_U0_ap_continue = tmp_channel_full_n;

assign tdf6_accum_2_U0_ap_start = accum1_out_0_t_empty_n;

assign tdf6_accum_2_U0_start_full_n = 1'b1;

assign tdf6_accum_2_U0_start_write = 1'b0;

assign tdf6_adjust_U0_ap_continue = outputs_0_full_n;

assign tdf6_adjust_U0_ap_start = sums_0_empty_n;

assign tdf6_adjust_U0_start_full_n = 1'b1;

assign tdf6_adjust_U0_start_write = 1'b0;

assign tdf6_dot_product_U0_ap_continue = products_0_i_full_n;

assign tdf6_dot_product_U0_ap_start = (weight_vecs_0_0_0_t_empty_n & ifmap_vec_0_0_t_empty_n);

assign tdf6_dot_product_U0_products_0_full_n = products_0_i_full_n;

assign tdf6_dot_product_U0_start_full_n = 1'b1;

assign tdf6_dot_product_U0_start_write = 1'b0;

assign tdf6_get_next_ijk_U0_ap_continue = 1'b1;

assign tdf6_get_next_ijk_U0_ap_start = ((ap_sync_reg_tdf6_get_next_ijk_U0_ap_ready ^ 1'b1) & ap_start);

assign tdf6_readFilters46_U0_ap_continue = weight_vecs_0_0_0_i_full_n;

assign tdf6_readFilters46_U0_ap_start = start_for_tdf6_readFilters46_U0_empty_n;

assign tdf6_readFilters46_U0_start_full_n = 1'b1;

assign tdf6_readFilters46_U0_start_write = 1'b0;

assign tdf6_readFilters46_U0_weight_vecs_0_0_0_full_n = weight_vecs_0_0_0_i_full_n;

assign tdf6_readInputs_U0_ap_continue = ifmap_vec_0_0_i_full_n;

assign tdf6_readInputs_U0_ap_start = ((ap_sync_reg_tdf6_readInputs_U0_ap_ready ^ 1'b1) & ap_start);

assign tdf6_readInputs_U0_ifmap_vec_0_0_full_n = ifmap_vec_0_0_i_full_n;

assign tdf6_readInputs_U0_in_data_full_n = in_data_empty_n;

assign tdf6_readInputs_U0_in_data_write = 1'b0;

assign tdf6_readInputs_U0_start_full_n = 1'b1;

assign tdf6_readInputs_U0_start_write = 1'b0;

assign tdf6_writeOutputs_unaligned_U0_ap_continue = ap_continue;

assign tdf6_writeOutputs_unaligned_U0_ap_start = outputs_0_empty_n;

assign tdf6_writeOutputs_unaligned_U0_out_data_full_n = out_data_full_n;

assign tdf6_writeOutputs_unaligned_U0_out_data_write = 1'b0;

assign tdf6_writeOutputs_unaligned_U0_start_full_n = 1'b1;

assign tdf6_writeOutputs_unaligned_U0_start_write = 1'b0;

endmodule //td_fused_top_dataflow_in_loop_TOP_LOOP37644
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37644_weight_vecs_0_0_0_memcore_ram (addr0, ce0, d0, we0, q0, addr1, ce1, d1, we1, q1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 8;
parameter MEM_SIZE = 256;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
output reg[DWIDTH-1:0] q1;
input clk;

reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];




always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1) 
            ram[addr1] <= d1; 
        q1 <= ram[addr1];
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37644_weight_vecs_0_0_0_memcore(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    q0,
    address1,
    ce1,
    we1,
    d1,
    q1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd256;
parameter AddressWidth = 32'd8;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;
output[DataWidth - 1:0] q1;



td_fused_top_dataflow_in_loop_TOP_LOOP37644_weight_vecs_0_0_0_memcore_ram td_fused_top_dataflow_in_loop_TOP_LOOP37644_weight_vecs_0_0_0_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 ),
    .q1( q1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_dataflow_in_loop_TOP_LOOP37644_weight_vecs_0_0_0
#(parameter
    DataWidth    = 16,
    AddressRange = 32,
    AddressWidth = 7,
    BufferCount  = 2,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire                    i_we0,
    input  wire [AddressWidth-1:0] i_address0,
    input  wire [DataWidth-1:0]    i_d0,
    output wire [DataWidth-1:0]    i_q0,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire                    t_we0,
    input  wire [AddressWidth-1:0] t_address0,
    input  wire [DataWidth-1:0]    t_d0,
    output wire [DataWidth-1:0]    t_q0
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
wire [AddressWidth+IndexWidth-1:0]   memcore_iaddr;
wire [AddressWidth+IndexWidth-1:0]   memcore_taddr;

//------------------------Instantiation------------------
assign memcore_iaddr = {i_address0, iptr};
assign memcore_taddr = {t_address0, tptr};
td_fused_top_dataflow_in_loop_TOP_LOOP37644_weight_vecs_0_0_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP37644_weight_vecs_0_0_0_memcore_U (
    .reset    ( reset ),
    .clk      ( clk ),
    .address0 ( memcore_iaddr ),
    .ce0      ( i_ce0 ),
    .we0      ( i_we0),
    .d0       ( i_d0 ),
    .q0       ( i_q0 ),
    .address1 ( memcore_taddr ),
    .ce1      ( t_ce0 ),
    .we1      ( t_we0),
    .d1       ( t_d0 ),
    .q1       ( t_q0 )

);

//------------------------Body---------------------------

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37738_accum1_out_0_memcore_ram (addr0, ce0, d0, we0, q0, addr1, ce1, d1, we1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 3;
parameter MEM_SIZE = 8;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
input clk;

reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];




always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1) 
            ram[addr1] <= d1; 
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37738_accum1_out_0_memcore(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    q0,
    address1,
    ce1,
    we1,
    d1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd8;
parameter AddressWidth = 32'd3;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;



td_fused_top_dataflow_in_loop_TOP_LOOP37738_accum1_out_0_memcore_ram td_fused_top_dataflow_in_loop_TOP_LOOP37738_accum1_out_0_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_dataflow_in_loop_TOP_LOOP37738_accum1_out_0
#(parameter
    DataWidth    = 16,
    AddressRange = 32,
    AddressWidth = 3,
    BufferCount  = 2,
    MemLatency   = 1,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire                    i_we0,
    input  wire [AddressWidth-1:0] i_address0,
    input  wire [DataWidth-1:0]    i_d0,
    output wire [DataWidth-1:0]    i_q0,
    input  wire                    i_ce1,
    input  wire                    i_we1,
    input  wire [AddressWidth-1:0] i_address1,
    input  wire [DataWidth-1:0]    i_d1,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire                    t_we0,
    input  wire [AddressWidth-1:0] t_address0,
    input  wire [DataWidth-1:0]    t_d0,
    output wire [DataWidth-1:0]    t_q0,
    input  wire                    t_ce1,
    input  wire                    t_we1,
    input  wire [AddressWidth-1:0] t_address1,
    input  wire [DataWidth-1:0]    t_d1
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth-1:0]   prev_iptr    = 1'b0; // previous initiator index
reg  [IndexWidth-1:0]   prev_tptr    = 1'b0; // previous target index
reg  [DataWidth-1:0]    reg_q0      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid0    = 1'b0; // buffer has valid data
reg  [DataWidth-1:0]    reg_q1      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid1    = 1'b0; // buffer has valid data
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
// buffer signals
wire [BufferCount-1:0] buf_ce0;
wire [BufferCount-1:0] buf_we0;
wire [AddressWidth-1:0] buf_a0_0, buf_a0_1;
wire [DataWidth-1:0] buf_d0_0, buf_d0_1;
wire [DataWidth-1:0] buf_q0_0, buf_q0_1;
wire [BufferCount-1:0] buf_ce1;
wire [BufferCount-1:0] buf_we1;
wire [AddressWidth-1:0] buf_a1_0, buf_a1_1;
wire [DataWidth-1:0] buf_d1_0, buf_d1_1;
//------------------------Instantiation------------------
//genvar i;
        td_fused_top_dataflow_in_loop_TOP_LOOP37738_accum1_out_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP37738_accum1_out_0_memcore_U_0 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_0 ),
            .ce0      ( buf_ce0[ 0 ] ),
            .we0      ( buf_we0[ 0 ] ),
            .d0       ( buf_d0_0 ),
            .q0       ( buf_q0_0 ),
            .address1 ( buf_a1_0 ),
            .ce1      ( buf_ce1[ 0 ] ),
            .we1      ( buf_we1[ 0 ] ),
            .d1       ( buf_d1_0 )
        );
        td_fused_top_dataflow_in_loop_TOP_LOOP37738_accum1_out_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP37738_accum1_out_0_memcore_U_1 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_1 ),
            .ce0      ( buf_ce0[ 1 ] ),
            .we0      ( buf_we0[ 1 ] ),
            .d0       ( buf_d0_1 ),
            .q0       ( buf_q0_1 ),
            .address1 ( buf_a1_1 ),
            .ce1      ( buf_ce1[ 1 ] ),
            .we1      ( buf_we1[ 1 ] ),
            .d1       ( buf_d1_1 )
        );

//++++++++++++++++++++++++buffer signals+++++++++++++++++
        assign buf_ce0[ 0 ] = (tptr ==  0  && empty_n) ? t_ce0
                             : (iptr ==  0 ) ? i_ce0 : 1'b0;
        assign buf_a0_0  = (tptr ==  0  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 0 ] = (tptr ==  0  && empty_n)  ? t_we0
                             : (iptr ==  0 ) ? i_we0 : 1'b0;
        assign buf_d0_0  = (tptr ==  0  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 0 ] = (tptr ==  0  && empty_n) ? t_ce1
                             : (iptr ==  0 ) ? i_ce1 : 1'b0;
        assign buf_a1_0  = (tptr ==  0  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 0 ] = (tptr ==  0  && empty_n)  ? t_we1
                             : (iptr ==  0 ) ? i_we1 : 1'b0;
        assign buf_d1_0  = (tptr ==  0  && empty_n) ? t_d1       : i_d1;
        assign buf_ce0[ 1 ] = (tptr ==  1  && empty_n) ? t_ce0
                             : (iptr ==  1 ) ? i_ce0 : 1'b0;
        assign buf_a0_1  = (tptr ==  1  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 1 ] = (tptr ==  1  && empty_n)  ? t_we0
                             : (iptr ==  1 ) ? i_we0 : 1'b0;
        assign buf_d0_1  = (tptr ==  1  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 1 ] = (tptr ==  1  && empty_n) ? t_ce1
                             : (iptr ==  1 ) ? i_ce1 : 1'b0;
        assign buf_a1_1  = (tptr ==  1  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 1 ] = (tptr ==  1  && empty_n)  ? t_we1
                             : (iptr ==  1 ) ? i_we1 : 1'b0;
        assign buf_d1_1  = (tptr ==  1  && empty_n) ? t_d1       : i_d1;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//------------------------Body---------------------------
assign i_q0      = (prev_iptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign t_q0      = reg_valid0 ? reg_q0 : (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// prev_iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_iptr <= 1'b0;
    else begin
        prev_iptr <= iptr;
    end
end

// prev_tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_tptr <= 1'b0;
    else begin
        prev_tptr <= tptr;
    end
end

// reg_q0 and reg_valid0
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q0     <= 1'b0;
        reg_valid0 <= 1'b0;
    end else if (!t_ce0 && !reg_valid0) begin
        reg_q0     <= (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
        reg_valid0 <= 1'b1;
    end else if (t_ce0) begin
        reg_valid0 <= 1'b0;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37738_ifmap_vec_memcore_ram (addr0, ce0, d0, we0, q0, addr1, ce1, d1, we1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 8;
parameter MEM_SIZE = 144;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
input clk;

reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];




always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1) 
            ram[addr1] <= d1; 
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37738_ifmap_vec_memcore(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    q0,
    address1,
    ce1,
    we1,
    d1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd144;
parameter AddressWidth = 32'd8;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;



td_fused_top_dataflow_in_loop_TOP_LOOP37738_ifmap_vec_memcore_ram td_fused_top_dataflow_in_loop_TOP_LOOP37738_ifmap_vec_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_dataflow_in_loop_TOP_LOOP37738_ifmap_vec
#(parameter
    DataWidth    = 16,
    AddressRange = 32,
    AddressWidth = 8,
    BufferCount  = 2,
    MemLatency   = 1,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire                    i_we0,
    input  wire [AddressWidth-1:0] i_address0,
    input  wire [DataWidth-1:0]    i_d0,
    output wire [DataWidth-1:0]    i_q0,
    input  wire                    i_ce1,
    input  wire                    i_we1,
    input  wire [AddressWidth-1:0] i_address1,
    input  wire [DataWidth-1:0]    i_d1,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire                    t_we0,
    input  wire [AddressWidth-1:0] t_address0,
    input  wire [DataWidth-1:0]    t_d0,
    output wire [DataWidth-1:0]    t_q0,
    input  wire                    t_ce1,
    input  wire                    t_we1,
    input  wire [AddressWidth-1:0] t_address1,
    input  wire [DataWidth-1:0]    t_d1
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth-1:0]   prev_iptr    = 1'b0; // previous initiator index
reg  [IndexWidth-1:0]   prev_tptr    = 1'b0; // previous target index
reg  [DataWidth-1:0]    reg_q0      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid0    = 1'b0; // buffer has valid data
reg  [DataWidth-1:0]    reg_q1      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid1    = 1'b0; // buffer has valid data
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
// buffer signals
wire [BufferCount-1:0] buf_ce0;
wire [BufferCount-1:0] buf_we0;
wire [AddressWidth-1:0] buf_a0_0, buf_a0_1;
wire [DataWidth-1:0] buf_d0_0, buf_d0_1;
wire [DataWidth-1:0] buf_q0_0, buf_q0_1;
wire [BufferCount-1:0] buf_ce1;
wire [BufferCount-1:0] buf_we1;
wire [AddressWidth-1:0] buf_a1_0, buf_a1_1;
wire [DataWidth-1:0] buf_d1_0, buf_d1_1;
//------------------------Instantiation------------------
//genvar i;
        td_fused_top_dataflow_in_loop_TOP_LOOP37738_ifmap_vec_memcore td_fused_top_dataflow_in_loop_TOP_LOOP37738_ifmap_vec_memcore_U_0 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_0 ),
            .ce0      ( buf_ce0[ 0 ] ),
            .we0      ( buf_we0[ 0 ] ),
            .d0       ( buf_d0_0 ),
            .q0       ( buf_q0_0 ),
            .address1 ( buf_a1_0 ),
            .ce1      ( buf_ce1[ 0 ] ),
            .we1      ( buf_we1[ 0 ] ),
            .d1       ( buf_d1_0 )
        );
        td_fused_top_dataflow_in_loop_TOP_LOOP37738_ifmap_vec_memcore td_fused_top_dataflow_in_loop_TOP_LOOP37738_ifmap_vec_memcore_U_1 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_1 ),
            .ce0      ( buf_ce0[ 1 ] ),
            .we0      ( buf_we0[ 1 ] ),
            .d0       ( buf_d0_1 ),
            .q0       ( buf_q0_1 ),
            .address1 ( buf_a1_1 ),
            .ce1      ( buf_ce1[ 1 ] ),
            .we1      ( buf_we1[ 1 ] ),
            .d1       ( buf_d1_1 )
        );

//++++++++++++++++++++++++buffer signals+++++++++++++++++
        assign buf_ce0[ 0 ] = (tptr ==  0  && empty_n) ? t_ce0
                             : (iptr ==  0 ) ? i_ce0 : 1'b0;
        assign buf_a0_0  = (tptr ==  0  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 0 ] = (tptr ==  0  && empty_n)  ? t_we0
                             : (iptr ==  0 ) ? i_we0 : 1'b0;
        assign buf_d0_0  = (tptr ==  0  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 0 ] = (tptr ==  0  && empty_n) ? t_ce1
                             : (iptr ==  0 ) ? i_ce1 : 1'b0;
        assign buf_a1_0  = (tptr ==  0  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 0 ] = (tptr ==  0  && empty_n)  ? t_we1
                             : (iptr ==  0 ) ? i_we1 : 1'b0;
        assign buf_d1_0  = (tptr ==  0  && empty_n) ? t_d1       : i_d1;
        assign buf_ce0[ 1 ] = (tptr ==  1  && empty_n) ? t_ce0
                             : (iptr ==  1 ) ? i_ce0 : 1'b0;
        assign buf_a0_1  = (tptr ==  1  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 1 ] = (tptr ==  1  && empty_n)  ? t_we0
                             : (iptr ==  1 ) ? i_we0 : 1'b0;
        assign buf_d0_1  = (tptr ==  1  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 1 ] = (tptr ==  1  && empty_n) ? t_ce1
                             : (iptr ==  1 ) ? i_ce1 : 1'b0;
        assign buf_a1_1  = (tptr ==  1  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 1 ] = (tptr ==  1  && empty_n)  ? t_we1
                             : (iptr ==  1 ) ? i_we1 : 1'b0;
        assign buf_d1_1  = (tptr ==  1  && empty_n) ? t_d1       : i_d1;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//------------------------Body---------------------------
assign i_q0      = (prev_iptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign t_q0      = reg_valid0 ? reg_q0 : (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// prev_iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_iptr <= 1'b0;
    else begin
        prev_iptr <= iptr;
    end
end

// prev_tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_tptr <= 1'b0;
    else begin
        prev_tptr <= tptr;
    end
end

// reg_q0 and reg_valid0
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q0     <= 1'b0;
        reg_valid0 <= 1'b0;
    end else if (!t_ce0 && !reg_valid0) begin
        reg_q0     <= (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
        reg_valid0 <= 1'b1;
    end else if (t_ce0) begin
        reg_valid0 <= 1'b0;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37738_products_0_memcore_ram (addr0, ce0, d0, we0, q0, addr1, ce1, q1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 8;
parameter MEM_SIZE = 144;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
output reg[DWIDTH-1:0] q1;
input clk;

reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];




always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        q1 <= ram[addr1];
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37738_products_0_memcore(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    q0,
    address1,
    ce1,
    q1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd144;
parameter AddressWidth = 32'd8;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
output[DataWidth - 1:0] q1;



td_fused_top_dataflow_in_loop_TOP_LOOP37738_products_0_memcore_ram td_fused_top_dataflow_in_loop_TOP_LOOP37738_products_0_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .q1( q1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_dataflow_in_loop_TOP_LOOP37738_products_0
#(parameter
    DataWidth    = 16,
    AddressRange = 32,
    AddressWidth = 8,
    BufferCount  = 2,
    MemLatency   = 1,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire                    i_we0,
    input  wire [AddressWidth-1:0] i_address0,
    input  wire [DataWidth-1:0]    i_d0,
    output wire [DataWidth-1:0]    i_q0,
    input  wire                    i_ce1,
    input  wire [AddressWidth-1:0] i_address1,
    output wire [DataWidth-1:0]    i_q1,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire                    t_we0,
    input  wire [AddressWidth-1:0] t_address0,
    input  wire [DataWidth-1:0]    t_d0,
    output wire [DataWidth-1:0]    t_q0,
    input  wire                    t_ce1,
    input  wire [AddressWidth-1:0] t_address1,
    output wire [DataWidth-1:0]    t_q1
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth-1:0]   prev_iptr    = 1'b0; // previous initiator index
reg  [IndexWidth-1:0]   prev_tptr    = 1'b0; // previous target index
reg  [DataWidth-1:0]    reg_q0      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid0    = 1'b0; // buffer has valid data
reg  [DataWidth-1:0]    reg_q1      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid1    = 1'b0; // buffer has valid data
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
// buffer signals
wire [BufferCount-1:0] buf_ce0;
wire [BufferCount-1:0] buf_we0;
wire [AddressWidth-1:0] buf_a0_0, buf_a0_1;
wire [DataWidth-1:0] buf_d0_0, buf_d0_1;
wire [DataWidth-1:0] buf_q0_0, buf_q0_1;
wire [BufferCount-1:0] buf_ce1;
wire [AddressWidth-1:0] buf_a1_0, buf_a1_1;
wire [DataWidth-1:0] buf_q1_0, buf_q1_1;
//------------------------Instantiation------------------
//genvar i;
        td_fused_top_dataflow_in_loop_TOP_LOOP37738_products_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP37738_products_0_memcore_U_0 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_0 ),
            .ce0      ( buf_ce0[ 0 ] ),
            .we0      ( buf_we0[ 0 ] ),
            .d0       ( buf_d0_0 ),
            .q0       ( buf_q0_0 ),
            .address1 ( buf_a1_0 ),
            .ce1      ( buf_ce1[ 0 ] ),
            .q1       ( buf_q1_0 )
        );
        td_fused_top_dataflow_in_loop_TOP_LOOP37738_products_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP37738_products_0_memcore_U_1 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_1 ),
            .ce0      ( buf_ce0[ 1 ] ),
            .we0      ( buf_we0[ 1 ] ),
            .d0       ( buf_d0_1 ),
            .q0       ( buf_q0_1 ),
            .address1 ( buf_a1_1 ),
            .ce1      ( buf_ce1[ 1 ] ),
            .q1       ( buf_q1_1 )
        );

//++++++++++++++++++++++++buffer signals+++++++++++++++++
        assign buf_ce0[ 0 ] = (tptr ==  0  && empty_n) ? t_ce0
                             : (iptr ==  0 ) ? i_ce0 : 1'b0;
        assign buf_a0_0  = (tptr ==  0  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 0 ] = (tptr ==  0  && empty_n)  ? t_we0
                             : (iptr ==  0 ) ? i_we0 : 1'b0;
        assign buf_d0_0  = (tptr ==  0  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 0 ] = (tptr ==  0  && empty_n) ? t_ce1
                             : (iptr ==  0 ) ? i_ce1 : 1'b0;
        assign buf_a1_0  = (tptr ==  0  && empty_n) ?  t_address1 : i_address1;
        assign buf_ce0[ 1 ] = (tptr ==  1  && empty_n) ? t_ce0
                             : (iptr ==  1 ) ? i_ce0 : 1'b0;
        assign buf_a0_1  = (tptr ==  1  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 1 ] = (tptr ==  1  && empty_n)  ? t_we0
                             : (iptr ==  1 ) ? i_we0 : 1'b0;
        assign buf_d0_1  = (tptr ==  1  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 1 ] = (tptr ==  1  && empty_n) ? t_ce1
                             : (iptr ==  1 ) ? i_ce1 : 1'b0;
        assign buf_a1_1  = (tptr ==  1  && empty_n) ?  t_address1 : i_address1;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//------------------------Body---------------------------
assign i_q0      = (prev_iptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign t_q0      = reg_valid0 ? reg_q0 : (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign i_q1      = (prev_iptr == 1'b1 ? buf_q1_1 : buf_q1_0);
assign t_q1      = reg_valid1 ? reg_q1 : (prev_tptr == 1'b1 ? buf_q1_1 : buf_q1_0);

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// prev_iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_iptr <= 1'b0;
    else begin
        prev_iptr <= iptr;
    end
end

// prev_tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_tptr <= 1'b0;
    else begin
        prev_tptr <= tptr;
    end
end

// reg_q0 and reg_valid0
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q0     <= 1'b0;
        reg_valid0 <= 1'b0;
    end else if (!t_ce0 && !reg_valid0) begin
        reg_q0     <= (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
        reg_valid0 <= 1'b1;
    end else if (t_ce0) begin
        reg_valid0 <= 1'b0;
    end
end

// reg_q1 and reg_valid1
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q1     <= 1'b0;
        reg_valid1 <= 1'b0;
    end else if (!t_ce1 && !reg_valid1) begin
        reg_q1     <= (prev_tptr == 1'b1 ? buf_q1_1 : buf_q1_0);
        reg_valid1 <= 1'b1;
    end else if (t_ce1) begin
        reg_valid1 <= 1'b0;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_dataflow_in_loop_TOP_LOOP37738 (
        ap_clk,
        ap_rst,
        in_data_address0,
        in_data_ce0,
        in_data_d0,
        in_data_q0,
        in_data_we0,
        in_data_address1,
        in_data_ce1,
        in_data_d1,
        in_data_q1,
        in_data_we1,
        filter_data_address0,
        filter_data_ce0,
        filter_data_d0,
        filter_data_q0,
        filter_data_we0,
        filter_data_address1,
        filter_data_ce1,
        filter_data_d1,
        filter_data_q1,
        filter_data_we1,
        adjustments_address0,
        adjustments_ce0,
        adjustments_d0,
        adjustments_q0,
        adjustments_we0,
        adjustments_address1,
        adjustments_ce1,
        adjustments_d1,
        adjustments_q1,
        adjustments_we1,
        out_data_address0,
        out_data_ce0,
        out_data_d0,
        out_data_q0,
        out_data_we0,
        out_data_address1,
        out_data_ce1,
        out_data_d1,
        out_data_q1,
        out_data_we1,
        ap_start,
        in_data_empty_n,
        in_data_read,
        out_data_full_n,
        out_data_write,
        ap_done,
        ap_ready,
        ap_idle,
        ap_continue
);


input   ap_clk;
input   ap_rst;
output  [13:0] in_data_address0;
output   in_data_ce0;
output  [63:0] in_data_d0;
input  [63:0] in_data_q0;
output   in_data_we0;
output  [13:0] in_data_address1;
output   in_data_ce1;
output  [63:0] in_data_d1;
input  [63:0] in_data_q1;
output   in_data_we1;
output  [14:0] filter_data_address0;
output   filter_data_ce0;
output  [15:0] filter_data_d0;
input  [15:0] filter_data_q0;
output   filter_data_we0;
output  [14:0] filter_data_address1;
output   filter_data_ce1;
output  [15:0] filter_data_d1;
input  [15:0] filter_data_q1;
output   filter_data_we1;
output  [6:0] adjustments_address0;
output   adjustments_ce0;
output  [47:0] adjustments_d0;
input  [47:0] adjustments_q0;
output   adjustments_we0;
output  [6:0] adjustments_address1;
output   adjustments_ce1;
output  [47:0] adjustments_d1;
input  [47:0] adjustments_q1;
output   adjustments_we1;
output  [14:0] out_data_address0;
output   out_data_ce0;
output  [63:0] out_data_d0;
input  [63:0] out_data_q0;
output   out_data_we0;
output  [14:0] out_data_address1;
output   out_data_ce1;
output  [63:0] out_data_d1;
input  [63:0] out_data_q1;
output   out_data_we1;
input   ap_start;
input   in_data_empty_n;
output   in_data_read;
input   out_data_full_n;
output   out_data_write;
output   ap_done;
output   ap_ready;
output   ap_idle;
input   ap_continue;

wire   [15:0] ifmap_vec_i_q0;
wire   [15:0] ifmap_vec_t_q0;
wire   [15:0] weight_vecs_0_i_q0;
wire   [15:0] weight_vecs_0_t_q0;
wire   [15:0] products_0_i_q0;
wire   [15:0] products_0_i_q1;
wire   [15:0] products_0_t_q0;
wire   [15:0] products_0_t_q1;
wire   [15:0] accum1_out_0_i_q0;
wire   [15:0] accum1_out_0_t_q0;
wire    tdf5_get_next_ijk_U0_ap_start;
wire    tdf5_get_next_ijk_U0_ap_done;
wire    tdf5_get_next_ijk_U0_ap_continue;
wire    tdf5_get_next_ijk_U0_ap_idle;
wire    tdf5_get_next_ijk_U0_ap_ready;
wire    tdf5_get_next_ijk_U0_start_out;
wire    tdf5_get_next_ijk_U0_start_write;
wire   [6:0] tdf5_get_next_ijk_U0_input_indices_2_out_din;
wire    tdf5_get_next_ijk_U0_input_indices_2_out_write;
wire   [6:0] tdf5_get_next_ijk_U0_input_indices_2_out1_din;
wire    tdf5_get_next_ijk_U0_input_indices_2_out1_write;
wire   [4:0] tdf5_get_next_ijk_U0_output_indices_0_din;
wire    tdf5_get_next_ijk_U0_output_indices_0_write;
wire   [9:0] tdf5_get_next_ijk_U0_output_indices_1_din;
wire    tdf5_get_next_ijk_U0_output_indices_1_write;
wire    tdf5_get_next_ijk_U0_resetMaximum_din;
wire    tdf5_get_next_ijk_U0_resetMaximum_write;
wire    tdf5_get_next_ijk_U0_storeOutput_din;
wire    tdf5_get_next_ijk_U0_storeOutput_write;
wire   [15:0] tdf5_get_next_ijk_U0_ap_return_0;
wire   [15:0] tdf5_get_next_ijk_U0_ap_return_1;
wire    ap_channel_done_input_indices_1;
wire    input_indices_1_full_n;
reg    ap_sync_reg_channel_write_input_indices_1;
wire    ap_sync_channel_write_input_indices_1;
wire    ap_channel_done_input_indices_0;
wire    input_indices_0_full_n;
reg    ap_sync_reg_channel_write_input_indices_0;
wire    ap_sync_channel_write_input_indices_0;
wire    tdf5_readInputs41_U0_ap_start;
wire    tdf5_readInputs41_U0_ap_done;
wire    tdf5_readInputs41_U0_ap_continue;
wire    tdf5_readInputs41_U0_ap_idle;
wire    tdf5_readInputs41_U0_ap_ready;
wire   [13:0] tdf5_readInputs41_U0_in_data_address0;
wire    tdf5_readInputs41_U0_in_data_ce0;
wire   [7:0] tdf5_readInputs41_U0_ifmap_vec_address0;
wire    tdf5_readInputs41_U0_ifmap_vec_ce0;
wire    tdf5_readInputs41_U0_ifmap_vec_we0;
wire   [15:0] tdf5_readInputs41_U0_ifmap_vec_d0;
wire   [7:0] tdf5_readInputs41_U0_ifmap_vec_address1;
wire    tdf5_readInputs41_U0_ifmap_vec_ce1;
wire    tdf5_readInputs41_U0_ifmap_vec_we1;
wire   [15:0] tdf5_readInputs41_U0_ifmap_vec_d1;
wire    tdf5_readInputs41_U0_in_data_full_n;
wire    tdf5_readInputs41_U0_in_data_write;
wire    ap_channel_done_ifmap_vec;
wire    tdf5_readInputs41_U0_ifmap_vec_full_n;
wire    tdf5_readFilters40_U0_ap_start;
wire    tdf5_readFilters40_U0_ap_done;
wire    tdf5_readFilters40_U0_ap_continue;
wire    tdf5_readFilters40_U0_ap_idle;
wire    tdf5_readFilters40_U0_ap_ready;
wire   [14:0] tdf5_readFilters40_U0_filter_data_address0;
wire    tdf5_readFilters40_U0_filter_data_ce0;
wire    tdf5_readFilters40_U0_input_indices_23_read;
wire   [7:0] tdf5_readFilters40_U0_weight_vecs_0_address0;
wire    tdf5_readFilters40_U0_weight_vecs_0_ce0;
wire    tdf5_readFilters40_U0_weight_vecs_0_we0;
wire   [15:0] tdf5_readFilters40_U0_weight_vecs_0_d0;
wire    ap_channel_done_weight_vecs_0;
wire    tdf5_readFilters40_U0_weight_vecs_0_full_n;
wire    tdf5_dot_product_U0_ap_start;
wire    tdf5_dot_product_U0_ap_done;
wire    tdf5_dot_product_U0_ap_continue;
wire    tdf5_dot_product_U0_ap_idle;
wire    tdf5_dot_product_U0_ap_ready;
wire   [7:0] tdf5_dot_product_U0_ifmap_vec_address0;
wire    tdf5_dot_product_U0_ifmap_vec_ce0;
wire   [7:0] tdf5_dot_product_U0_weight_vecs_0_address0;
wire    tdf5_dot_product_U0_weight_vecs_0_ce0;
wire   [7:0] tdf5_dot_product_U0_products_0_address0;
wire    tdf5_dot_product_U0_products_0_ce0;
wire    tdf5_dot_product_U0_products_0_we0;
wire   [15:0] tdf5_dot_product_U0_products_0_d0;
wire    ap_channel_done_products_0;
wire    tdf5_dot_product_U0_products_0_full_n;
wire    tdf5_accum_1_U0_ap_start;
wire    tdf5_accum_1_U0_ap_done;
wire    tdf5_accum_1_U0_ap_continue;
wire    tdf5_accum_1_U0_ap_idle;
wire    tdf5_accum_1_U0_ap_ready;
wire   [7:0] tdf5_accum_1_U0_accum_in_0_address0;
wire    tdf5_accum_1_U0_accum_in_0_ce0;
wire   [7:0] tdf5_accum_1_U0_accum_in_0_address1;
wire    tdf5_accum_1_U0_accum_in_0_ce1;
wire   [2:0] tdf5_accum_1_U0_accum_out_address0;
wire    tdf5_accum_1_U0_accum_out_ce0;
wire    tdf5_accum_1_U0_accum_out_we0;
wire   [15:0] tdf5_accum_1_U0_accum_out_d0;
wire   [2:0] tdf5_accum_1_U0_accum_out_address1;
wire    tdf5_accum_1_U0_accum_out_ce1;
wire    tdf5_accum_1_U0_accum_out_we1;
wire   [15:0] tdf5_accum_1_U0_accum_out_d1;
wire    ap_channel_done_accum1_out_0;
wire    tdf5_accum_1_U0_accum_out_full_n;
wire    tdf5_accum_2_U0_ap_start;
wire    tdf5_accum_2_U0_ap_done;
wire    tdf5_accum_2_U0_ap_continue;
wire    tdf5_accum_2_U0_ap_idle;
wire    tdf5_accum_2_U0_ap_ready;
wire   [15:0] tdf5_accum_2_U0_accum_in_10;
wire    tdf5_accum_2_U0_accum_in_10_ap_vld;
wire   [2:0] tdf5_accum_2_U0_accum_in_address0;
wire    tdf5_accum_2_U0_accum_in_ce0;
wire    ap_channel_done_tmp_channel;
wire    tmp_channel_full_n;
wire    Block_entry_proc_proc408_U0_ap_start;
wire    Block_entry_proc_proc408_U0_ap_done;
wire    Block_entry_proc_proc408_U0_ap_continue;
wire    Block_entry_proc_proc408_U0_ap_idle;
wire    Block_entry_proc_proc408_U0_ap_ready;
wire   [15:0] Block_entry_proc_proc408_U0_ap_return;
wire    ap_channel_done_sums_0;
wire    sums_0_full_n;
wire    tdf5_adjust_U0_ap_start;
wire    tdf5_adjust_U0_ap_done;
wire    tdf5_adjust_U0_ap_continue;
wire    tdf5_adjust_U0_ap_idle;
wire    tdf5_adjust_U0_ap_ready;
wire   [6:0] tdf5_adjust_U0_adjustments_address0;
wire    tdf5_adjust_U0_adjustments_ce0;
wire    tdf5_adjust_U0_input_indices_23_read;
wire   [15:0] tdf5_adjust_U0_ap_return;
wire    ap_channel_done_outputs_0;
wire    outputs_0_full_n;
wire    tdf5_poolOutputs_U0_ap_start;
wire    tdf5_poolOutputs_U0_ap_done;
wire    tdf5_poolOutputs_U0_ap_continue;
wire    tdf5_poolOutputs_U0_ap_idle;
wire    tdf5_poolOutputs_U0_ap_ready;
wire    tdf5_poolOutputs_U0_output_indices_04_read;
wire    tdf5_poolOutputs_U0_output_indices_15_read;
wire    tdf5_poolOutputs_U0_resetMaximum6_read;
wire    tdf5_poolOutputs_U0_storeOutput7_read;
wire   [14:0] tdf5_poolOutputs_U0_out_data_address1;
wire    tdf5_poolOutputs_U0_out_data_ce1;
wire    tdf5_poolOutputs_U0_out_data_we1;
wire   [63:0] tdf5_poolOutputs_U0_out_data_d1;
wire    tdf5_poolOutputs_U0_out_data_full_n;
wire    tdf5_poolOutputs_U0_out_data_write;
wire    ap_sync_continue;
wire    ifmap_vec_i_full_n;
wire    ifmap_vec_t_empty_n;
wire    weight_vecs_0_i_full_n;
wire    weight_vecs_0_t_empty_n;
wire    products_0_i_full_n;
wire    products_0_t_empty_n;
wire   [15:0] products_0_t_d1;
wire    products_0_t_we1;
wire    accum1_out_0_i_full_n;
wire    accum1_out_0_t_empty_n;
wire    input_indices_23_c_full_n;
wire   [6:0] input_indices_23_c_dout;
wire    input_indices_23_c_empty_n;
wire    input_indices_23_c1_full_n;
wire   [6:0] input_indices_23_c1_dout;
wire    input_indices_23_c1_empty_n;
wire    output_indices_04_c_full_n;
wire   [4:0] output_indices_04_c_dout;
wire    output_indices_04_c_empty_n;
wire    output_indices_15_c_full_n;
wire   [9:0] output_indices_15_c_dout;
wire    output_indices_15_c_empty_n;
wire   [0:0] resetMaximum6_c_din;
wire    resetMaximum6_c_full_n;
wire   [0:0] resetMaximum6_c_dout;
wire    resetMaximum6_c_empty_n;
wire   [0:0] storeOutput7_c_din;
wire    storeOutput7_c_full_n;
wire   [0:0] storeOutput7_c_dout;
wire    storeOutput7_c_empty_n;
wire   [15:0] input_indices_0_dout;
wire    input_indices_0_empty_n;
wire   [15:0] input_indices_1_dout;
wire    input_indices_1_empty_n;
wire   [15:0] tmp_channel_dout;
wire    tmp_channel_empty_n;
wire   [15:0] sums_0_dout;
wire    sums_0_empty_n;
wire   [15:0] outputs_0_dout;
wire    outputs_0_empty_n;
wire    ap_sync_done;
wire    ap_sync_ready;
reg    ap_sync_reg_tdf5_get_next_ijk_U0_ap_ready;
wire    ap_sync_tdf5_get_next_ijk_U0_ap_ready;
reg    ap_sync_reg_tdf5_readInputs41_U0_ap_ready;
wire    ap_sync_tdf5_readInputs41_U0_ap_ready;
wire   [0:0] start_for_tdf5_readFilters40_U0_din;
wire    start_for_tdf5_readFilters40_U0_full_n;
wire   [0:0] start_for_tdf5_readFilters40_U0_dout;
wire    start_for_tdf5_readFilters40_U0_empty_n;
wire    tdf5_readInputs41_U0_start_full_n;
wire    tdf5_readInputs41_U0_start_write;
wire    tdf5_readFilters40_U0_start_full_n;
wire    tdf5_readFilters40_U0_start_write;
wire    tdf5_dot_product_U0_start_full_n;
wire    tdf5_dot_product_U0_start_write;
wire    tdf5_accum_1_U0_start_full_n;
wire    tdf5_accum_1_U0_start_write;
wire    tdf5_accum_2_U0_start_full_n;
wire    tdf5_accum_2_U0_start_write;
wire    Block_entry_proc_proc408_U0_start_full_n;
wire    Block_entry_proc_proc408_U0_start_write;
wire    tdf5_adjust_U0_start_full_n;
wire    tdf5_adjust_U0_start_write;
wire    tdf5_poolOutputs_U0_start_full_n;
wire    tdf5_poolOutputs_U0_start_write;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_sync_reg_channel_write_input_indices_1 = 1'b0;
#0 ap_sync_reg_channel_write_input_indices_0 = 1'b0;
#0 ap_sync_reg_tdf5_get_next_ijk_U0_ap_ready = 1'b0;
#0 ap_sync_reg_tdf5_readInputs41_U0_ap_ready = 1'b0;
end

td_fused_top_dataflow_in_loop_TOP_LOOP37738_ifmap_vec #(
    .DataWidth( 16 ),
    .AddressRange( 144 ),
    .AddressWidth( 8 ))
ifmap_vec_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf5_readInputs41_U0_ap_done),
    .i_full_n(ifmap_vec_i_full_n),
    .i_ce0(tdf5_readInputs41_U0_ifmap_vec_ce0),
    .i_we0(tdf5_readInputs41_U0_ifmap_vec_we0),
    .i_address0(tdf5_readInputs41_U0_ifmap_vec_address0),
    .i_d0(tdf5_readInputs41_U0_ifmap_vec_d0),
    .i_q0(ifmap_vec_i_q0),
    .i_ce1(tdf5_readInputs41_U0_ifmap_vec_ce1),
    .i_we1(tdf5_readInputs41_U0_ifmap_vec_we1),
    .i_address1(tdf5_readInputs41_U0_ifmap_vec_address1),
    .i_d1(tdf5_readInputs41_U0_ifmap_vec_d1),
    .t_ce(1'b1),
    .t_read(tdf5_dot_product_U0_ap_ready),
    .t_empty_n(ifmap_vec_t_empty_n),
    .t_ce0(tdf5_dot_product_U0_ifmap_vec_ce0),
    .t_we0(1'b0),
    .t_address0(tdf5_dot_product_U0_ifmap_vec_address0),
    .t_d0(16'd0),
    .t_q0(ifmap_vec_t_q0),
    .t_ce1(1'b0),
    .t_we1(1'b0),
    .t_address1(8'd0),
    .t_d1(16'd0)
);

td_fused_top_dataflow_in_loop_TOP_LOOP37738_weight_vecs_0 #(
    .DataWidth( 16 ),
    .AddressRange( 144 ),
    .AddressWidth( 8 ))
weight_vecs_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf5_readFilters40_U0_ap_done),
    .i_full_n(weight_vecs_0_i_full_n),
    .i_ce0(tdf5_readFilters40_U0_weight_vecs_0_ce0),
    .i_we0(tdf5_readFilters40_U0_weight_vecs_0_we0),
    .i_address0(tdf5_readFilters40_U0_weight_vecs_0_address0),
    .i_d0(tdf5_readFilters40_U0_weight_vecs_0_d0),
    .i_q0(weight_vecs_0_i_q0),
    .t_ce(1'b1),
    .t_read(tdf5_dot_product_U0_ap_ready),
    .t_empty_n(weight_vecs_0_t_empty_n),
    .t_ce0(tdf5_dot_product_U0_weight_vecs_0_ce0),
    .t_we0(1'b0),
    .t_address0(tdf5_dot_product_U0_weight_vecs_0_address0),
    .t_d0(16'd0),
    .t_q0(weight_vecs_0_t_q0)
);

td_fused_top_dataflow_in_loop_TOP_LOOP37738_products_0 #(
    .DataWidth( 16 ),
    .AddressRange( 144 ),
    .AddressWidth( 8 ))
products_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf5_dot_product_U0_ap_done),
    .i_full_n(products_0_i_full_n),
    .i_ce0(tdf5_dot_product_U0_products_0_ce0),
    .i_we0(tdf5_dot_product_U0_products_0_we0),
    .i_address0(tdf5_dot_product_U0_products_0_address0),
    .i_d0(tdf5_dot_product_U0_products_0_d0),
    .i_q0(products_0_i_q0),
    .i_ce1(1'b0),
    .i_address1(8'd0),
    .i_q1(products_0_i_q1),
    .t_ce(1'b1),
    .t_read(tdf5_accum_1_U0_ap_ready),
    .t_empty_n(products_0_t_empty_n),
    .t_ce0(tdf5_accum_1_U0_accum_in_0_ce0),
    .t_we0(1'b0),
    .t_address0(tdf5_accum_1_U0_accum_in_0_address0),
    .t_d0(16'd0),
    .t_q0(products_0_t_q0),
    .t_ce1(tdf5_accum_1_U0_accum_in_0_ce1),
    .t_address1(tdf5_accum_1_U0_accum_in_0_address1),
    .t_q1(products_0_t_q1)
);

td_fused_top_dataflow_in_loop_TOP_LOOP37738_accum1_out_0 #(
    .DataWidth( 16 ),
    .AddressRange( 8 ),
    .AddressWidth( 3 ))
accum1_out_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf5_accum_1_U0_ap_done),
    .i_full_n(accum1_out_0_i_full_n),
    .i_ce0(tdf5_accum_1_U0_accum_out_ce0),
    .i_we0(tdf5_accum_1_U0_accum_out_we0),
    .i_address0(tdf5_accum_1_U0_accum_out_address0),
    .i_d0(tdf5_accum_1_U0_accum_out_d0),
    .i_q0(accum1_out_0_i_q0),
    .i_ce1(tdf5_accum_1_U0_accum_out_ce1),
    .i_we1(tdf5_accum_1_U0_accum_out_we1),
    .i_address1(tdf5_accum_1_U0_accum_out_address1),
    .i_d1(tdf5_accum_1_U0_accum_out_d1),
    .t_ce(1'b1),
    .t_read(tdf5_accum_2_U0_ap_ready),
    .t_empty_n(accum1_out_0_t_empty_n),
    .t_ce0(tdf5_accum_2_U0_accum_in_ce0),
    .t_we0(1'b0),
    .t_address0(tdf5_accum_2_U0_accum_in_address0),
    .t_d0(16'd0),
    .t_q0(accum1_out_0_t_q0),
    .t_ce1(1'b0),
    .t_we1(1'b0),
    .t_address1(3'd0),
    .t_d1(16'd0)
);

td_fused_top_tdf5_get_next_ijk tdf5_get_next_ijk_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf5_get_next_ijk_U0_ap_start),
    .start_full_n(start_for_tdf5_readFilters40_U0_full_n),
    .ap_done(tdf5_get_next_ijk_U0_ap_done),
    .ap_continue(tdf5_get_next_ijk_U0_ap_continue),
    .ap_idle(tdf5_get_next_ijk_U0_ap_idle),
    .ap_ready(tdf5_get_next_ijk_U0_ap_ready),
    .start_out(tdf5_get_next_ijk_U0_start_out),
    .start_write(tdf5_get_next_ijk_U0_start_write),
    .input_indices_2_out_din(tdf5_get_next_ijk_U0_input_indices_2_out_din),
    .input_indices_2_out_full_n(input_indices_23_c_full_n),
    .input_indices_2_out_write(tdf5_get_next_ijk_U0_input_indices_2_out_write),
    .input_indices_2_out1_din(tdf5_get_next_ijk_U0_input_indices_2_out1_din),
    .input_indices_2_out1_full_n(input_indices_23_c1_full_n),
    .input_indices_2_out1_write(tdf5_get_next_ijk_U0_input_indices_2_out1_write),
    .output_indices_0_din(tdf5_get_next_ijk_U0_output_indices_0_din),
    .output_indices_0_full_n(output_indices_04_c_full_n),
    .output_indices_0_write(tdf5_get_next_ijk_U0_output_indices_0_write),
    .output_indices_1_din(tdf5_get_next_ijk_U0_output_indices_1_din),
    .output_indices_1_full_n(output_indices_15_c_full_n),
    .output_indices_1_write(tdf5_get_next_ijk_U0_output_indices_1_write),
    .resetMaximum_din(tdf5_get_next_ijk_U0_resetMaximum_din),
    .resetMaximum_full_n(resetMaximum6_c_full_n),
    .resetMaximum_write(tdf5_get_next_ijk_U0_resetMaximum_write),
    .storeOutput_din(tdf5_get_next_ijk_U0_storeOutput_din),
    .storeOutput_full_n(storeOutput7_c_full_n),
    .storeOutput_write(tdf5_get_next_ijk_U0_storeOutput_write),
    .ap_return_0(tdf5_get_next_ijk_U0_ap_return_0),
    .ap_return_1(tdf5_get_next_ijk_U0_ap_return_1)
);

td_fused_top_tdf5_readInputs41 tdf5_readInputs41_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf5_readInputs41_U0_ap_start),
    .ap_done(tdf5_readInputs41_U0_ap_done),
    .ap_continue(tdf5_readInputs41_U0_ap_continue),
    .ap_idle(tdf5_readInputs41_U0_ap_idle),
    .ap_ready(tdf5_readInputs41_U0_ap_ready),
    .in_data_address0(tdf5_readInputs41_U0_in_data_address0),
    .in_data_ce0(tdf5_readInputs41_U0_in_data_ce0),
    .in_data_q0(in_data_q0),
    .i_15(input_indices_0_dout),
    .j_15(input_indices_1_dout),
    .ifmap_vec_address0(tdf5_readInputs41_U0_ifmap_vec_address0),
    .ifmap_vec_ce0(tdf5_readInputs41_U0_ifmap_vec_ce0),
    .ifmap_vec_we0(tdf5_readInputs41_U0_ifmap_vec_we0),
    .ifmap_vec_d0(tdf5_readInputs41_U0_ifmap_vec_d0),
    .ifmap_vec_address1(tdf5_readInputs41_U0_ifmap_vec_address1),
    .ifmap_vec_ce1(tdf5_readInputs41_U0_ifmap_vec_ce1),
    .ifmap_vec_we1(tdf5_readInputs41_U0_ifmap_vec_we1),
    .ifmap_vec_d1(tdf5_readInputs41_U0_ifmap_vec_d1)
);

td_fused_top_tdf5_readFilters40 tdf5_readFilters40_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf5_readFilters40_U0_ap_start),
    .ap_done(tdf5_readFilters40_U0_ap_done),
    .ap_continue(tdf5_readFilters40_U0_ap_continue),
    .ap_idle(tdf5_readFilters40_U0_ap_idle),
    .ap_ready(tdf5_readFilters40_U0_ap_ready),
    .filter_data_address0(tdf5_readFilters40_U0_filter_data_address0),
    .filter_data_ce0(tdf5_readFilters40_U0_filter_data_ce0),
    .filter_data_q0(filter_data_q0),
    .input_indices_23_dout(input_indices_23_c_dout),
    .input_indices_23_empty_n(input_indices_23_c_empty_n),
    .input_indices_23_read(tdf5_readFilters40_U0_input_indices_23_read),
    .weight_vecs_0_address0(tdf5_readFilters40_U0_weight_vecs_0_address0),
    .weight_vecs_0_ce0(tdf5_readFilters40_U0_weight_vecs_0_ce0),
    .weight_vecs_0_we0(tdf5_readFilters40_U0_weight_vecs_0_we0),
    .weight_vecs_0_d0(tdf5_readFilters40_U0_weight_vecs_0_d0)
);

td_fused_top_tdf5_dot_product tdf5_dot_product_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf5_dot_product_U0_ap_start),
    .ap_done(tdf5_dot_product_U0_ap_done),
    .ap_continue(tdf5_dot_product_U0_ap_continue),
    .ap_idle(tdf5_dot_product_U0_ap_idle),
    .ap_ready(tdf5_dot_product_U0_ap_ready),
    .ifmap_vec_address0(tdf5_dot_product_U0_ifmap_vec_address0),
    .ifmap_vec_ce0(tdf5_dot_product_U0_ifmap_vec_ce0),
    .ifmap_vec_q0(ifmap_vec_t_q0),
    .weight_vecs_0_address0(tdf5_dot_product_U0_weight_vecs_0_address0),
    .weight_vecs_0_ce0(tdf5_dot_product_U0_weight_vecs_0_ce0),
    .weight_vecs_0_q0(weight_vecs_0_t_q0),
    .products_0_address0(tdf5_dot_product_U0_products_0_address0),
    .products_0_ce0(tdf5_dot_product_U0_products_0_ce0),
    .products_0_we0(tdf5_dot_product_U0_products_0_we0),
    .products_0_d0(tdf5_dot_product_U0_products_0_d0)
);

td_fused_top_tdf5_accum_1 tdf5_accum_1_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf5_accum_1_U0_ap_start),
    .ap_done(tdf5_accum_1_U0_ap_done),
    .ap_continue(tdf5_accum_1_U0_ap_continue),
    .ap_idle(tdf5_accum_1_U0_ap_idle),
    .ap_ready(tdf5_accum_1_U0_ap_ready),
    .accum_in_0_address0(tdf5_accum_1_U0_accum_in_0_address0),
    .accum_in_0_ce0(tdf5_accum_1_U0_accum_in_0_ce0),
    .accum_in_0_q0(products_0_t_q0),
    .accum_in_0_address1(tdf5_accum_1_U0_accum_in_0_address1),
    .accum_in_0_ce1(tdf5_accum_1_U0_accum_in_0_ce1),
    .accum_in_0_q1(products_0_t_q1),
    .accum_out_address0(tdf5_accum_1_U0_accum_out_address0),
    .accum_out_ce0(tdf5_accum_1_U0_accum_out_ce0),
    .accum_out_we0(tdf5_accum_1_U0_accum_out_we0),
    .accum_out_d0(tdf5_accum_1_U0_accum_out_d0),
    .accum_out_address1(tdf5_accum_1_U0_accum_out_address1),
    .accum_out_ce1(tdf5_accum_1_U0_accum_out_ce1),
    .accum_out_we1(tdf5_accum_1_U0_accum_out_we1),
    .accum_out_d1(tdf5_accum_1_U0_accum_out_d1)
);

td_fused_top_tdf5_accum_2 tdf5_accum_2_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf5_accum_2_U0_ap_start),
    .ap_done(tdf5_accum_2_U0_ap_done),
    .ap_continue(tdf5_accum_2_U0_ap_continue),
    .ap_idle(tdf5_accum_2_U0_ap_idle),
    .ap_ready(tdf5_accum_2_U0_ap_ready),
    .accum_in_10(tdf5_accum_2_U0_accum_in_10),
    .accum_in_10_ap_vld(tdf5_accum_2_U0_accum_in_10_ap_vld),
    .accum_in_address0(tdf5_accum_2_U0_accum_in_address0),
    .accum_in_ce0(tdf5_accum_2_U0_accum_in_ce0),
    .accum_in_q0(accum1_out_0_t_q0)
);

td_fused_top_Block_entry_proc_proc408 Block_entry_proc_proc408_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(Block_entry_proc_proc408_U0_ap_start),
    .ap_done(Block_entry_proc_proc408_U0_ap_done),
    .ap_continue(Block_entry_proc_proc408_U0_ap_continue),
    .ap_idle(Block_entry_proc_proc408_U0_ap_idle),
    .ap_ready(Block_entry_proc_proc408_U0_ap_ready),
    .tmp(tmp_channel_dout),
    .ap_return(Block_entry_proc_proc408_U0_ap_return)
);

td_fused_top_tdf5_adjust tdf5_adjust_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf5_adjust_U0_ap_start),
    .ap_done(tdf5_adjust_U0_ap_done),
    .ap_continue(tdf5_adjust_U0_ap_continue),
    .ap_idle(tdf5_adjust_U0_ap_idle),
    .ap_ready(tdf5_adjust_U0_ap_ready),
    .sums_read(sums_0_dout),
    .adjustments_address0(tdf5_adjust_U0_adjustments_address0),
    .adjustments_ce0(tdf5_adjust_U0_adjustments_ce0),
    .adjustments_q0(adjustments_q0),
    .input_indices_23_dout(input_indices_23_c1_dout),
    .input_indices_23_empty_n(input_indices_23_c1_empty_n),
    .input_indices_23_read(tdf5_adjust_U0_input_indices_23_read),
    .ap_return(tdf5_adjust_U0_ap_return)
);

td_fused_top_tdf5_poolOutputs tdf5_poolOutputs_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf5_poolOutputs_U0_ap_start),
    .ap_done(tdf5_poolOutputs_U0_ap_done),
    .ap_continue(tdf5_poolOutputs_U0_ap_continue),
    .ap_idle(tdf5_poolOutputs_U0_ap_idle),
    .ap_ready(tdf5_poolOutputs_U0_ap_ready),
    .output_indices_04_dout(output_indices_04_c_dout),
    .output_indices_04_empty_n(output_indices_04_c_empty_n),
    .output_indices_04_read(tdf5_poolOutputs_U0_output_indices_04_read),
    .output_indices_15_dout(output_indices_15_c_dout),
    .output_indices_15_empty_n(output_indices_15_c_empty_n),
    .output_indices_15_read(tdf5_poolOutputs_U0_output_indices_15_read),
    .resetMaximum6_dout(resetMaximum6_c_dout),
    .resetMaximum6_empty_n(resetMaximum6_c_empty_n),
    .resetMaximum6_read(tdf5_poolOutputs_U0_resetMaximum6_read),
    .storeOutput7_dout(storeOutput7_c_dout),
    .storeOutput7_empty_n(storeOutput7_c_empty_n),
    .storeOutput7_read(tdf5_poolOutputs_U0_storeOutput7_read),
    .p_read(outputs_0_dout),
    .out_data_address1(tdf5_poolOutputs_U0_out_data_address1),
    .out_data_ce1(tdf5_poolOutputs_U0_out_data_ce1),
    .out_data_we1(tdf5_poolOutputs_U0_out_data_we1),
    .out_data_d1(tdf5_poolOutputs_U0_out_data_d1)
);

td_fused_top_fifo_w7_d2_S_x input_indices_23_c_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(input_indices_23_c_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf5_readFilters40_U0_input_indices_23_read),
    .if_dout(input_indices_23_c_dout),
    .if_full_n(input_indices_23_c_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf5_get_next_ijk_U0_input_indices_2_out_write),
    .if_din(tdf5_get_next_ijk_U0_input_indices_2_out_din)
);

td_fused_top_fifo_w7_d7_S input_indices_23_c1_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(input_indices_23_c1_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf5_adjust_U0_input_indices_23_read),
    .if_dout(input_indices_23_c1_dout),
    .if_full_n(input_indices_23_c1_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf5_get_next_ijk_U0_input_indices_2_out1_write),
    .if_din(tdf5_get_next_ijk_U0_input_indices_2_out1_din)
);

td_fused_top_fifo_w5_d8_S output_indices_04_c_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(output_indices_04_c_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf5_poolOutputs_U0_output_indices_04_read),
    .if_dout(output_indices_04_c_dout),
    .if_full_n(output_indices_04_c_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf5_get_next_ijk_U0_output_indices_0_write),
    .if_din(tdf5_get_next_ijk_U0_output_indices_0_din)
);

td_fused_top_fifo_w10_d8_S output_indices_15_c_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(output_indices_15_c_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf5_poolOutputs_U0_output_indices_15_read),
    .if_dout(output_indices_15_c_dout),
    .if_full_n(output_indices_15_c_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf5_get_next_ijk_U0_output_indices_1_write),
    .if_din(tdf5_get_next_ijk_U0_output_indices_1_din)
);

td_fused_top_fifo_w1_d8_S_x resetMaximum6_c_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(resetMaximum6_c_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf5_poolOutputs_U0_resetMaximum6_read),
    .if_dout(resetMaximum6_c_dout),
    .if_full_n(resetMaximum6_c_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf5_get_next_ijk_U0_resetMaximum_write),
    .if_din(resetMaximum6_c_din)
);

td_fused_top_fifo_w1_d8_S_x storeOutput7_c_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(storeOutput7_c_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf5_poolOutputs_U0_storeOutput7_read),
    .if_dout(storeOutput7_c_dout),
    .if_full_n(storeOutput7_c_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf5_get_next_ijk_U0_storeOutput_write),
    .if_din(storeOutput7_c_din)
);

td_fused_top_fifo_w16_d2_S_x2 input_indices_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(input_indices_0_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf5_readInputs41_U0_ap_ready),
    .if_dout(input_indices_0_dout),
    .if_full_n(input_indices_0_full_n),
    .if_write_ce(1'b1),
    .if_write(ap_channel_done_input_indices_0),
    .if_din(tdf5_get_next_ijk_U0_ap_return_0)
);

td_fused_top_fifo_w16_d2_S_x2 input_indices_1_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(input_indices_1_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf5_readInputs41_U0_ap_ready),
    .if_dout(input_indices_1_dout),
    .if_full_n(input_indices_1_full_n),
    .if_write_ce(1'b1),
    .if_write(ap_channel_done_input_indices_1),
    .if_din(tdf5_get_next_ijk_U0_ap_return_1)
);

td_fused_top_fifo_w16_d2_S_x2 tmp_channel_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(tmp_channel_empty_n),
    .if_read_ce(1'b1),
    .if_read(Block_entry_proc_proc408_U0_ap_ready),
    .if_dout(tmp_channel_dout),
    .if_full_n(tmp_channel_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf5_accum_2_U0_ap_done),
    .if_din(tdf5_accum_2_U0_accum_in_10)
);

td_fused_top_fifo_w16_d2_S_x2 sums_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(sums_0_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf5_adjust_U0_ap_ready),
    .if_dout(sums_0_dout),
    .if_full_n(sums_0_full_n),
    .if_write_ce(1'b1),
    .if_write(Block_entry_proc_proc408_U0_ap_done),
    .if_din(Block_entry_proc_proc408_U0_ap_return)
);

td_fused_top_fifo_w16_d2_S_x2 outputs_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(outputs_0_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf5_poolOutputs_U0_ap_ready),
    .if_dout(outputs_0_dout),
    .if_full_n(outputs_0_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf5_adjust_U0_ap_done),
    .if_din(tdf5_adjust_U0_ap_return)
);

td_fused_top_start_for_tdf5_readFilters40_U0 start_for_tdf5_readFilters40_U0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(start_for_tdf5_readFilters40_U0_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf5_readFilters40_U0_ap_ready),
    .if_dout(start_for_tdf5_readFilters40_U0_dout),
    .if_full_n(start_for_tdf5_readFilters40_U0_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf5_get_next_ijk_U0_start_write),
    .if_din(start_for_tdf5_readFilters40_U0_din)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_sync_reg_channel_write_input_indices_0 <= 1'b0;
    end else begin
        if (((tdf5_get_next_ijk_U0_ap_done & tdf5_get_next_ijk_U0_ap_continue) == 1'b1)) begin
            ap_sync_reg_channel_write_input_indices_0 <= 1'b0;
        end else begin
            ap_sync_reg_channel_write_input_indices_0 <= ap_sync_channel_write_input_indices_0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_sync_reg_channel_write_input_indices_1 <= 1'b0;
    end else begin
        if (((tdf5_get_next_ijk_U0_ap_done & tdf5_get_next_ijk_U0_ap_continue) == 1'b1)) begin
            ap_sync_reg_channel_write_input_indices_1 <= 1'b0;
        end else begin
            ap_sync_reg_channel_write_input_indices_1 <= ap_sync_channel_write_input_indices_1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_sync_reg_tdf5_get_next_ijk_U0_ap_ready <= 1'b0;
    end else begin
        if (((ap_sync_ready & ap_start) == 1'b1)) begin
            ap_sync_reg_tdf5_get_next_ijk_U0_ap_ready <= 1'b0;
        end else begin
            ap_sync_reg_tdf5_get_next_ijk_U0_ap_ready <= ap_sync_tdf5_get_next_ijk_U0_ap_ready;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_sync_reg_tdf5_readInputs41_U0_ap_ready <= 1'b0;
    end else begin
        if (((ap_sync_ready & ap_start) == 1'b1)) begin
            ap_sync_reg_tdf5_readInputs41_U0_ap_ready <= 1'b0;
        end else begin
            ap_sync_reg_tdf5_readInputs41_U0_ap_ready <= ap_sync_tdf5_readInputs41_U0_ap_ready;
        end
    end
end

assign Block_entry_proc_proc408_U0_ap_continue = sums_0_full_n;

assign Block_entry_proc_proc408_U0_ap_start = tmp_channel_empty_n;

assign Block_entry_proc_proc408_U0_start_full_n = 1'b1;

assign Block_entry_proc_proc408_U0_start_write = 1'b0;

assign adjustments_address0 = tdf5_adjust_U0_adjustments_address0;

assign adjustments_address1 = 7'd0;

assign adjustments_ce0 = tdf5_adjust_U0_adjustments_ce0;

assign adjustments_ce1 = 1'b0;

assign adjustments_d0 = 48'd0;

assign adjustments_d1 = 48'd0;

assign adjustments_we0 = 1'b0;

assign adjustments_we1 = 1'b0;

assign ap_channel_done_accum1_out_0 = tdf5_accum_1_U0_ap_done;

assign ap_channel_done_ifmap_vec = tdf5_readInputs41_U0_ap_done;

assign ap_channel_done_input_indices_0 = (tdf5_get_next_ijk_U0_ap_done & (ap_sync_reg_channel_write_input_indices_0 ^ 1'b1));

assign ap_channel_done_input_indices_1 = (tdf5_get_next_ijk_U0_ap_done & (ap_sync_reg_channel_write_input_indices_1 ^ 1'b1));

assign ap_channel_done_outputs_0 = tdf5_adjust_U0_ap_done;

assign ap_channel_done_products_0 = tdf5_dot_product_U0_ap_done;

assign ap_channel_done_sums_0 = Block_entry_proc_proc408_U0_ap_done;

assign ap_channel_done_tmp_channel = tdf5_accum_2_U0_ap_done;

assign ap_channel_done_weight_vecs_0 = tdf5_readFilters40_U0_ap_done;

assign ap_done = tdf5_poolOutputs_U0_ap_done;

assign ap_idle = (tdf5_readInputs41_U0_ap_idle & tdf5_readFilters40_U0_ap_idle & tdf5_poolOutputs_U0_ap_idle & tdf5_get_next_ijk_U0_ap_idle & tdf5_dot_product_U0_ap_idle & tdf5_adjust_U0_ap_idle & tdf5_accum_2_U0_ap_idle & tdf5_accum_1_U0_ap_idle & (outputs_0_empty_n ^ 1'b1) & (sums_0_empty_n ^ 1'b1) & (tmp_channel_empty_n ^ 1'b1) & (input_indices_1_empty_n ^ 1'b1) & (input_indices_0_empty_n ^ 1'b1) & (products_0_t_empty_n ^ 1'b1) & (weight_vecs_0_t_empty_n ^ 1'b1) & (ifmap_vec_t_empty_n ^ 1'b1) & (1'b1 ^ accum1_out_0_t_empty_n) & Block_entry_proc_proc408_U0_ap_idle);

assign ap_ready = ap_sync_ready;

assign ap_sync_channel_write_input_indices_0 = ((input_indices_0_full_n & ap_channel_done_input_indices_0) | ap_sync_reg_channel_write_input_indices_0);

assign ap_sync_channel_write_input_indices_1 = ((input_indices_1_full_n & ap_channel_done_input_indices_1) | ap_sync_reg_channel_write_input_indices_1);

assign ap_sync_continue = ap_continue;

assign ap_sync_done = tdf5_poolOutputs_U0_ap_done;

assign ap_sync_ready = (ap_sync_tdf5_readInputs41_U0_ap_ready & ap_sync_tdf5_get_next_ijk_U0_ap_ready);

assign ap_sync_tdf5_get_next_ijk_U0_ap_ready = (tdf5_get_next_ijk_U0_ap_ready | ap_sync_reg_tdf5_get_next_ijk_U0_ap_ready);

assign ap_sync_tdf5_readInputs41_U0_ap_ready = (tdf5_readInputs41_U0_ap_ready | ap_sync_reg_tdf5_readInputs41_U0_ap_ready);

assign filter_data_address0 = tdf5_readFilters40_U0_filter_data_address0;

assign filter_data_address1 = 15'd0;

assign filter_data_ce0 = tdf5_readFilters40_U0_filter_data_ce0;

assign filter_data_ce1 = 1'b0;

assign filter_data_d0 = 16'd0;

assign filter_data_d1 = 16'd0;

assign filter_data_we0 = 1'b0;

assign filter_data_we1 = 1'b0;

assign in_data_address0 = tdf5_readInputs41_U0_in_data_address0;

assign in_data_address1 = 14'd0;

assign in_data_ce0 = tdf5_readInputs41_U0_in_data_ce0;

assign in_data_ce1 = 1'b0;

assign in_data_d0 = 64'd0;

assign in_data_d1 = 64'd0;

assign in_data_read = tdf5_readInputs41_U0_in_data_write;

assign in_data_we0 = 1'b0;

assign in_data_we1 = 1'b0;

assign out_data_address0 = 15'd0;

assign out_data_address1 = tdf5_poolOutputs_U0_out_data_address1;

assign out_data_ce0 = 1'b0;

assign out_data_ce1 = tdf5_poolOutputs_U0_out_data_ce1;

assign out_data_d0 = 64'd0;

assign out_data_d1 = tdf5_poolOutputs_U0_out_data_d1;

assign out_data_we0 = 1'b0;

assign out_data_we1 = tdf5_poolOutputs_U0_out_data_we1;

assign out_data_write = tdf5_poolOutputs_U0_out_data_write;

assign products_0_t_d1 = 16'd0;

assign products_0_t_we1 = 1'b0;

assign resetMaximum6_c_din = tdf5_get_next_ijk_U0_resetMaximum_din;

assign start_for_tdf5_readFilters40_U0_din = 1'b1;

assign storeOutput7_c_din = tdf5_get_next_ijk_U0_storeOutput_din;

assign tdf5_accum_1_U0_accum_out_full_n = accum1_out_0_i_full_n;

assign tdf5_accum_1_U0_ap_continue = accum1_out_0_i_full_n;

assign tdf5_accum_1_U0_ap_start = products_0_t_empty_n;

assign tdf5_accum_1_U0_start_full_n = 1'b1;

assign tdf5_accum_1_U0_start_write = 1'b0;

assign tdf5_accum_2_U0_ap_continue = tmp_channel_full_n;

assign tdf5_accum_2_U0_ap_start = accum1_out_0_t_empty_n;

assign tdf5_accum_2_U0_start_full_n = 1'b1;

assign tdf5_accum_2_U0_start_write = 1'b0;

assign tdf5_adjust_U0_ap_continue = outputs_0_full_n;

assign tdf5_adjust_U0_ap_start = sums_0_empty_n;

assign tdf5_adjust_U0_start_full_n = 1'b1;

assign tdf5_adjust_U0_start_write = 1'b0;

assign tdf5_dot_product_U0_ap_continue = products_0_i_full_n;

assign tdf5_dot_product_U0_ap_start = (weight_vecs_0_t_empty_n & ifmap_vec_t_empty_n);

assign tdf5_dot_product_U0_products_0_full_n = products_0_i_full_n;

assign tdf5_dot_product_U0_start_full_n = 1'b1;

assign tdf5_dot_product_U0_start_write = 1'b0;

assign tdf5_get_next_ijk_U0_ap_continue = (ap_sync_channel_write_input_indices_1 & ap_sync_channel_write_input_indices_0);

assign tdf5_get_next_ijk_U0_ap_start = ((ap_sync_reg_tdf5_get_next_ijk_U0_ap_ready ^ 1'b1) & ap_start);

assign tdf5_poolOutputs_U0_ap_continue = ap_continue;

assign tdf5_poolOutputs_U0_ap_start = outputs_0_empty_n;

assign tdf5_poolOutputs_U0_out_data_full_n = out_data_full_n;

assign tdf5_poolOutputs_U0_out_data_write = 1'b0;

assign tdf5_poolOutputs_U0_start_full_n = 1'b1;

assign tdf5_poolOutputs_U0_start_write = 1'b0;

assign tdf5_readFilters40_U0_ap_continue = weight_vecs_0_i_full_n;

assign tdf5_readFilters40_U0_ap_start = start_for_tdf5_readFilters40_U0_empty_n;

assign tdf5_readFilters40_U0_start_full_n = 1'b1;

assign tdf5_readFilters40_U0_start_write = 1'b0;

assign tdf5_readFilters40_U0_weight_vecs_0_full_n = weight_vecs_0_i_full_n;

assign tdf5_readInputs41_U0_ap_continue = ifmap_vec_i_full_n;

assign tdf5_readInputs41_U0_ap_start = (input_indices_1_empty_n & input_indices_0_empty_n & (ap_sync_reg_tdf5_readInputs41_U0_ap_ready ^ 1'b1) & ap_start);

assign tdf5_readInputs41_U0_ifmap_vec_full_n = ifmap_vec_i_full_n;

assign tdf5_readInputs41_U0_in_data_full_n = in_data_empty_n;

assign tdf5_readInputs41_U0_in_data_write = 1'b0;

assign tdf5_readInputs41_U0_start_full_n = 1'b1;

assign tdf5_readInputs41_U0_start_write = 1'b0;

endmodule //td_fused_top_dataflow_in_loop_TOP_LOOP37738
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37738_weight_vecs_0_memcore_ram (addr0, ce0, d0, we0, q0, addr1, ce1, d1, we1, q1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 9;
parameter MEM_SIZE = 288;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
output reg[DWIDTH-1:0] q1;
input clk;

reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];




always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1) 
            ram[addr1] <= d1; 
        q1 <= ram[addr1];
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37738_weight_vecs_0_memcore(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    q0,
    address1,
    ce1,
    we1,
    d1,
    q1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd288;
parameter AddressWidth = 32'd9;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;
output[DataWidth - 1:0] q1;



td_fused_top_dataflow_in_loop_TOP_LOOP37738_weight_vecs_0_memcore_ram td_fused_top_dataflow_in_loop_TOP_LOOP37738_weight_vecs_0_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 ),
    .q1( q1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_dataflow_in_loop_TOP_LOOP37738_weight_vecs_0
#(parameter
    DataWidth    = 16,
    AddressRange = 32,
    AddressWidth = 8,
    BufferCount  = 2,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire                    i_we0,
    input  wire [AddressWidth-1:0] i_address0,
    input  wire [DataWidth-1:0]    i_d0,
    output wire [DataWidth-1:0]    i_q0,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire                    t_we0,
    input  wire [AddressWidth-1:0] t_address0,
    input  wire [DataWidth-1:0]    t_d0,
    output wire [DataWidth-1:0]    t_q0
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
wire [AddressWidth+IndexWidth-1:0]   memcore_iaddr;
wire [AddressWidth+IndexWidth-1:0]   memcore_taddr;

//------------------------Instantiation------------------
assign memcore_iaddr = {i_address0, iptr};
assign memcore_taddr = {t_address0, tptr};
td_fused_top_dataflow_in_loop_TOP_LOOP37738_weight_vecs_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP37738_weight_vecs_0_memcore_U (
    .reset    ( reset ),
    .clk      ( clk ),
    .address0 ( memcore_iaddr ),
    .ce0      ( i_ce0 ),
    .we0      ( i_we0),
    .d0       ( i_d0 ),
    .q0       ( i_q0 ),
    .address1 ( memcore_taddr ),
    .ce1      ( t_ce0 ),
    .we1      ( t_we0),
    .d1       ( t_d0 ),
    .q1       ( t_q0 )

);

//------------------------Body---------------------------

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37832_accum1_out_0_memcore_ram (addr0, ce0, d0, we0, q0, addr1, ce1, d1, we1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 3;
parameter MEM_SIZE = 8;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
input clk;

reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];




always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1) 
            ram[addr1] <= d1; 
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37832_accum1_out_0_memcore(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    q0,
    address1,
    ce1,
    we1,
    d1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd8;
parameter AddressWidth = 32'd3;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;



td_fused_top_dataflow_in_loop_TOP_LOOP37832_accum1_out_0_memcore_ram td_fused_top_dataflow_in_loop_TOP_LOOP37832_accum1_out_0_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_dataflow_in_loop_TOP_LOOP37832_accum1_out_0
#(parameter
    DataWidth    = 16,
    AddressRange = 32,
    AddressWidth = 3,
    BufferCount  = 2,
    MemLatency   = 1,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire                    i_we0,
    input  wire [AddressWidth-1:0] i_address0,
    input  wire [DataWidth-1:0]    i_d0,
    output wire [DataWidth-1:0]    i_q0,
    input  wire                    i_ce1,
    input  wire                    i_we1,
    input  wire [AddressWidth-1:0] i_address1,
    input  wire [DataWidth-1:0]    i_d1,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire                    t_we0,
    input  wire [AddressWidth-1:0] t_address0,
    input  wire [DataWidth-1:0]    t_d0,
    output wire [DataWidth-1:0]    t_q0,
    input  wire                    t_ce1,
    input  wire                    t_we1,
    input  wire [AddressWidth-1:0] t_address1,
    input  wire [DataWidth-1:0]    t_d1
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth-1:0]   prev_iptr    = 1'b0; // previous initiator index
reg  [IndexWidth-1:0]   prev_tptr    = 1'b0; // previous target index
reg  [DataWidth-1:0]    reg_q0      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid0    = 1'b0; // buffer has valid data
reg  [DataWidth-1:0]    reg_q1      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid1    = 1'b0; // buffer has valid data
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
// buffer signals
wire [BufferCount-1:0] buf_ce0;
wire [BufferCount-1:0] buf_we0;
wire [AddressWidth-1:0] buf_a0_0, buf_a0_1;
wire [DataWidth-1:0] buf_d0_0, buf_d0_1;
wire [DataWidth-1:0] buf_q0_0, buf_q0_1;
wire [BufferCount-1:0] buf_ce1;
wire [BufferCount-1:0] buf_we1;
wire [AddressWidth-1:0] buf_a1_0, buf_a1_1;
wire [DataWidth-1:0] buf_d1_0, buf_d1_1;
//------------------------Instantiation------------------
//genvar i;
        td_fused_top_dataflow_in_loop_TOP_LOOP37832_accum1_out_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP37832_accum1_out_0_memcore_U_0 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_0 ),
            .ce0      ( buf_ce0[ 0 ] ),
            .we0      ( buf_we0[ 0 ] ),
            .d0       ( buf_d0_0 ),
            .q0       ( buf_q0_0 ),
            .address1 ( buf_a1_0 ),
            .ce1      ( buf_ce1[ 0 ] ),
            .we1      ( buf_we1[ 0 ] ),
            .d1       ( buf_d1_0 )
        );
        td_fused_top_dataflow_in_loop_TOP_LOOP37832_accum1_out_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP37832_accum1_out_0_memcore_U_1 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_1 ),
            .ce0      ( buf_ce0[ 1 ] ),
            .we0      ( buf_we0[ 1 ] ),
            .d0       ( buf_d0_1 ),
            .q0       ( buf_q0_1 ),
            .address1 ( buf_a1_1 ),
            .ce1      ( buf_ce1[ 1 ] ),
            .we1      ( buf_we1[ 1 ] ),
            .d1       ( buf_d1_1 )
        );

//++++++++++++++++++++++++buffer signals+++++++++++++++++
        assign buf_ce0[ 0 ] = (tptr ==  0  && empty_n) ? t_ce0
                             : (iptr ==  0 ) ? i_ce0 : 1'b0;
        assign buf_a0_0  = (tptr ==  0  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 0 ] = (tptr ==  0  && empty_n)  ? t_we0
                             : (iptr ==  0 ) ? i_we0 : 1'b0;
        assign buf_d0_0  = (tptr ==  0  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 0 ] = (tptr ==  0  && empty_n) ? t_ce1
                             : (iptr ==  0 ) ? i_ce1 : 1'b0;
        assign buf_a1_0  = (tptr ==  0  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 0 ] = (tptr ==  0  && empty_n)  ? t_we1
                             : (iptr ==  0 ) ? i_we1 : 1'b0;
        assign buf_d1_0  = (tptr ==  0  && empty_n) ? t_d1       : i_d1;
        assign buf_ce0[ 1 ] = (tptr ==  1  && empty_n) ? t_ce0
                             : (iptr ==  1 ) ? i_ce0 : 1'b0;
        assign buf_a0_1  = (tptr ==  1  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 1 ] = (tptr ==  1  && empty_n)  ? t_we0
                             : (iptr ==  1 ) ? i_we0 : 1'b0;
        assign buf_d0_1  = (tptr ==  1  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 1 ] = (tptr ==  1  && empty_n) ? t_ce1
                             : (iptr ==  1 ) ? i_ce1 : 1'b0;
        assign buf_a1_1  = (tptr ==  1  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 1 ] = (tptr ==  1  && empty_n)  ? t_we1
                             : (iptr ==  1 ) ? i_we1 : 1'b0;
        assign buf_d1_1  = (tptr ==  1  && empty_n) ? t_d1       : i_d1;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//------------------------Body---------------------------
assign i_q0      = (prev_iptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign t_q0      = reg_valid0 ? reg_q0 : (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// prev_iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_iptr <= 1'b0;
    else begin
        prev_iptr <= iptr;
    end
end

// prev_tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_tptr <= 1'b0;
    else begin
        prev_tptr <= tptr;
    end
end

// reg_q0 and reg_valid0
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q0     <= 1'b0;
        reg_valid0 <= 1'b0;
    end else if (!t_ce0 && !reg_valid0) begin
        reg_q0     <= (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
        reg_valid0 <= 1'b1;
    end else if (t_ce0) begin
        reg_valid0 <= 1'b0;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37832_ifmap_vec_memcore_ram (addr0, ce0, d0, we0, q0, addr1, ce1, d1, we1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 8;
parameter MEM_SIZE = 144;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
input clk;

reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];




always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1) 
            ram[addr1] <= d1; 
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37832_ifmap_vec_memcore(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    q0,
    address1,
    ce1,
    we1,
    d1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd144;
parameter AddressWidth = 32'd8;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;



td_fused_top_dataflow_in_loop_TOP_LOOP37832_ifmap_vec_memcore_ram td_fused_top_dataflow_in_loop_TOP_LOOP37832_ifmap_vec_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_dataflow_in_loop_TOP_LOOP37832_ifmap_vec
#(parameter
    DataWidth    = 16,
    AddressRange = 32,
    AddressWidth = 8,
    BufferCount  = 2,
    MemLatency   = 1,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire                    i_we0,
    input  wire [AddressWidth-1:0] i_address0,
    input  wire [DataWidth-1:0]    i_d0,
    output wire [DataWidth-1:0]    i_q0,
    input  wire                    i_ce1,
    input  wire                    i_we1,
    input  wire [AddressWidth-1:0] i_address1,
    input  wire [DataWidth-1:0]    i_d1,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire                    t_we0,
    input  wire [AddressWidth-1:0] t_address0,
    input  wire [DataWidth-1:0]    t_d0,
    output wire [DataWidth-1:0]    t_q0,
    input  wire                    t_ce1,
    input  wire                    t_we1,
    input  wire [AddressWidth-1:0] t_address1,
    input  wire [DataWidth-1:0]    t_d1
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth-1:0]   prev_iptr    = 1'b0; // previous initiator index
reg  [IndexWidth-1:0]   prev_tptr    = 1'b0; // previous target index
reg  [DataWidth-1:0]    reg_q0      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid0    = 1'b0; // buffer has valid data
reg  [DataWidth-1:0]    reg_q1      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid1    = 1'b0; // buffer has valid data
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
// buffer signals
wire [BufferCount-1:0] buf_ce0;
wire [BufferCount-1:0] buf_we0;
wire [AddressWidth-1:0] buf_a0_0, buf_a0_1;
wire [DataWidth-1:0] buf_d0_0, buf_d0_1;
wire [DataWidth-1:0] buf_q0_0, buf_q0_1;
wire [BufferCount-1:0] buf_ce1;
wire [BufferCount-1:0] buf_we1;
wire [AddressWidth-1:0] buf_a1_0, buf_a1_1;
wire [DataWidth-1:0] buf_d1_0, buf_d1_1;
//------------------------Instantiation------------------
//genvar i;
        td_fused_top_dataflow_in_loop_TOP_LOOP37832_ifmap_vec_memcore td_fused_top_dataflow_in_loop_TOP_LOOP37832_ifmap_vec_memcore_U_0 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_0 ),
            .ce0      ( buf_ce0[ 0 ] ),
            .we0      ( buf_we0[ 0 ] ),
            .d0       ( buf_d0_0 ),
            .q0       ( buf_q0_0 ),
            .address1 ( buf_a1_0 ),
            .ce1      ( buf_ce1[ 0 ] ),
            .we1      ( buf_we1[ 0 ] ),
            .d1       ( buf_d1_0 )
        );
        td_fused_top_dataflow_in_loop_TOP_LOOP37832_ifmap_vec_memcore td_fused_top_dataflow_in_loop_TOP_LOOP37832_ifmap_vec_memcore_U_1 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_1 ),
            .ce0      ( buf_ce0[ 1 ] ),
            .we0      ( buf_we0[ 1 ] ),
            .d0       ( buf_d0_1 ),
            .q0       ( buf_q0_1 ),
            .address1 ( buf_a1_1 ),
            .ce1      ( buf_ce1[ 1 ] ),
            .we1      ( buf_we1[ 1 ] ),
            .d1       ( buf_d1_1 )
        );

//++++++++++++++++++++++++buffer signals+++++++++++++++++
        assign buf_ce0[ 0 ] = (tptr ==  0  && empty_n) ? t_ce0
                             : (iptr ==  0 ) ? i_ce0 : 1'b0;
        assign buf_a0_0  = (tptr ==  0  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 0 ] = (tptr ==  0  && empty_n)  ? t_we0
                             : (iptr ==  0 ) ? i_we0 : 1'b0;
        assign buf_d0_0  = (tptr ==  0  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 0 ] = (tptr ==  0  && empty_n) ? t_ce1
                             : (iptr ==  0 ) ? i_ce1 : 1'b0;
        assign buf_a1_0  = (tptr ==  0  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 0 ] = (tptr ==  0  && empty_n)  ? t_we1
                             : (iptr ==  0 ) ? i_we1 : 1'b0;
        assign buf_d1_0  = (tptr ==  0  && empty_n) ? t_d1       : i_d1;
        assign buf_ce0[ 1 ] = (tptr ==  1  && empty_n) ? t_ce0
                             : (iptr ==  1 ) ? i_ce0 : 1'b0;
        assign buf_a0_1  = (tptr ==  1  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 1 ] = (tptr ==  1  && empty_n)  ? t_we0
                             : (iptr ==  1 ) ? i_we0 : 1'b0;
        assign buf_d0_1  = (tptr ==  1  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 1 ] = (tptr ==  1  && empty_n) ? t_ce1
                             : (iptr ==  1 ) ? i_ce1 : 1'b0;
        assign buf_a1_1  = (tptr ==  1  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 1 ] = (tptr ==  1  && empty_n)  ? t_we1
                             : (iptr ==  1 ) ? i_we1 : 1'b0;
        assign buf_d1_1  = (tptr ==  1  && empty_n) ? t_d1       : i_d1;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//------------------------Body---------------------------
assign i_q0      = (prev_iptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign t_q0      = reg_valid0 ? reg_q0 : (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// prev_iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_iptr <= 1'b0;
    else begin
        prev_iptr <= iptr;
    end
end

// prev_tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_tptr <= 1'b0;
    else begin
        prev_tptr <= tptr;
    end
end

// reg_q0 and reg_valid0
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q0     <= 1'b0;
        reg_valid0 <= 1'b0;
    end else if (!t_ce0 && !reg_valid0) begin
        reg_q0     <= (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
        reg_valid0 <= 1'b1;
    end else if (t_ce0) begin
        reg_valid0 <= 1'b0;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37832_l2_products_memcore_ram (addr0, ce0, d0, we0, q0, addr1, ce1, d1, we1, q1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 5;
parameter MEM_SIZE = 32;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
output reg[DWIDTH-1:0] q1;
input clk;

 reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];




always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1) 
            ram[addr1] <= d1; 
        q1 <= ram[addr1];
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37832_l2_products_memcore(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    q0,
    address1,
    ce1,
    we1,
    d1,
    q1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd32;
parameter AddressWidth = 32'd5;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;
output[DataWidth - 1:0] q1;



td_fused_top_dataflow_in_loop_TOP_LOOP37832_l2_products_memcore_ram td_fused_top_dataflow_in_loop_TOP_LOOP37832_l2_products_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 ),
    .q1( q1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_dataflow_in_loop_TOP_LOOP37832_l2_products
#(parameter
    DataWidth    = 16,
    AddressRange = 32,
    AddressWidth = 4,
    BufferCount  = 2,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire                    i_we0,
    input  wire [AddressWidth-1:0] i_address0,
    input  wire [DataWidth-1:0]    i_d0,
    output wire [DataWidth-1:0]    i_q0,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire                    t_we0,
    input  wire [AddressWidth-1:0] t_address0,
    input  wire [DataWidth-1:0]    t_d0,
    output wire [DataWidth-1:0]    t_q0
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
wire [AddressWidth+IndexWidth-1:0]   memcore_iaddr;
wire [AddressWidth+IndexWidth-1:0]   memcore_taddr;

//------------------------Instantiation------------------
assign memcore_iaddr = {i_address0, iptr};
assign memcore_taddr = {t_address0, tptr};
td_fused_top_dataflow_in_loop_TOP_LOOP37832_l2_products_memcore td_fused_top_dataflow_in_loop_TOP_LOOP37832_l2_products_memcore_U (
    .reset    ( reset ),
    .clk      ( clk ),
    .address0 ( memcore_iaddr ),
    .ce0      ( i_ce0 ),
    .we0      ( i_we0),
    .d0       ( i_d0 ),
    .q0       ( i_q0 ),
    .address1 ( memcore_taddr ),
    .ce1      ( t_ce0 ),
    .we1      ( t_we0),
    .d1       ( t_d0 ),
    .q1       ( t_q0 )

);

//------------------------Body---------------------------

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37832_products_0_memcore_ram (addr0, ce0, d0, we0, q0, addr1, ce1, q1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 8;
parameter MEM_SIZE = 144;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
output reg[DWIDTH-1:0] q1;
input clk;

reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];




always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        q1 <= ram[addr1];
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37832_products_0_memcore(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    q0,
    address1,
    ce1,
    q1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd144;
parameter AddressWidth = 32'd8;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
output[DataWidth - 1:0] q1;



td_fused_top_dataflow_in_loop_TOP_LOOP37832_products_0_memcore_ram td_fused_top_dataflow_in_loop_TOP_LOOP37832_products_0_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .q1( q1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_dataflow_in_loop_TOP_LOOP37832_products_0
#(parameter
    DataWidth    = 16,
    AddressRange = 32,
    AddressWidth = 8,
    BufferCount  = 2,
    MemLatency   = 1,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire                    i_we0,
    input  wire [AddressWidth-1:0] i_address0,
    input  wire [DataWidth-1:0]    i_d0,
    output wire [DataWidth-1:0]    i_q0,
    input  wire                    i_ce1,
    input  wire [AddressWidth-1:0] i_address1,
    output wire [DataWidth-1:0]    i_q1,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire                    t_we0,
    input  wire [AddressWidth-1:0] t_address0,
    input  wire [DataWidth-1:0]    t_d0,
    output wire [DataWidth-1:0]    t_q0,
    input  wire                    t_ce1,
    input  wire [AddressWidth-1:0] t_address1,
    output wire [DataWidth-1:0]    t_q1
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth-1:0]   prev_iptr    = 1'b0; // previous initiator index
reg  [IndexWidth-1:0]   prev_tptr    = 1'b0; // previous target index
reg  [DataWidth-1:0]    reg_q0      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid0    = 1'b0; // buffer has valid data
reg  [DataWidth-1:0]    reg_q1      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid1    = 1'b0; // buffer has valid data
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
// buffer signals
wire [BufferCount-1:0] buf_ce0;
wire [BufferCount-1:0] buf_we0;
wire [AddressWidth-1:0] buf_a0_0, buf_a0_1;
wire [DataWidth-1:0] buf_d0_0, buf_d0_1;
wire [DataWidth-1:0] buf_q0_0, buf_q0_1;
wire [BufferCount-1:0] buf_ce1;
wire [AddressWidth-1:0] buf_a1_0, buf_a1_1;
wire [DataWidth-1:0] buf_q1_0, buf_q1_1;
//------------------------Instantiation------------------
//genvar i;
        td_fused_top_dataflow_in_loop_TOP_LOOP37832_products_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP37832_products_0_memcore_U_0 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_0 ),
            .ce0      ( buf_ce0[ 0 ] ),
            .we0      ( buf_we0[ 0 ] ),
            .d0       ( buf_d0_0 ),
            .q0       ( buf_q0_0 ),
            .address1 ( buf_a1_0 ),
            .ce1      ( buf_ce1[ 0 ] ),
            .q1       ( buf_q1_0 )
        );
        td_fused_top_dataflow_in_loop_TOP_LOOP37832_products_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP37832_products_0_memcore_U_1 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_1 ),
            .ce0      ( buf_ce0[ 1 ] ),
            .we0      ( buf_we0[ 1 ] ),
            .d0       ( buf_d0_1 ),
            .q0       ( buf_q0_1 ),
            .address1 ( buf_a1_1 ),
            .ce1      ( buf_ce1[ 1 ] ),
            .q1       ( buf_q1_1 )
        );

//++++++++++++++++++++++++buffer signals+++++++++++++++++
        assign buf_ce0[ 0 ] = (tptr ==  0  && empty_n) ? t_ce0
                             : (iptr ==  0 ) ? i_ce0 : 1'b0;
        assign buf_a0_0  = (tptr ==  0  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 0 ] = (tptr ==  0  && empty_n)  ? t_we0
                             : (iptr ==  0 ) ? i_we0 : 1'b0;
        assign buf_d0_0  = (tptr ==  0  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 0 ] = (tptr ==  0  && empty_n) ? t_ce1
                             : (iptr ==  0 ) ? i_ce1 : 1'b0;
        assign buf_a1_0  = (tptr ==  0  && empty_n) ?  t_address1 : i_address1;
        assign buf_ce0[ 1 ] = (tptr ==  1  && empty_n) ? t_ce0
                             : (iptr ==  1 ) ? i_ce0 : 1'b0;
        assign buf_a0_1  = (tptr ==  1  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 1 ] = (tptr ==  1  && empty_n)  ? t_we0
                             : (iptr ==  1 ) ? i_we0 : 1'b0;
        assign buf_d0_1  = (tptr ==  1  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 1 ] = (tptr ==  1  && empty_n) ? t_ce1
                             : (iptr ==  1 ) ? i_ce1 : 1'b0;
        assign buf_a1_1  = (tptr ==  1  && empty_n) ?  t_address1 : i_address1;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//------------------------Body---------------------------
assign i_q0      = (prev_iptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign t_q0      = reg_valid0 ? reg_q0 : (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign i_q1      = (prev_iptr == 1'b1 ? buf_q1_1 : buf_q1_0);
assign t_q1      = reg_valid1 ? reg_q1 : (prev_tptr == 1'b1 ? buf_q1_1 : buf_q1_0);

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// prev_iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_iptr <= 1'b0;
    else begin
        prev_iptr <= iptr;
    end
end

// prev_tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_tptr <= 1'b0;
    else begin
        prev_tptr <= tptr;
    end
end

// reg_q0 and reg_valid0
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q0     <= 1'b0;
        reg_valid0 <= 1'b0;
    end else if (!t_ce0 && !reg_valid0) begin
        reg_q0     <= (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
        reg_valid0 <= 1'b1;
    end else if (t_ce0) begin
        reg_valid0 <= 1'b0;
    end
end

// reg_q1 and reg_valid1
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q1     <= 1'b0;
        reg_valid1 <= 1'b0;
    end else if (!t_ce1 && !reg_valid1) begin
        reg_q1     <= (prev_tptr == 1'b1 ? buf_q1_1 : buf_q1_0);
        reg_valid1 <= 1'b1;
    end else if (t_ce1) begin
        reg_valid1 <= 1'b0;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_dataflow_in_loop_TOP_LOOP37832 (
        ap_clk,
        ap_rst,
        in_data_address0,
        in_data_ce0,
        in_data_d0,
        in_data_q0,
        in_data_we0,
        in_data_address1,
        in_data_ce1,
        in_data_d1,
        in_data_q1,
        in_data_we1,
        l1_filter_data_address0,
        l1_filter_data_ce0,
        l1_filter_data_d0,
        l1_filter_data_q0,
        l1_filter_data_we0,
        l1_filter_data_address1,
        l1_filter_data_ce1,
        l1_filter_data_d1,
        l1_filter_data_q1,
        l1_filter_data_we1,
        l1_adjustments_address0,
        l1_adjustments_ce0,
        l1_adjustments_d0,
        l1_adjustments_q0,
        l1_adjustments_we0,
        l1_adjustments_address1,
        l1_adjustments_ce1,
        l1_adjustments_d1,
        l1_adjustments_q1,
        l1_adjustments_we1,
        l2_filter_data_address0,
        l2_filter_data_ce0,
        l2_filter_data_d0,
        l2_filter_data_q0,
        l2_filter_data_we0,
        l2_filter_data_address1,
        l2_filter_data_ce1,
        l2_filter_data_d1,
        l2_filter_data_q1,
        l2_filter_data_we1,
        out_data_address0,
        out_data_ce0,
        out_data_d0,
        out_data_q0,
        out_data_we0,
        out_data_address1,
        out_data_ce1,
        out_data_d1,
        out_data_q1,
        out_data_we1,
        l2_adjustments_address0,
        l2_adjustments_ce0,
        l2_adjustments_d0,
        l2_adjustments_q0,
        l2_adjustments_we0,
        l2_adjustments_address1,
        l2_adjustments_ce1,
        l2_adjustments_d1,
        l2_adjustments_q1,
        l2_adjustments_we1,
        ap_start,
        in_data_empty_n,
        in_data_read,
        out_data_full_n,
        out_data_write,
        ap_done,
        ap_ready,
        ap_idle,
        ap_continue
);


input   ap_clk;
input   ap_rst;
output  [13:0] in_data_address0;
output   in_data_ce0;
output  [63:0] in_data_d0;
input  [63:0] in_data_q0;
output   in_data_we0;
output  [13:0] in_data_address1;
output   in_data_ce1;
output  [63:0] in_data_d1;
input  [63:0] in_data_q1;
output   in_data_we1;
output  [14:0] l1_filter_data_address0;
output   l1_filter_data_ce0;
output  [15:0] l1_filter_data_d0;
input  [15:0] l1_filter_data_q0;
output   l1_filter_data_we0;
output  [14:0] l1_filter_data_address1;
output   l1_filter_data_ce1;
output  [15:0] l1_filter_data_d1;
input  [15:0] l1_filter_data_q1;
output   l1_filter_data_we1;
output  [6:0] l1_adjustments_address0;
output   l1_adjustments_ce0;
output  [47:0] l1_adjustments_d0;
input  [47:0] l1_adjustments_q0;
output   l1_adjustments_we0;
output  [6:0] l1_adjustments_address1;
output   l1_adjustments_ce1;
output  [47:0] l1_adjustments_d1;
input  [47:0] l1_adjustments_q1;
output   l1_adjustments_we1;
output  [10:0] l2_filter_data_address0;
output   l2_filter_data_ce0;
output  [15:0] l2_filter_data_d0;
input  [15:0] l2_filter_data_q0;
output   l2_filter_data_we0;
output  [10:0] l2_filter_data_address1;
output   l2_filter_data_ce1;
output  [15:0] l2_filter_data_d1;
input  [15:0] l2_filter_data_q1;
output   l2_filter_data_we1;
output  [13:0] out_data_address0;
output   out_data_ce0;
output  [63:0] out_data_d0;
input  [63:0] out_data_q0;
output   out_data_we0;
output  [13:0] out_data_address1;
output   out_data_ce1;
output  [63:0] out_data_d1;
input  [63:0] out_data_q1;
output   out_data_we1;
output  [3:0] l2_adjustments_address0;
output   l2_adjustments_ce0;
output  [47:0] l2_adjustments_d0;
input  [47:0] l2_adjustments_q0;
output   l2_adjustments_we0;
output  [3:0] l2_adjustments_address1;
output   l2_adjustments_ce1;
output  [47:0] l2_adjustments_d1;
input  [47:0] l2_adjustments_q1;
output   l2_adjustments_we1;
input   ap_start;
input   in_data_empty_n;
output   in_data_read;
input   out_data_full_n;
output   out_data_write;
output   ap_done;
output   ap_ready;
output   ap_idle;
input   ap_continue;

wire   [15:0] ifmap_vec_i_q0;
wire   [15:0] ifmap_vec_t_q0;
wire   [15:0] weight_vecs_0_i_q0;
wire   [15:0] weight_vecs_0_t_q0;
wire   [15:0] products_0_i_q0;
wire   [15:0] products_0_i_q1;
wire   [15:0] products_0_t_q0;
wire   [15:0] products_0_t_q1;
wire   [15:0] accum1_out_0_i_q0;
wire   [15:0] accum1_out_0_t_q0;
wire   [15:0] l2_products_i_q0;
wire   [15:0] l2_products_t_q0;
wire    tdf4_get_next_ijk_U0_ap_start;
wire    tdf4_get_next_ijk_U0_ap_done;
wire    tdf4_get_next_ijk_U0_ap_continue;
wire    tdf4_get_next_ijk_U0_ap_idle;
wire    tdf4_get_next_ijk_U0_ap_ready;
wire    tdf4_get_next_ijk_U0_start_out;
wire    tdf4_get_next_ijk_U0_start_write;
wire   [15:0] tdf4_get_next_ijk_U0_indices_0_din;
wire    tdf4_get_next_ijk_U0_indices_0_write;
wire   [15:0] tdf4_get_next_ijk_U0_indices_1_din;
wire    tdf4_get_next_ijk_U0_indices_1_write;
wire   [6:0] tdf4_get_next_ijk_U0_indices_2_out_din;
wire    tdf4_get_next_ijk_U0_indices_2_out_write;
wire   [10:0] tdf4_get_next_ijk_U0_indices_2_out1_din;
wire    tdf4_get_next_ijk_U0_indices_2_out1_write;
wire    tdf4_get_next_ijk_U0_write_r_din;
wire    tdf4_get_next_ijk_U0_write_r_write;
wire    tdf4_readInputs37_U0_ap_start;
wire    tdf4_readInputs37_U0_ap_done;
wire    tdf4_readInputs37_U0_ap_continue;
wire    tdf4_readInputs37_U0_ap_idle;
wire    tdf4_readInputs37_U0_ap_ready;
wire   [13:0] tdf4_readInputs37_U0_in_data_address0;
wire    tdf4_readInputs37_U0_in_data_ce0;
wire    tdf4_readInputs37_U0_indices_01_read;
wire    tdf4_readInputs37_U0_indices_12_read;
wire   [7:0] tdf4_readInputs37_U0_ifmap_vec_address0;
wire    tdf4_readInputs37_U0_ifmap_vec_ce0;
wire    tdf4_readInputs37_U0_ifmap_vec_we0;
wire   [15:0] tdf4_readInputs37_U0_ifmap_vec_d0;
wire   [7:0] tdf4_readInputs37_U0_ifmap_vec_address1;
wire    tdf4_readInputs37_U0_ifmap_vec_ce1;
wire    tdf4_readInputs37_U0_ifmap_vec_we1;
wire   [15:0] tdf4_readInputs37_U0_ifmap_vec_d1;
wire   [5:0] tdf4_readInputs37_U0_indices_01_out_din;
wire    tdf4_readInputs37_U0_indices_01_out_write;
wire   [11:0] tdf4_readInputs37_U0_indices_12_out_din;
wire    tdf4_readInputs37_U0_indices_12_out_write;
wire    tdf4_readInputs37_U0_in_data_full_n;
wire    tdf4_readInputs37_U0_in_data_write;
wire    ap_channel_done_ifmap_vec;
wire    tdf4_readInputs37_U0_ifmap_vec_full_n;
wire    tdf4_readFilters36_U0_ap_start;
wire    tdf4_readFilters36_U0_ap_done;
wire    tdf4_readFilters36_U0_ap_continue;
wire    tdf4_readFilters36_U0_ap_idle;
wire    tdf4_readFilters36_U0_ap_ready;
wire   [14:0] tdf4_readFilters36_U0_filter_data_address0;
wire    tdf4_readFilters36_U0_filter_data_ce0;
wire    tdf4_readFilters36_U0_indices_23_read;
wire   [7:0] tdf4_readFilters36_U0_weight_vecs_0_address0;
wire    tdf4_readFilters36_U0_weight_vecs_0_ce0;
wire    tdf4_readFilters36_U0_weight_vecs_0_we0;
wire   [15:0] tdf4_readFilters36_U0_weight_vecs_0_d0;
wire    ap_channel_done_weight_vecs_0;
wire    tdf4_readFilters36_U0_weight_vecs_0_full_n;
wire    tdf4_dot_product_U0_ap_start;
wire    tdf4_dot_product_U0_ap_done;
wire    tdf4_dot_product_U0_ap_continue;
wire    tdf4_dot_product_U0_ap_idle;
wire    tdf4_dot_product_U0_ap_ready;
wire   [7:0] tdf4_dot_product_U0_ifmap_vec_address0;
wire    tdf4_dot_product_U0_ifmap_vec_ce0;
wire   [7:0] tdf4_dot_product_U0_weight_vecs_0_address0;
wire    tdf4_dot_product_U0_weight_vecs_0_ce0;
wire   [7:0] tdf4_dot_product_U0_products_0_address0;
wire    tdf4_dot_product_U0_products_0_ce0;
wire    tdf4_dot_product_U0_products_0_we0;
wire   [15:0] tdf4_dot_product_U0_products_0_d0;
wire    ap_channel_done_products_0;
wire    tdf4_dot_product_U0_products_0_full_n;
wire    tdf4_accum_1_U0_ap_start;
wire    tdf4_accum_1_U0_ap_done;
wire    tdf4_accum_1_U0_ap_continue;
wire    tdf4_accum_1_U0_ap_idle;
wire    tdf4_accum_1_U0_ap_ready;
wire   [7:0] tdf4_accum_1_U0_accum_in_0_address0;
wire    tdf4_accum_1_U0_accum_in_0_ce0;
wire   [7:0] tdf4_accum_1_U0_accum_in_0_address1;
wire    tdf4_accum_1_U0_accum_in_0_ce1;
wire   [2:0] tdf4_accum_1_U0_accum_out_address0;
wire    tdf4_accum_1_U0_accum_out_ce0;
wire    tdf4_accum_1_U0_accum_out_we0;
wire   [15:0] tdf4_accum_1_U0_accum_out_d0;
wire   [2:0] tdf4_accum_1_U0_accum_out_address1;
wire    tdf4_accum_1_U0_accum_out_ce1;
wire    tdf4_accum_1_U0_accum_out_we1;
wire   [15:0] tdf4_accum_1_U0_accum_out_d1;
wire    ap_channel_done_accum1_out_0;
wire    tdf4_accum_1_U0_accum_out_full_n;
wire    tdf4_accum_2_U0_ap_start;
wire    tdf4_accum_2_U0_ap_done;
wire    tdf4_accum_2_U0_ap_continue;
wire    tdf4_accum_2_U0_ap_idle;
wire    tdf4_accum_2_U0_ap_ready;
wire   [15:0] tdf4_accum_2_U0_accum_in_12;
wire    tdf4_accum_2_U0_accum_in_12_ap_vld;
wire   [2:0] tdf4_accum_2_U0_accum_in_address0;
wire    tdf4_accum_2_U0_accum_in_ce0;
wire    ap_channel_done_tmp_channel;
wire    tmp_channel_full_n;
wire    Block_entry_proc_proc403_U0_ap_start;
wire    Block_entry_proc_proc403_U0_ap_done;
wire    Block_entry_proc_proc403_U0_ap_continue;
wire    Block_entry_proc_proc403_U0_ap_idle;
wire    Block_entry_proc_proc403_U0_ap_ready;
wire   [15:0] Block_entry_proc_proc403_U0_ap_return;
wire    ap_channel_done_sums_0;
wire    sums_0_full_n;
wire    tdf4_adjust_U0_ap_start;
wire    tdf4_adjust_U0_ap_done;
wire    tdf4_adjust_U0_ap_continue;
wire    tdf4_adjust_U0_ap_idle;
wire    tdf4_adjust_U0_ap_ready;
wire   [6:0] tdf4_adjust_U0_adjustments_address0;
wire    tdf4_adjust_U0_adjustments_ce0;
wire    tdf4_adjust_U0_indices_23_read;
wire   [10:0] tdf4_adjust_U0_indices_23_out_din;
wire    tdf4_adjust_U0_indices_23_out_write;
wire   [15:0] tdf4_adjust_U0_ap_return;
wire    ap_channel_done_intermediate_fmaps_0;
wire    intermediate_fmaps_0_full_n;
wire    tdf4_l2_multiply34_U0_ap_start;
wire    tdf4_l2_multiply34_U0_ap_done;
wire    tdf4_l2_multiply34_U0_ap_continue;
wire    tdf4_l2_multiply34_U0_ap_idle;
wire    tdf4_l2_multiply34_U0_ap_ready;
wire   [10:0] tdf4_l2_multiply34_U0_l2_filter_data_address0;
wire    tdf4_l2_multiply34_U0_l2_filter_data_ce0;
wire   [3:0] tdf4_l2_multiply34_U0_l2_products_address0;
wire    tdf4_l2_multiply34_U0_l2_products_ce0;
wire    tdf4_l2_multiply34_U0_l2_products_we0;
wire   [15:0] tdf4_l2_multiply34_U0_l2_products_d0;
wire    tdf4_l2_multiply34_U0_indices_23_read;
wire    ap_channel_done_l2_products;
wire    tdf4_l2_multiply34_U0_l2_products_full_n;
wire    tdf4_l2_writeOutputs_133_U0_ap_start;
wire    tdf4_l2_writeOutputs_133_U0_ap_done;
wire    tdf4_l2_writeOutputs_133_U0_ap_continue;
wire    tdf4_l2_writeOutputs_133_U0_ap_idle;
wire    tdf4_l2_writeOutputs_133_U0_ap_ready;
wire    tdf4_l2_writeOutputs_133_U0_indices_01_read;
wire    tdf4_l2_writeOutputs_133_U0_indices_12_read;
wire    tdf4_l2_writeOutputs_133_U0_write4_read;
wire   [3:0] tdf4_l2_writeOutputs_133_U0_l2_partial_sums_address0;
wire    tdf4_l2_writeOutputs_133_U0_l2_partial_sums_ce0;
wire   [13:0] tdf4_l2_writeOutputs_133_U0_out_data_address1;
wire    tdf4_l2_writeOutputs_133_U0_out_data_ce1;
wire    tdf4_l2_writeOutputs_133_U0_out_data_we1;
wire   [63:0] tdf4_l2_writeOutputs_133_U0_out_data_d1;
wire   [3:0] tdf4_l2_writeOutputs_133_U0_l2_adjustments_address0;
wire    tdf4_l2_writeOutputs_133_U0_l2_adjustments_ce0;
wire    tdf4_l2_writeOutputs_133_U0_out_data_full_n;
wire    tdf4_l2_writeOutputs_133_U0_out_data_write;
wire    ap_sync_continue;
wire    ifmap_vec_i_full_n;
wire    ifmap_vec_t_empty_n;
wire    weight_vecs_0_i_full_n;
wire    weight_vecs_0_t_empty_n;
wire    products_0_i_full_n;
wire    products_0_t_empty_n;
wire   [15:0] products_0_t_d1;
wire    products_0_t_we1;
wire    accum1_out_0_i_full_n;
wire    accum1_out_0_t_empty_n;
wire    l2_products_i_full_n;
wire    l2_products_t_empty_n;
wire    indices_01_c_full_n;
wire   [15:0] indices_01_c_dout;
wire    indices_01_c_empty_n;
wire    indices_12_c_full_n;
wire   [15:0] indices_12_c_dout;
wire    indices_12_c_empty_n;
wire    indices_23_c_full_n;
wire   [6:0] indices_23_c_dout;
wire    indices_23_c_empty_n;
wire    indices_23_c1_full_n;
wire   [10:0] indices_23_c1_dout;
wire    indices_23_c1_empty_n;
wire   [0:0] write4_c_din;
wire    write4_c_full_n;
wire   [0:0] write4_c_dout;
wire    write4_c_empty_n;
wire    indices_01_c2_full_n;
wire   [5:0] indices_01_c2_dout;
wire    indices_01_c2_empty_n;
wire    indices_12_c3_full_n;
wire   [11:0] indices_12_c3_dout;
wire    indices_12_c3_empty_n;
wire   [15:0] tmp_channel_dout;
wire    tmp_channel_empty_n;
wire   [15:0] sums_0_dout;
wire    sums_0_empty_n;
wire    indices_23_c4_full_n;
wire   [10:0] indices_23_c4_dout;
wire    indices_23_c4_empty_n;
wire   [15:0] intermediate_fmaps_0_dout;
wire    intermediate_fmaps_0_empty_n;
wire    ap_sync_done;
wire    ap_sync_ready;
reg    ap_sync_reg_tdf4_get_next_ijk_U0_ap_ready;
wire    ap_sync_tdf4_get_next_ijk_U0_ap_ready;
reg    ap_sync_reg_tdf4_readInputs37_U0_ap_ready;
wire    ap_sync_tdf4_readInputs37_U0_ap_ready;
wire   [0:0] start_for_tdf4_readFilters36_U0_din;
wire    start_for_tdf4_readFilters36_U0_full_n;
wire   [0:0] start_for_tdf4_readFilters36_U0_dout;
wire    start_for_tdf4_readFilters36_U0_empty_n;
wire    tdf4_readInputs37_U0_start_full_n;
wire    tdf4_readInputs37_U0_start_write;
wire    tdf4_readFilters36_U0_start_full_n;
wire    tdf4_readFilters36_U0_start_write;
wire    tdf4_dot_product_U0_start_full_n;
wire    tdf4_dot_product_U0_start_write;
wire    tdf4_accum_1_U0_start_full_n;
wire    tdf4_accum_1_U0_start_write;
wire    tdf4_accum_2_U0_start_full_n;
wire    tdf4_accum_2_U0_start_write;
wire    Block_entry_proc_proc403_U0_start_full_n;
wire    Block_entry_proc_proc403_U0_start_write;
wire    tdf4_adjust_U0_start_full_n;
wire    tdf4_adjust_U0_start_write;
wire    tdf4_l2_multiply34_U0_start_full_n;
wire    tdf4_l2_multiply34_U0_start_write;
wire    tdf4_l2_writeOutputs_133_U0_start_full_n;
wire    tdf4_l2_writeOutputs_133_U0_start_write;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_sync_reg_tdf4_get_next_ijk_U0_ap_ready = 1'b0;
#0 ap_sync_reg_tdf4_readInputs37_U0_ap_ready = 1'b0;
end

td_fused_top_dataflow_in_loop_TOP_LOOP37832_ifmap_vec #(
    .DataWidth( 16 ),
    .AddressRange( 144 ),
    .AddressWidth( 8 ))
ifmap_vec_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf4_readInputs37_U0_ap_done),
    .i_full_n(ifmap_vec_i_full_n),
    .i_ce0(tdf4_readInputs37_U0_ifmap_vec_ce0),
    .i_we0(tdf4_readInputs37_U0_ifmap_vec_we0),
    .i_address0(tdf4_readInputs37_U0_ifmap_vec_address0),
    .i_d0(tdf4_readInputs37_U0_ifmap_vec_d0),
    .i_q0(ifmap_vec_i_q0),
    .i_ce1(tdf4_readInputs37_U0_ifmap_vec_ce1),
    .i_we1(tdf4_readInputs37_U0_ifmap_vec_we1),
    .i_address1(tdf4_readInputs37_U0_ifmap_vec_address1),
    .i_d1(tdf4_readInputs37_U0_ifmap_vec_d1),
    .t_ce(1'b1),
    .t_read(tdf4_dot_product_U0_ap_ready),
    .t_empty_n(ifmap_vec_t_empty_n),
    .t_ce0(tdf4_dot_product_U0_ifmap_vec_ce0),
    .t_we0(1'b0),
    .t_address0(tdf4_dot_product_U0_ifmap_vec_address0),
    .t_d0(16'd0),
    .t_q0(ifmap_vec_t_q0),
    .t_ce1(1'b0),
    .t_we1(1'b0),
    .t_address1(8'd0),
    .t_d1(16'd0)
);

td_fused_top_dataflow_in_loop_TOP_LOOP37832_weight_vecs_0 #(
    .DataWidth( 16 ),
    .AddressRange( 144 ),
    .AddressWidth( 8 ))
weight_vecs_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf4_readFilters36_U0_ap_done),
    .i_full_n(weight_vecs_0_i_full_n),
    .i_ce0(tdf4_readFilters36_U0_weight_vecs_0_ce0),
    .i_we0(tdf4_readFilters36_U0_weight_vecs_0_we0),
    .i_address0(tdf4_readFilters36_U0_weight_vecs_0_address0),
    .i_d0(tdf4_readFilters36_U0_weight_vecs_0_d0),
    .i_q0(weight_vecs_0_i_q0),
    .t_ce(1'b1),
    .t_read(tdf4_dot_product_U0_ap_ready),
    .t_empty_n(weight_vecs_0_t_empty_n),
    .t_ce0(tdf4_dot_product_U0_weight_vecs_0_ce0),
    .t_we0(1'b0),
    .t_address0(tdf4_dot_product_U0_weight_vecs_0_address0),
    .t_d0(16'd0),
    .t_q0(weight_vecs_0_t_q0)
);

td_fused_top_dataflow_in_loop_TOP_LOOP37832_products_0 #(
    .DataWidth( 16 ),
    .AddressRange( 144 ),
    .AddressWidth( 8 ))
products_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf4_dot_product_U0_ap_done),
    .i_full_n(products_0_i_full_n),
    .i_ce0(tdf4_dot_product_U0_products_0_ce0),
    .i_we0(tdf4_dot_product_U0_products_0_we0),
    .i_address0(tdf4_dot_product_U0_products_0_address0),
    .i_d0(tdf4_dot_product_U0_products_0_d0),
    .i_q0(products_0_i_q0),
    .i_ce1(1'b0),
    .i_address1(8'd0),
    .i_q1(products_0_i_q1),
    .t_ce(1'b1),
    .t_read(tdf4_accum_1_U0_ap_ready),
    .t_empty_n(products_0_t_empty_n),
    .t_ce0(tdf4_accum_1_U0_accum_in_0_ce0),
    .t_we0(1'b0),
    .t_address0(tdf4_accum_1_U0_accum_in_0_address0),
    .t_d0(16'd0),
    .t_q0(products_0_t_q0),
    .t_ce1(tdf4_accum_1_U0_accum_in_0_ce1),
    .t_address1(tdf4_accum_1_U0_accum_in_0_address1),
    .t_q1(products_0_t_q1)
);

td_fused_top_dataflow_in_loop_TOP_LOOP37832_accum1_out_0 #(
    .DataWidth( 16 ),
    .AddressRange( 8 ),
    .AddressWidth( 3 ))
accum1_out_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf4_accum_1_U0_ap_done),
    .i_full_n(accum1_out_0_i_full_n),
    .i_ce0(tdf4_accum_1_U0_accum_out_ce0),
    .i_we0(tdf4_accum_1_U0_accum_out_we0),
    .i_address0(tdf4_accum_1_U0_accum_out_address0),
    .i_d0(tdf4_accum_1_U0_accum_out_d0),
    .i_q0(accum1_out_0_i_q0),
    .i_ce1(tdf4_accum_1_U0_accum_out_ce1),
    .i_we1(tdf4_accum_1_U0_accum_out_we1),
    .i_address1(tdf4_accum_1_U0_accum_out_address1),
    .i_d1(tdf4_accum_1_U0_accum_out_d1),
    .t_ce(1'b1),
    .t_read(tdf4_accum_2_U0_ap_ready),
    .t_empty_n(accum1_out_0_t_empty_n),
    .t_ce0(tdf4_accum_2_U0_accum_in_ce0),
    .t_we0(1'b0),
    .t_address0(tdf4_accum_2_U0_accum_in_address0),
    .t_d0(16'd0),
    .t_q0(accum1_out_0_t_q0),
    .t_ce1(1'b0),
    .t_we1(1'b0),
    .t_address1(3'd0),
    .t_d1(16'd0)
);

td_fused_top_dataflow_in_loop_TOP_LOOP37832_l2_products #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
l2_products_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf4_l2_multiply34_U0_ap_done),
    .i_full_n(l2_products_i_full_n),
    .i_ce0(tdf4_l2_multiply34_U0_l2_products_ce0),
    .i_we0(tdf4_l2_multiply34_U0_l2_products_we0),
    .i_address0(tdf4_l2_multiply34_U0_l2_products_address0),
    .i_d0(tdf4_l2_multiply34_U0_l2_products_d0),
    .i_q0(l2_products_i_q0),
    .t_ce(1'b1),
    .t_read(tdf4_l2_writeOutputs_133_U0_ap_ready),
    .t_empty_n(l2_products_t_empty_n),
    .t_ce0(tdf4_l2_writeOutputs_133_U0_l2_partial_sums_ce0),
    .t_we0(1'b0),
    .t_address0(tdf4_l2_writeOutputs_133_U0_l2_partial_sums_address0),
    .t_d0(16'd0),
    .t_q0(l2_products_t_q0)
);

td_fused_top_tdf4_get_next_ijk tdf4_get_next_ijk_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf4_get_next_ijk_U0_ap_start),
    .start_full_n(start_for_tdf4_readFilters36_U0_full_n),
    .ap_done(tdf4_get_next_ijk_U0_ap_done),
    .ap_continue(tdf4_get_next_ijk_U0_ap_continue),
    .ap_idle(tdf4_get_next_ijk_U0_ap_idle),
    .ap_ready(tdf4_get_next_ijk_U0_ap_ready),
    .start_out(tdf4_get_next_ijk_U0_start_out),
    .start_write(tdf4_get_next_ijk_U0_start_write),
    .indices_0_din(tdf4_get_next_ijk_U0_indices_0_din),
    .indices_0_full_n(indices_01_c_full_n),
    .indices_0_write(tdf4_get_next_ijk_U0_indices_0_write),
    .indices_1_din(tdf4_get_next_ijk_U0_indices_1_din),
    .indices_1_full_n(indices_12_c_full_n),
    .indices_1_write(tdf4_get_next_ijk_U0_indices_1_write),
    .indices_2_out_din(tdf4_get_next_ijk_U0_indices_2_out_din),
    .indices_2_out_full_n(indices_23_c_full_n),
    .indices_2_out_write(tdf4_get_next_ijk_U0_indices_2_out_write),
    .indices_2_out1_din(tdf4_get_next_ijk_U0_indices_2_out1_din),
    .indices_2_out1_full_n(indices_23_c1_full_n),
    .indices_2_out1_write(tdf4_get_next_ijk_U0_indices_2_out1_write),
    .write_r_din(tdf4_get_next_ijk_U0_write_r_din),
    .write_r_full_n(write4_c_full_n),
    .write_r_write(tdf4_get_next_ijk_U0_write_r_write)
);

td_fused_top_tdf4_readInputs37 tdf4_readInputs37_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf4_readInputs37_U0_ap_start),
    .ap_done(tdf4_readInputs37_U0_ap_done),
    .ap_continue(tdf4_readInputs37_U0_ap_continue),
    .ap_idle(tdf4_readInputs37_U0_ap_idle),
    .ap_ready(tdf4_readInputs37_U0_ap_ready),
    .in_data_address0(tdf4_readInputs37_U0_in_data_address0),
    .in_data_ce0(tdf4_readInputs37_U0_in_data_ce0),
    .in_data_q0(in_data_q0),
    .indices_01_dout(indices_01_c_dout),
    .indices_01_empty_n(indices_01_c_empty_n),
    .indices_01_read(tdf4_readInputs37_U0_indices_01_read),
    .indices_12_dout(indices_12_c_dout),
    .indices_12_empty_n(indices_12_c_empty_n),
    .indices_12_read(tdf4_readInputs37_U0_indices_12_read),
    .ifmap_vec_address0(tdf4_readInputs37_U0_ifmap_vec_address0),
    .ifmap_vec_ce0(tdf4_readInputs37_U0_ifmap_vec_ce0),
    .ifmap_vec_we0(tdf4_readInputs37_U0_ifmap_vec_we0),
    .ifmap_vec_d0(tdf4_readInputs37_U0_ifmap_vec_d0),
    .ifmap_vec_address1(tdf4_readInputs37_U0_ifmap_vec_address1),
    .ifmap_vec_ce1(tdf4_readInputs37_U0_ifmap_vec_ce1),
    .ifmap_vec_we1(tdf4_readInputs37_U0_ifmap_vec_we1),
    .ifmap_vec_d1(tdf4_readInputs37_U0_ifmap_vec_d1),
    .indices_01_out_din(tdf4_readInputs37_U0_indices_01_out_din),
    .indices_01_out_full_n(indices_01_c2_full_n),
    .indices_01_out_write(tdf4_readInputs37_U0_indices_01_out_write),
    .indices_12_out_din(tdf4_readInputs37_U0_indices_12_out_din),
    .indices_12_out_full_n(indices_12_c3_full_n),
    .indices_12_out_write(tdf4_readInputs37_U0_indices_12_out_write)
);

td_fused_top_tdf4_readFilters36 tdf4_readFilters36_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf4_readFilters36_U0_ap_start),
    .ap_done(tdf4_readFilters36_U0_ap_done),
    .ap_continue(tdf4_readFilters36_U0_ap_continue),
    .ap_idle(tdf4_readFilters36_U0_ap_idle),
    .ap_ready(tdf4_readFilters36_U0_ap_ready),
    .filter_data_address0(tdf4_readFilters36_U0_filter_data_address0),
    .filter_data_ce0(tdf4_readFilters36_U0_filter_data_ce0),
    .filter_data_q0(l1_filter_data_q0),
    .indices_23_dout(indices_23_c_dout),
    .indices_23_empty_n(indices_23_c_empty_n),
    .indices_23_read(tdf4_readFilters36_U0_indices_23_read),
    .weight_vecs_0_address0(tdf4_readFilters36_U0_weight_vecs_0_address0),
    .weight_vecs_0_ce0(tdf4_readFilters36_U0_weight_vecs_0_ce0),
    .weight_vecs_0_we0(tdf4_readFilters36_U0_weight_vecs_0_we0),
    .weight_vecs_0_d0(tdf4_readFilters36_U0_weight_vecs_0_d0)
);

td_fused_top_tdf4_dot_product tdf4_dot_product_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf4_dot_product_U0_ap_start),
    .ap_done(tdf4_dot_product_U0_ap_done),
    .ap_continue(tdf4_dot_product_U0_ap_continue),
    .ap_idle(tdf4_dot_product_U0_ap_idle),
    .ap_ready(tdf4_dot_product_U0_ap_ready),
    .ifmap_vec_address0(tdf4_dot_product_U0_ifmap_vec_address0),
    .ifmap_vec_ce0(tdf4_dot_product_U0_ifmap_vec_ce0),
    .ifmap_vec_q0(ifmap_vec_t_q0),
    .weight_vecs_0_address0(tdf4_dot_product_U0_weight_vecs_0_address0),
    .weight_vecs_0_ce0(tdf4_dot_product_U0_weight_vecs_0_ce0),
    .weight_vecs_0_q0(weight_vecs_0_t_q0),
    .products_0_address0(tdf4_dot_product_U0_products_0_address0),
    .products_0_ce0(tdf4_dot_product_U0_products_0_ce0),
    .products_0_we0(tdf4_dot_product_U0_products_0_we0),
    .products_0_d0(tdf4_dot_product_U0_products_0_d0)
);

td_fused_top_tdf4_accum_1 tdf4_accum_1_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf4_accum_1_U0_ap_start),
    .ap_done(tdf4_accum_1_U0_ap_done),
    .ap_continue(tdf4_accum_1_U0_ap_continue),
    .ap_idle(tdf4_accum_1_U0_ap_idle),
    .ap_ready(tdf4_accum_1_U0_ap_ready),
    .accum_in_0_address0(tdf4_accum_1_U0_accum_in_0_address0),
    .accum_in_0_ce0(tdf4_accum_1_U0_accum_in_0_ce0),
    .accum_in_0_q0(products_0_t_q0),
    .accum_in_0_address1(tdf4_accum_1_U0_accum_in_0_address1),
    .accum_in_0_ce1(tdf4_accum_1_U0_accum_in_0_ce1),
    .accum_in_0_q1(products_0_t_q1),
    .accum_out_address0(tdf4_accum_1_U0_accum_out_address0),
    .accum_out_ce0(tdf4_accum_1_U0_accum_out_ce0),
    .accum_out_we0(tdf4_accum_1_U0_accum_out_we0),
    .accum_out_d0(tdf4_accum_1_U0_accum_out_d0),
    .accum_out_address1(tdf4_accum_1_U0_accum_out_address1),
    .accum_out_ce1(tdf4_accum_1_U0_accum_out_ce1),
    .accum_out_we1(tdf4_accum_1_U0_accum_out_we1),
    .accum_out_d1(tdf4_accum_1_U0_accum_out_d1)
);

td_fused_top_tdf4_accum_2 tdf4_accum_2_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf4_accum_2_U0_ap_start),
    .ap_done(tdf4_accum_2_U0_ap_done),
    .ap_continue(tdf4_accum_2_U0_ap_continue),
    .ap_idle(tdf4_accum_2_U0_ap_idle),
    .ap_ready(tdf4_accum_2_U0_ap_ready),
    .accum_in_12(tdf4_accum_2_U0_accum_in_12),
    .accum_in_12_ap_vld(tdf4_accum_2_U0_accum_in_12_ap_vld),
    .accum_in_address0(tdf4_accum_2_U0_accum_in_address0),
    .accum_in_ce0(tdf4_accum_2_U0_accum_in_ce0),
    .accum_in_q0(accum1_out_0_t_q0)
);

td_fused_top_Block_entry_proc_proc403 Block_entry_proc_proc403_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(Block_entry_proc_proc403_U0_ap_start),
    .ap_done(Block_entry_proc_proc403_U0_ap_done),
    .ap_continue(Block_entry_proc_proc403_U0_ap_continue),
    .ap_idle(Block_entry_proc_proc403_U0_ap_idle),
    .ap_ready(Block_entry_proc_proc403_U0_ap_ready),
    .tmp(tmp_channel_dout),
    .ap_return(Block_entry_proc_proc403_U0_ap_return)
);

td_fused_top_tdf4_adjust tdf4_adjust_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf4_adjust_U0_ap_start),
    .ap_done(tdf4_adjust_U0_ap_done),
    .ap_continue(tdf4_adjust_U0_ap_continue),
    .ap_idle(tdf4_adjust_U0_ap_idle),
    .ap_ready(tdf4_adjust_U0_ap_ready),
    .sums_read(sums_0_dout),
    .adjustments_address0(tdf4_adjust_U0_adjustments_address0),
    .adjustments_ce0(tdf4_adjust_U0_adjustments_ce0),
    .adjustments_q0(l1_adjustments_q0),
    .indices_23_dout(indices_23_c1_dout),
    .indices_23_empty_n(indices_23_c1_empty_n),
    .indices_23_read(tdf4_adjust_U0_indices_23_read),
    .indices_23_out_din(tdf4_adjust_U0_indices_23_out_din),
    .indices_23_out_full_n(indices_23_c4_full_n),
    .indices_23_out_write(tdf4_adjust_U0_indices_23_out_write),
    .ap_return(tdf4_adjust_U0_ap_return)
);

td_fused_top_tdf4_l2_multiply34 tdf4_l2_multiply34_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf4_l2_multiply34_U0_ap_start),
    .ap_done(tdf4_l2_multiply34_U0_ap_done),
    .ap_continue(tdf4_l2_multiply34_U0_ap_continue),
    .ap_idle(tdf4_l2_multiply34_U0_ap_idle),
    .ap_ready(tdf4_l2_multiply34_U0_ap_ready),
    .intermediate_fmaps_read(intermediate_fmaps_0_dout),
    .l2_filter_data_address0(tdf4_l2_multiply34_U0_l2_filter_data_address0),
    .l2_filter_data_ce0(tdf4_l2_multiply34_U0_l2_filter_data_ce0),
    .l2_filter_data_q0(l2_filter_data_q0),
    .l2_products_address0(tdf4_l2_multiply34_U0_l2_products_address0),
    .l2_products_ce0(tdf4_l2_multiply34_U0_l2_products_ce0),
    .l2_products_we0(tdf4_l2_multiply34_U0_l2_products_we0),
    .l2_products_d0(tdf4_l2_multiply34_U0_l2_products_d0),
    .indices_23_dout(indices_23_c4_dout),
    .indices_23_empty_n(indices_23_c4_empty_n),
    .indices_23_read(tdf4_l2_multiply34_U0_indices_23_read)
);

td_fused_top_tdf4_l2_writeOutputs_133 tdf4_l2_writeOutputs_133_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf4_l2_writeOutputs_133_U0_ap_start),
    .ap_done(tdf4_l2_writeOutputs_133_U0_ap_done),
    .ap_continue(tdf4_l2_writeOutputs_133_U0_ap_continue),
    .ap_idle(tdf4_l2_writeOutputs_133_U0_ap_idle),
    .ap_ready(tdf4_l2_writeOutputs_133_U0_ap_ready),
    .indices_01_dout(indices_01_c2_dout),
    .indices_01_empty_n(indices_01_c2_empty_n),
    .indices_01_read(tdf4_l2_writeOutputs_133_U0_indices_01_read),
    .indices_12_dout(indices_12_c3_dout),
    .indices_12_empty_n(indices_12_c3_empty_n),
    .indices_12_read(tdf4_l2_writeOutputs_133_U0_indices_12_read),
    .write4_dout(write4_c_dout),
    .write4_empty_n(write4_c_empty_n),
    .write4_read(tdf4_l2_writeOutputs_133_U0_write4_read),
    .l2_partial_sums_address0(tdf4_l2_writeOutputs_133_U0_l2_partial_sums_address0),
    .l2_partial_sums_ce0(tdf4_l2_writeOutputs_133_U0_l2_partial_sums_ce0),
    .l2_partial_sums_q0(l2_products_t_q0),
    .out_data_address1(tdf4_l2_writeOutputs_133_U0_out_data_address1),
    .out_data_ce1(tdf4_l2_writeOutputs_133_U0_out_data_ce1),
    .out_data_we1(tdf4_l2_writeOutputs_133_U0_out_data_we1),
    .out_data_d1(tdf4_l2_writeOutputs_133_U0_out_data_d1),
    .l2_adjustments_address0(tdf4_l2_writeOutputs_133_U0_l2_adjustments_address0),
    .l2_adjustments_ce0(tdf4_l2_writeOutputs_133_U0_l2_adjustments_ce0),
    .l2_adjustments_q0(l2_adjustments_q0)
);

td_fused_top_fifo_w16_d2_S_x1 indices_01_c_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(indices_01_c_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf4_readInputs37_U0_indices_01_read),
    .if_dout(indices_01_c_dout),
    .if_full_n(indices_01_c_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf4_get_next_ijk_U0_indices_0_write),
    .if_din(tdf4_get_next_ijk_U0_indices_0_din)
);

td_fused_top_fifo_w16_d2_S_x1 indices_12_c_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(indices_12_c_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf4_readInputs37_U0_indices_12_read),
    .if_dout(indices_12_c_dout),
    .if_full_n(indices_12_c_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf4_get_next_ijk_U0_indices_1_write),
    .if_din(tdf4_get_next_ijk_U0_indices_1_din)
);

td_fused_top_fifo_w7_d2_S indices_23_c_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(indices_23_c_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf4_readFilters36_U0_indices_23_read),
    .if_dout(indices_23_c_dout),
    .if_full_n(indices_23_c_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf4_get_next_ijk_U0_indices_2_out_write),
    .if_din(tdf4_get_next_ijk_U0_indices_2_out_din)
);

td_fused_top_fifo_w11_d7_S indices_23_c1_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(indices_23_c1_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf4_adjust_U0_indices_23_read),
    .if_dout(indices_23_c1_dout),
    .if_full_n(indices_23_c1_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf4_get_next_ijk_U0_indices_2_out1_write),
    .if_din(tdf4_get_next_ijk_U0_indices_2_out1_din)
);

td_fused_top_fifo_w1_d9_S_x write4_c_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(write4_c_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf4_l2_writeOutputs_133_U0_write4_read),
    .if_dout(write4_c_dout),
    .if_full_n(write4_c_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf4_get_next_ijk_U0_write_r_write),
    .if_din(write4_c_din)
);

td_fused_top_fifo_w6_d8_S_x indices_01_c2_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(indices_01_c2_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf4_l2_writeOutputs_133_U0_indices_01_read),
    .if_dout(indices_01_c2_dout),
    .if_full_n(indices_01_c2_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf4_readInputs37_U0_indices_01_out_write),
    .if_din(tdf4_readInputs37_U0_indices_01_out_din)
);

td_fused_top_fifo_w12_d8_S_x indices_12_c3_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(indices_12_c3_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf4_l2_writeOutputs_133_U0_indices_12_read),
    .if_dout(indices_12_c3_dout),
    .if_full_n(indices_12_c3_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf4_readInputs37_U0_indices_12_out_write),
    .if_din(tdf4_readInputs37_U0_indices_12_out_din)
);

td_fused_top_fifo_w16_d2_S_x1 tmp_channel_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(tmp_channel_empty_n),
    .if_read_ce(1'b1),
    .if_read(Block_entry_proc_proc403_U0_ap_ready),
    .if_dout(tmp_channel_dout),
    .if_full_n(tmp_channel_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf4_accum_2_U0_ap_done),
    .if_din(tdf4_accum_2_U0_accum_in_12)
);

td_fused_top_fifo_w16_d2_S_x1 sums_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(sums_0_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf4_adjust_U0_ap_ready),
    .if_dout(sums_0_dout),
    .if_full_n(sums_0_full_n),
    .if_write_ce(1'b1),
    .if_write(Block_entry_proc_proc403_U0_ap_done),
    .if_din(Block_entry_proc_proc403_U0_ap_return)
);

td_fused_top_fifo_w11_d2_S indices_23_c4_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(indices_23_c4_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf4_l2_multiply34_U0_indices_23_read),
    .if_dout(indices_23_c4_dout),
    .if_full_n(indices_23_c4_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf4_adjust_U0_indices_23_out_write),
    .if_din(tdf4_adjust_U0_indices_23_out_din)
);

td_fused_top_fifo_w16_d2_S_x1 intermediate_fmaps_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(intermediate_fmaps_0_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf4_l2_multiply34_U0_ap_ready),
    .if_dout(intermediate_fmaps_0_dout),
    .if_full_n(intermediate_fmaps_0_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf4_adjust_U0_ap_done),
    .if_din(tdf4_adjust_U0_ap_return)
);

td_fused_top_start_for_tdf4_readFilters36_U0 start_for_tdf4_readFilters36_U0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(start_for_tdf4_readFilters36_U0_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf4_readFilters36_U0_ap_ready),
    .if_dout(start_for_tdf4_readFilters36_U0_dout),
    .if_full_n(start_for_tdf4_readFilters36_U0_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf4_get_next_ijk_U0_start_write),
    .if_din(start_for_tdf4_readFilters36_U0_din)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_sync_reg_tdf4_get_next_ijk_U0_ap_ready <= 1'b0;
    end else begin
        if (((ap_sync_ready & ap_start) == 1'b1)) begin
            ap_sync_reg_tdf4_get_next_ijk_U0_ap_ready <= 1'b0;
        end else begin
            ap_sync_reg_tdf4_get_next_ijk_U0_ap_ready <= ap_sync_tdf4_get_next_ijk_U0_ap_ready;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_sync_reg_tdf4_readInputs37_U0_ap_ready <= 1'b0;
    end else begin
        if (((ap_sync_ready & ap_start) == 1'b1)) begin
            ap_sync_reg_tdf4_readInputs37_U0_ap_ready <= 1'b0;
        end else begin
            ap_sync_reg_tdf4_readInputs37_U0_ap_ready <= ap_sync_tdf4_readInputs37_U0_ap_ready;
        end
    end
end

assign Block_entry_proc_proc403_U0_ap_continue = sums_0_full_n;

assign Block_entry_proc_proc403_U0_ap_start = tmp_channel_empty_n;

assign Block_entry_proc_proc403_U0_start_full_n = 1'b1;

assign Block_entry_proc_proc403_U0_start_write = 1'b0;

assign ap_channel_done_accum1_out_0 = tdf4_accum_1_U0_ap_done;

assign ap_channel_done_ifmap_vec = tdf4_readInputs37_U0_ap_done;

assign ap_channel_done_intermediate_fmaps_0 = tdf4_adjust_U0_ap_done;

assign ap_channel_done_l2_products = tdf4_l2_multiply34_U0_ap_done;

assign ap_channel_done_products_0 = tdf4_dot_product_U0_ap_done;

assign ap_channel_done_sums_0 = Block_entry_proc_proc403_U0_ap_done;

assign ap_channel_done_tmp_channel = tdf4_accum_2_U0_ap_done;

assign ap_channel_done_weight_vecs_0 = tdf4_readFilters36_U0_ap_done;

assign ap_done = tdf4_l2_writeOutputs_133_U0_ap_done;

assign ap_idle = (tdf4_readInputs37_U0_ap_idle & tdf4_readFilters36_U0_ap_idle & tdf4_l2_writeOutputs_133_U0_ap_idle & tdf4_l2_multiply34_U0_ap_idle & tdf4_get_next_ijk_U0_ap_idle & tdf4_dot_product_U0_ap_idle & tdf4_adjust_U0_ap_idle & tdf4_accum_2_U0_ap_idle & tdf4_accum_1_U0_ap_idle & (intermediate_fmaps_0_empty_n ^ 1'b1) & (sums_0_empty_n ^ 1'b1) & (tmp_channel_empty_n ^ 1'b1) & (l2_products_t_empty_n ^ 1'b1) & (products_0_t_empty_n ^ 1'b1) & (weight_vecs_0_t_empty_n ^ 1'b1) & (ifmap_vec_t_empty_n ^ 1'b1) & (1'b1 ^ accum1_out_0_t_empty_n) & Block_entry_proc_proc403_U0_ap_idle);

assign ap_ready = ap_sync_ready;

assign ap_sync_continue = ap_continue;

assign ap_sync_done = tdf4_l2_writeOutputs_133_U0_ap_done;

assign ap_sync_ready = (ap_sync_tdf4_readInputs37_U0_ap_ready & ap_sync_tdf4_get_next_ijk_U0_ap_ready);

assign ap_sync_tdf4_get_next_ijk_U0_ap_ready = (tdf4_get_next_ijk_U0_ap_ready | ap_sync_reg_tdf4_get_next_ijk_U0_ap_ready);

assign ap_sync_tdf4_readInputs37_U0_ap_ready = (tdf4_readInputs37_U0_ap_ready | ap_sync_reg_tdf4_readInputs37_U0_ap_ready);

assign in_data_address0 = tdf4_readInputs37_U0_in_data_address0;

assign in_data_address1 = 14'd0;

assign in_data_ce0 = tdf4_readInputs37_U0_in_data_ce0;

assign in_data_ce1 = 1'b0;

assign in_data_d0 = 64'd0;

assign in_data_d1 = 64'd0;

assign in_data_read = tdf4_readInputs37_U0_in_data_write;

assign in_data_we0 = 1'b0;

assign in_data_we1 = 1'b0;

assign l1_adjustments_address0 = tdf4_adjust_U0_adjustments_address0;

assign l1_adjustments_address1 = 7'd0;

assign l1_adjustments_ce0 = tdf4_adjust_U0_adjustments_ce0;

assign l1_adjustments_ce1 = 1'b0;

assign l1_adjustments_d0 = 48'd0;

assign l1_adjustments_d1 = 48'd0;

assign l1_adjustments_we0 = 1'b0;

assign l1_adjustments_we1 = 1'b0;

assign l1_filter_data_address0 = tdf4_readFilters36_U0_filter_data_address0;

assign l1_filter_data_address1 = 15'd0;

assign l1_filter_data_ce0 = tdf4_readFilters36_U0_filter_data_ce0;

assign l1_filter_data_ce1 = 1'b0;

assign l1_filter_data_d0 = 16'd0;

assign l1_filter_data_d1 = 16'd0;

assign l1_filter_data_we0 = 1'b0;

assign l1_filter_data_we1 = 1'b0;

assign l2_adjustments_address0 = tdf4_l2_writeOutputs_133_U0_l2_adjustments_address0;

assign l2_adjustments_address1 = 4'd0;

assign l2_adjustments_ce0 = tdf4_l2_writeOutputs_133_U0_l2_adjustments_ce0;

assign l2_adjustments_ce1 = 1'b0;

assign l2_adjustments_d0 = 48'd0;

assign l2_adjustments_d1 = 48'd0;

assign l2_adjustments_we0 = 1'b0;

assign l2_adjustments_we1 = 1'b0;

assign l2_filter_data_address0 = tdf4_l2_multiply34_U0_l2_filter_data_address0;

assign l2_filter_data_address1 = 11'd0;

assign l2_filter_data_ce0 = tdf4_l2_multiply34_U0_l2_filter_data_ce0;

assign l2_filter_data_ce1 = 1'b0;

assign l2_filter_data_d0 = 16'd0;

assign l2_filter_data_d1 = 16'd0;

assign l2_filter_data_we0 = 1'b0;

assign l2_filter_data_we1 = 1'b0;

assign out_data_address0 = 14'd0;

assign out_data_address1 = tdf4_l2_writeOutputs_133_U0_out_data_address1;

assign out_data_ce0 = 1'b0;

assign out_data_ce1 = tdf4_l2_writeOutputs_133_U0_out_data_ce1;

assign out_data_d0 = 64'd0;

assign out_data_d1 = tdf4_l2_writeOutputs_133_U0_out_data_d1;

assign out_data_we0 = 1'b0;

assign out_data_we1 = tdf4_l2_writeOutputs_133_U0_out_data_we1;

assign out_data_write = tdf4_l2_writeOutputs_133_U0_out_data_write;

assign products_0_t_d1 = 16'd0;

assign products_0_t_we1 = 1'b0;

assign start_for_tdf4_readFilters36_U0_din = 1'b1;

assign tdf4_accum_1_U0_accum_out_full_n = accum1_out_0_i_full_n;

assign tdf4_accum_1_U0_ap_continue = accum1_out_0_i_full_n;

assign tdf4_accum_1_U0_ap_start = products_0_t_empty_n;

assign tdf4_accum_1_U0_start_full_n = 1'b1;

assign tdf4_accum_1_U0_start_write = 1'b0;

assign tdf4_accum_2_U0_ap_continue = tmp_channel_full_n;

assign tdf4_accum_2_U0_ap_start = accum1_out_0_t_empty_n;

assign tdf4_accum_2_U0_start_full_n = 1'b1;

assign tdf4_accum_2_U0_start_write = 1'b0;

assign tdf4_adjust_U0_ap_continue = intermediate_fmaps_0_full_n;

assign tdf4_adjust_U0_ap_start = sums_0_empty_n;

assign tdf4_adjust_U0_start_full_n = 1'b1;

assign tdf4_adjust_U0_start_write = 1'b0;

assign tdf4_dot_product_U0_ap_continue = products_0_i_full_n;

assign tdf4_dot_product_U0_ap_start = (weight_vecs_0_t_empty_n & ifmap_vec_t_empty_n);

assign tdf4_dot_product_U0_products_0_full_n = products_0_i_full_n;

assign tdf4_dot_product_U0_start_full_n = 1'b1;

assign tdf4_dot_product_U0_start_write = 1'b0;

assign tdf4_get_next_ijk_U0_ap_continue = 1'b1;

assign tdf4_get_next_ijk_U0_ap_start = ((ap_sync_reg_tdf4_get_next_ijk_U0_ap_ready ^ 1'b1) & ap_start);

assign tdf4_l2_multiply34_U0_ap_continue = l2_products_i_full_n;

assign tdf4_l2_multiply34_U0_ap_start = intermediate_fmaps_0_empty_n;

assign tdf4_l2_multiply34_U0_l2_products_full_n = l2_products_i_full_n;

assign tdf4_l2_multiply34_U0_start_full_n = 1'b1;

assign tdf4_l2_multiply34_U0_start_write = 1'b0;

assign tdf4_l2_writeOutputs_133_U0_ap_continue = ap_continue;

assign tdf4_l2_writeOutputs_133_U0_ap_start = l2_products_t_empty_n;

assign tdf4_l2_writeOutputs_133_U0_out_data_full_n = out_data_full_n;

assign tdf4_l2_writeOutputs_133_U0_out_data_write = 1'b0;

assign tdf4_l2_writeOutputs_133_U0_start_full_n = 1'b1;

assign tdf4_l2_writeOutputs_133_U0_start_write = 1'b0;

assign tdf4_readFilters36_U0_ap_continue = weight_vecs_0_i_full_n;

assign tdf4_readFilters36_U0_ap_start = start_for_tdf4_readFilters36_U0_empty_n;

assign tdf4_readFilters36_U0_start_full_n = 1'b1;

assign tdf4_readFilters36_U0_start_write = 1'b0;

assign tdf4_readFilters36_U0_weight_vecs_0_full_n = weight_vecs_0_i_full_n;

assign tdf4_readInputs37_U0_ap_continue = ifmap_vec_i_full_n;

assign tdf4_readInputs37_U0_ap_start = ((ap_sync_reg_tdf4_readInputs37_U0_ap_ready ^ 1'b1) & ap_start);

assign tdf4_readInputs37_U0_ifmap_vec_full_n = ifmap_vec_i_full_n;

assign tdf4_readInputs37_U0_in_data_full_n = in_data_empty_n;

assign tdf4_readInputs37_U0_in_data_write = 1'b0;

assign tdf4_readInputs37_U0_start_full_n = 1'b1;

assign tdf4_readInputs37_U0_start_write = 1'b0;

assign write4_c_din = tdf4_get_next_ijk_U0_write_r_din;

endmodule //td_fused_top_dataflow_in_loop_TOP_LOOP37832
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37832_weight_vecs_0_memcore_ram (addr0, ce0, d0, we0, q0, addr1, ce1, d1, we1, q1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 9;
parameter MEM_SIZE = 288;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
output reg[DWIDTH-1:0] q1;
input clk;

reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];




always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1) 
            ram[addr1] <= d1; 
        q1 <= ram[addr1];
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37832_weight_vecs_0_memcore(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    q0,
    address1,
    ce1,
    we1,
    d1,
    q1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd288;
parameter AddressWidth = 32'd9;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;
output[DataWidth - 1:0] q1;



td_fused_top_dataflow_in_loop_TOP_LOOP37832_weight_vecs_0_memcore_ram td_fused_top_dataflow_in_loop_TOP_LOOP37832_weight_vecs_0_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 ),
    .q1( q1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_dataflow_in_loop_TOP_LOOP37832_weight_vecs_0
#(parameter
    DataWidth    = 16,
    AddressRange = 32,
    AddressWidth = 8,
    BufferCount  = 2,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire                    i_we0,
    input  wire [AddressWidth-1:0] i_address0,
    input  wire [DataWidth-1:0]    i_d0,
    output wire [DataWidth-1:0]    i_q0,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire                    t_we0,
    input  wire [AddressWidth-1:0] t_address0,
    input  wire [DataWidth-1:0]    t_d0,
    output wire [DataWidth-1:0]    t_q0
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
wire [AddressWidth+IndexWidth-1:0]   memcore_iaddr;
wire [AddressWidth+IndexWidth-1:0]   memcore_taddr;

//------------------------Instantiation------------------
assign memcore_iaddr = {i_address0, iptr};
assign memcore_taddr = {t_address0, tptr};
td_fused_top_dataflow_in_loop_TOP_LOOP37832_weight_vecs_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP37832_weight_vecs_0_memcore_U (
    .reset    ( reset ),
    .clk      ( clk ),
    .address0 ( memcore_iaddr ),
    .ce0      ( i_ce0 ),
    .we0      ( i_we0),
    .d0       ( i_d0 ),
    .q0       ( i_q0 ),
    .address1 ( memcore_taddr ),
    .ce1      ( t_ce0 ),
    .we1      ( t_we0),
    .d1       ( t_d0 ),
    .q1       ( t_q0 )

);

//------------------------Body---------------------------

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37928_accum1_out_0_memcore_ram (addr0, ce0, d0, we0, q0, addr1, ce1, d1, we1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 3;
parameter MEM_SIZE = 8;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
input clk;

reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];




always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1) 
            ram[addr1] <= d1; 
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37928_accum1_out_0_memcore(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    q0,
    address1,
    ce1,
    we1,
    d1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd8;
parameter AddressWidth = 32'd3;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;



td_fused_top_dataflow_in_loop_TOP_LOOP37928_accum1_out_0_memcore_ram td_fused_top_dataflow_in_loop_TOP_LOOP37928_accum1_out_0_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_dataflow_in_loop_TOP_LOOP37928_accum1_out_0
#(parameter
    DataWidth    = 16,
    AddressRange = 32,
    AddressWidth = 3,
    BufferCount  = 2,
    MemLatency   = 1,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire                    i_we0,
    input  wire [AddressWidth-1:0] i_address0,
    input  wire [DataWidth-1:0]    i_d0,
    output wire [DataWidth-1:0]    i_q0,
    input  wire                    i_ce1,
    input  wire                    i_we1,
    input  wire [AddressWidth-1:0] i_address1,
    input  wire [DataWidth-1:0]    i_d1,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire                    t_we0,
    input  wire [AddressWidth-1:0] t_address0,
    input  wire [DataWidth-1:0]    t_d0,
    output wire [DataWidth-1:0]    t_q0,
    input  wire                    t_ce1,
    input  wire                    t_we1,
    input  wire [AddressWidth-1:0] t_address1,
    input  wire [DataWidth-1:0]    t_d1
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth-1:0]   prev_iptr    = 1'b0; // previous initiator index
reg  [IndexWidth-1:0]   prev_tptr    = 1'b0; // previous target index
reg  [DataWidth-1:0]    reg_q0      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid0    = 1'b0; // buffer has valid data
reg  [DataWidth-1:0]    reg_q1      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid1    = 1'b0; // buffer has valid data
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
// buffer signals
wire [BufferCount-1:0] buf_ce0;
wire [BufferCount-1:0] buf_we0;
wire [AddressWidth-1:0] buf_a0_0, buf_a0_1;
wire [DataWidth-1:0] buf_d0_0, buf_d0_1;
wire [DataWidth-1:0] buf_q0_0, buf_q0_1;
wire [BufferCount-1:0] buf_ce1;
wire [BufferCount-1:0] buf_we1;
wire [AddressWidth-1:0] buf_a1_0, buf_a1_1;
wire [DataWidth-1:0] buf_d1_0, buf_d1_1;
//------------------------Instantiation------------------
//genvar i;
        td_fused_top_dataflow_in_loop_TOP_LOOP37928_accum1_out_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP37928_accum1_out_0_memcore_U_0 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_0 ),
            .ce0      ( buf_ce0[ 0 ] ),
            .we0      ( buf_we0[ 0 ] ),
            .d0       ( buf_d0_0 ),
            .q0       ( buf_q0_0 ),
            .address1 ( buf_a1_0 ),
            .ce1      ( buf_ce1[ 0 ] ),
            .we1      ( buf_we1[ 0 ] ),
            .d1       ( buf_d1_0 )
        );
        td_fused_top_dataflow_in_loop_TOP_LOOP37928_accum1_out_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP37928_accum1_out_0_memcore_U_1 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_1 ),
            .ce0      ( buf_ce0[ 1 ] ),
            .we0      ( buf_we0[ 1 ] ),
            .d0       ( buf_d0_1 ),
            .q0       ( buf_q0_1 ),
            .address1 ( buf_a1_1 ),
            .ce1      ( buf_ce1[ 1 ] ),
            .we1      ( buf_we1[ 1 ] ),
            .d1       ( buf_d1_1 )
        );

//++++++++++++++++++++++++buffer signals+++++++++++++++++
        assign buf_ce0[ 0 ] = (tptr ==  0  && empty_n) ? t_ce0
                             : (iptr ==  0 ) ? i_ce0 : 1'b0;
        assign buf_a0_0  = (tptr ==  0  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 0 ] = (tptr ==  0  && empty_n)  ? t_we0
                             : (iptr ==  0 ) ? i_we0 : 1'b0;
        assign buf_d0_0  = (tptr ==  0  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 0 ] = (tptr ==  0  && empty_n) ? t_ce1
                             : (iptr ==  0 ) ? i_ce1 : 1'b0;
        assign buf_a1_0  = (tptr ==  0  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 0 ] = (tptr ==  0  && empty_n)  ? t_we1
                             : (iptr ==  0 ) ? i_we1 : 1'b0;
        assign buf_d1_0  = (tptr ==  0  && empty_n) ? t_d1       : i_d1;
        assign buf_ce0[ 1 ] = (tptr ==  1  && empty_n) ? t_ce0
                             : (iptr ==  1 ) ? i_ce0 : 1'b0;
        assign buf_a0_1  = (tptr ==  1  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 1 ] = (tptr ==  1  && empty_n)  ? t_we0
                             : (iptr ==  1 ) ? i_we0 : 1'b0;
        assign buf_d0_1  = (tptr ==  1  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 1 ] = (tptr ==  1  && empty_n) ? t_ce1
                             : (iptr ==  1 ) ? i_ce1 : 1'b0;
        assign buf_a1_1  = (tptr ==  1  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 1 ] = (tptr ==  1  && empty_n)  ? t_we1
                             : (iptr ==  1 ) ? i_we1 : 1'b0;
        assign buf_d1_1  = (tptr ==  1  && empty_n) ? t_d1       : i_d1;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//------------------------Body---------------------------
assign i_q0      = (prev_iptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign t_q0      = reg_valid0 ? reg_q0 : (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// prev_iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_iptr <= 1'b0;
    else begin
        prev_iptr <= iptr;
    end
end

// prev_tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_tptr <= 1'b0;
    else begin
        prev_tptr <= tptr;
    end
end

// reg_q0 and reg_valid0
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q0     <= 1'b0;
        reg_valid0 <= 1'b0;
    end else if (!t_ce0 && !reg_valid0) begin
        reg_q0     <= (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
        reg_valid0 <= 1'b1;
    end else if (t_ce0) begin
        reg_valid0 <= 1'b0;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37928_ifmap_vec_0_0_memcore_ram (addr0, ce0, d0, we0, q0, addr1, ce1, d1, we1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 5;
parameter MEM_SIZE = 32;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
input clk;

reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];




always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1) 
            ram[addr1] <= d1; 
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37928_ifmap_vec_0_0_memcore(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    q0,
    address1,
    ce1,
    we1,
    d1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd32;
parameter AddressWidth = 32'd5;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;



td_fused_top_dataflow_in_loop_TOP_LOOP37928_ifmap_vec_0_0_memcore_ram td_fused_top_dataflow_in_loop_TOP_LOOP37928_ifmap_vec_0_0_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_dataflow_in_loop_TOP_LOOP37928_ifmap_vec_0_0
#(parameter
    DataWidth    = 16,
    AddressRange = 32,
    AddressWidth = 5,
    BufferCount  = 2,
    MemLatency   = 1,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire                    i_we0,
    input  wire [AddressWidth-1:0] i_address0,
    input  wire [DataWidth-1:0]    i_d0,
    output wire [DataWidth-1:0]    i_q0,
    input  wire                    i_ce1,
    input  wire                    i_we1,
    input  wire [AddressWidth-1:0] i_address1,
    input  wire [DataWidth-1:0]    i_d1,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire                    t_we0,
    input  wire [AddressWidth-1:0] t_address0,
    input  wire [DataWidth-1:0]    t_d0,
    output wire [DataWidth-1:0]    t_q0,
    input  wire                    t_ce1,
    input  wire                    t_we1,
    input  wire [AddressWidth-1:0] t_address1,
    input  wire [DataWidth-1:0]    t_d1
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth-1:0]   prev_iptr    = 1'b0; // previous initiator index
reg  [IndexWidth-1:0]   prev_tptr    = 1'b0; // previous target index
reg  [DataWidth-1:0]    reg_q0      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid0    = 1'b0; // buffer has valid data
reg  [DataWidth-1:0]    reg_q1      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid1    = 1'b0; // buffer has valid data
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
// buffer signals
wire [BufferCount-1:0] buf_ce0;
wire [BufferCount-1:0] buf_we0;
wire [AddressWidth-1:0] buf_a0_0, buf_a0_1;
wire [DataWidth-1:0] buf_d0_0, buf_d0_1;
wire [DataWidth-1:0] buf_q0_0, buf_q0_1;
wire [BufferCount-1:0] buf_ce1;
wire [BufferCount-1:0] buf_we1;
wire [AddressWidth-1:0] buf_a1_0, buf_a1_1;
wire [DataWidth-1:0] buf_d1_0, buf_d1_1;
//------------------------Instantiation------------------
//genvar i;
        td_fused_top_dataflow_in_loop_TOP_LOOP37928_ifmap_vec_0_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP37928_ifmap_vec_0_0_memcore_U_0 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_0 ),
            .ce0      ( buf_ce0[ 0 ] ),
            .we0      ( buf_we0[ 0 ] ),
            .d0       ( buf_d0_0 ),
            .q0       ( buf_q0_0 ),
            .address1 ( buf_a1_0 ),
            .ce1      ( buf_ce1[ 0 ] ),
            .we1      ( buf_we1[ 0 ] ),
            .d1       ( buf_d1_0 )
        );
        td_fused_top_dataflow_in_loop_TOP_LOOP37928_ifmap_vec_0_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP37928_ifmap_vec_0_0_memcore_U_1 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_1 ),
            .ce0      ( buf_ce0[ 1 ] ),
            .we0      ( buf_we0[ 1 ] ),
            .d0       ( buf_d0_1 ),
            .q0       ( buf_q0_1 ),
            .address1 ( buf_a1_1 ),
            .ce1      ( buf_ce1[ 1 ] ),
            .we1      ( buf_we1[ 1 ] ),
            .d1       ( buf_d1_1 )
        );

//++++++++++++++++++++++++buffer signals+++++++++++++++++
        assign buf_ce0[ 0 ] = (tptr ==  0  && empty_n) ? t_ce0
                             : (iptr ==  0 ) ? i_ce0 : 1'b0;
        assign buf_a0_0  = (tptr ==  0  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 0 ] = (tptr ==  0  && empty_n)  ? t_we0
                             : (iptr ==  0 ) ? i_we0 : 1'b0;
        assign buf_d0_0  = (tptr ==  0  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 0 ] = (tptr ==  0  && empty_n) ? t_ce1
                             : (iptr ==  0 ) ? i_ce1 : 1'b0;
        assign buf_a1_0  = (tptr ==  0  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 0 ] = (tptr ==  0  && empty_n)  ? t_we1
                             : (iptr ==  0 ) ? i_we1 : 1'b0;
        assign buf_d1_0  = (tptr ==  0  && empty_n) ? t_d1       : i_d1;
        assign buf_ce0[ 1 ] = (tptr ==  1  && empty_n) ? t_ce0
                             : (iptr ==  1 ) ? i_ce0 : 1'b0;
        assign buf_a0_1  = (tptr ==  1  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 1 ] = (tptr ==  1  && empty_n)  ? t_we0
                             : (iptr ==  1 ) ? i_we0 : 1'b0;
        assign buf_d0_1  = (tptr ==  1  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 1 ] = (tptr ==  1  && empty_n) ? t_ce1
                             : (iptr ==  1 ) ? i_ce1 : 1'b0;
        assign buf_a1_1  = (tptr ==  1  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 1 ] = (tptr ==  1  && empty_n)  ? t_we1
                             : (iptr ==  1 ) ? i_we1 : 1'b0;
        assign buf_d1_1  = (tptr ==  1  && empty_n) ? t_d1       : i_d1;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//------------------------Body---------------------------
assign i_q0      = (prev_iptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign t_q0      = reg_valid0 ? reg_q0 : (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// prev_iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_iptr <= 1'b0;
    else begin
        prev_iptr <= iptr;
    end
end

// prev_tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_tptr <= 1'b0;
    else begin
        prev_tptr <= tptr;
    end
end

// reg_q0 and reg_valid0
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q0     <= 1'b0;
        reg_valid0 <= 1'b0;
    end else if (!t_ce0 && !reg_valid0) begin
        reg_q0     <= (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
        reg_valid0 <= 1'b1;
    end else if (t_ce0) begin
        reg_valid0 <= 1'b0;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37928_products_0_memcore_ram (addr0, ce0, d0, we0, q0, addr1, ce1, q1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 5;
parameter MEM_SIZE = 32;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
output reg[DWIDTH-1:0] q1;
input clk;

reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];




always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        q1 <= ram[addr1];
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37928_products_0_memcore(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    q0,
    address1,
    ce1,
    q1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd32;
parameter AddressWidth = 32'd5;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
output[DataWidth - 1:0] q1;



td_fused_top_dataflow_in_loop_TOP_LOOP37928_products_0_memcore_ram td_fused_top_dataflow_in_loop_TOP_LOOP37928_products_0_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .q1( q1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_dataflow_in_loop_TOP_LOOP37928_products_0
#(parameter
    DataWidth    = 16,
    AddressRange = 32,
    AddressWidth = 5,
    BufferCount  = 2,
    MemLatency   = 1,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire                    i_we0,
    input  wire [AddressWidth-1:0] i_address0,
    input  wire [DataWidth-1:0]    i_d0,
    output wire [DataWidth-1:0]    i_q0,
    input  wire                    i_ce1,
    input  wire [AddressWidth-1:0] i_address1,
    output wire [DataWidth-1:0]    i_q1,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire                    t_we0,
    input  wire [AddressWidth-1:0] t_address0,
    input  wire [DataWidth-1:0]    t_d0,
    output wire [DataWidth-1:0]    t_q0,
    input  wire                    t_ce1,
    input  wire [AddressWidth-1:0] t_address1,
    output wire [DataWidth-1:0]    t_q1
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth-1:0]   prev_iptr    = 1'b0; // previous initiator index
reg  [IndexWidth-1:0]   prev_tptr    = 1'b0; // previous target index
reg  [DataWidth-1:0]    reg_q0      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid0    = 1'b0; // buffer has valid data
reg  [DataWidth-1:0]    reg_q1      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid1    = 1'b0; // buffer has valid data
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
// buffer signals
wire [BufferCount-1:0] buf_ce0;
wire [BufferCount-1:0] buf_we0;
wire [AddressWidth-1:0] buf_a0_0, buf_a0_1;
wire [DataWidth-1:0] buf_d0_0, buf_d0_1;
wire [DataWidth-1:0] buf_q0_0, buf_q0_1;
wire [BufferCount-1:0] buf_ce1;
wire [AddressWidth-1:0] buf_a1_0, buf_a1_1;
wire [DataWidth-1:0] buf_q1_0, buf_q1_1;
//------------------------Instantiation------------------
//genvar i;
        td_fused_top_dataflow_in_loop_TOP_LOOP37928_products_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP37928_products_0_memcore_U_0 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_0 ),
            .ce0      ( buf_ce0[ 0 ] ),
            .we0      ( buf_we0[ 0 ] ),
            .d0       ( buf_d0_0 ),
            .q0       ( buf_q0_0 ),
            .address1 ( buf_a1_0 ),
            .ce1      ( buf_ce1[ 0 ] ),
            .q1       ( buf_q1_0 )
        );
        td_fused_top_dataflow_in_loop_TOP_LOOP37928_products_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP37928_products_0_memcore_U_1 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_1 ),
            .ce0      ( buf_ce0[ 1 ] ),
            .we0      ( buf_we0[ 1 ] ),
            .d0       ( buf_d0_1 ),
            .q0       ( buf_q0_1 ),
            .address1 ( buf_a1_1 ),
            .ce1      ( buf_ce1[ 1 ] ),
            .q1       ( buf_q1_1 )
        );

//++++++++++++++++++++++++buffer signals+++++++++++++++++
        assign buf_ce0[ 0 ] = (tptr ==  0  && empty_n) ? t_ce0
                             : (iptr ==  0 ) ? i_ce0 : 1'b0;
        assign buf_a0_0  = (tptr ==  0  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 0 ] = (tptr ==  0  && empty_n)  ? t_we0
                             : (iptr ==  0 ) ? i_we0 : 1'b0;
        assign buf_d0_0  = (tptr ==  0  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 0 ] = (tptr ==  0  && empty_n) ? t_ce1
                             : (iptr ==  0 ) ? i_ce1 : 1'b0;
        assign buf_a1_0  = (tptr ==  0  && empty_n) ?  t_address1 : i_address1;
        assign buf_ce0[ 1 ] = (tptr ==  1  && empty_n) ? t_ce0
                             : (iptr ==  1 ) ? i_ce0 : 1'b0;
        assign buf_a0_1  = (tptr ==  1  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 1 ] = (tptr ==  1  && empty_n)  ? t_we0
                             : (iptr ==  1 ) ? i_we0 : 1'b0;
        assign buf_d0_1  = (tptr ==  1  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 1 ] = (tptr ==  1  && empty_n) ? t_ce1
                             : (iptr ==  1 ) ? i_ce1 : 1'b0;
        assign buf_a1_1  = (tptr ==  1  && empty_n) ?  t_address1 : i_address1;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//------------------------Body---------------------------
assign i_q0      = (prev_iptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign t_q0      = reg_valid0 ? reg_q0 : (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign i_q1      = (prev_iptr == 1'b1 ? buf_q1_1 : buf_q1_0);
assign t_q1      = reg_valid1 ? reg_q1 : (prev_tptr == 1'b1 ? buf_q1_1 : buf_q1_0);

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// prev_iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_iptr <= 1'b0;
    else begin
        prev_iptr <= iptr;
    end
end

// prev_tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_tptr <= 1'b0;
    else begin
        prev_tptr <= tptr;
    end
end

// reg_q0 and reg_valid0
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q0     <= 1'b0;
        reg_valid0 <= 1'b0;
    end else if (!t_ce0 && !reg_valid0) begin
        reg_q0     <= (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
        reg_valid0 <= 1'b1;
    end else if (t_ce0) begin
        reg_valid0 <= 1'b0;
    end
end

// reg_q1 and reg_valid1
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q1     <= 1'b0;
        reg_valid1 <= 1'b0;
    end else if (!t_ce1 && !reg_valid1) begin
        reg_q1     <= (prev_tptr == 1'b1 ? buf_q1_1 : buf_q1_0);
        reg_valid1 <= 1'b1;
    end else if (t_ce1) begin
        reg_valid1 <= 1'b0;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_dataflow_in_loop_TOP_LOOP37928 (
        ap_clk,
        ap_rst,
        in_data_address0,
        in_data_ce0,
        in_data_d0,
        in_data_q0,
        in_data_we0,
        in_data_address1,
        in_data_ce1,
        in_data_d1,
        in_data_q1,
        in_data_we1,
        filter_data_address0,
        filter_data_ce0,
        filter_data_d0,
        filter_data_q0,
        filter_data_we0,
        filter_data_address1,
        filter_data_ce1,
        filter_data_d1,
        filter_data_q1,
        filter_data_we1,
        adjustments_address0,
        adjustments_ce0,
        adjustments_d0,
        adjustments_q0,
        adjustments_we0,
        adjustments_address1,
        adjustments_ce1,
        adjustments_d1,
        adjustments_q1,
        adjustments_we1,
        out_data_address0,
        out_data_ce0,
        out_data_d0,
        out_data_q0,
        out_data_we0,
        out_data_address1,
        out_data_ce1,
        out_data_d1,
        out_data_q1,
        out_data_we1,
        ap_start,
        in_data_empty_n,
        in_data_read,
        out_data_full_n,
        out_data_write,
        ap_done,
        ap_ready,
        ap_idle,
        ap_continue
);


input   ap_clk;
input   ap_rst;
output  [14:0] in_data_address0;
output   in_data_ce0;
output  [63:0] in_data_d0;
input  [63:0] in_data_q0;
output   in_data_we0;
output  [14:0] in_data_address1;
output   in_data_ce1;
output  [63:0] in_data_d1;
input  [63:0] in_data_q1;
output   in_data_we1;
output  [8:0] filter_data_address0;
output   filter_data_ce0;
output  [15:0] filter_data_d0;
input  [15:0] filter_data_q0;
output   filter_data_we0;
output  [8:0] filter_data_address1;
output   filter_data_ce1;
output  [15:0] filter_data_d1;
input  [15:0] filter_data_q1;
output   filter_data_we1;
output  [3:0] adjustments_address0;
output   adjustments_ce0;
output  [47:0] adjustments_d0;
input  [47:0] adjustments_q0;
output   adjustments_we0;
output  [3:0] adjustments_address1;
output   adjustments_ce1;
output  [47:0] adjustments_d1;
input  [47:0] adjustments_q1;
output   adjustments_we1;
output  [13:0] out_data_address0;
output   out_data_ce0;
output  [63:0] out_data_d0;
input  [63:0] out_data_q0;
output   out_data_we0;
output  [13:0] out_data_address1;
output   out_data_ce1;
output  [63:0] out_data_d1;
input  [63:0] out_data_q1;
output   out_data_we1;
input   ap_start;
input   in_data_empty_n;
output   in_data_read;
input   out_data_full_n;
output   out_data_write;
output   ap_done;
output   ap_ready;
output   ap_idle;
input   ap_continue;

wire   [15:0] ifmap_vec_0_0_i_q0;
wire   [15:0] ifmap_vec_0_0_t_q0;
wire   [15:0] weight_vecs_0_0_0_i_q0;
wire   [15:0] weight_vecs_0_0_0_t_q0;
wire   [15:0] products_0_i_q0;
wire   [15:0] products_0_i_q1;
wire   [15:0] products_0_t_q0;
wire   [15:0] products_0_t_q1;
wire   [15:0] accum1_out_0_i_q0;
wire   [15:0] accum1_out_0_t_q0;
wire    tdf3_get_next_ijk_U0_ap_start;
wire    tdf3_get_next_ijk_U0_ap_done;
wire    tdf3_get_next_ijk_U0_ap_continue;
wire    tdf3_get_next_ijk_U0_ap_idle;
wire    tdf3_get_next_ijk_U0_ap_ready;
wire    tdf3_get_next_ijk_U0_start_out;
wire    tdf3_get_next_ijk_U0_start_write;
wire   [15:0] tdf3_get_next_ijk_U0_indices_0_din;
wire    tdf3_get_next_ijk_U0_indices_0_write;
wire   [15:0] tdf3_get_next_ijk_U0_indices_1_din;
wire    tdf3_get_next_ijk_U0_indices_1_write;
wire   [3:0] tdf3_get_next_ijk_U0_indices_2_out_din;
wire    tdf3_get_next_ijk_U0_indices_2_out_write;
wire   [3:0] tdf3_get_next_ijk_U0_indices_2_out1_din;
wire    tdf3_get_next_ijk_U0_indices_2_out1_write;
wire    tdf3_readInputs_U0_ap_start;
wire    tdf3_readInputs_U0_ap_done;
wire    tdf3_readInputs_U0_ap_continue;
wire    tdf3_readInputs_U0_ap_idle;
wire    tdf3_readInputs_U0_ap_ready;
wire   [14:0] tdf3_readInputs_U0_in_data_address0;
wire    tdf3_readInputs_U0_in_data_ce0;
wire    tdf3_readInputs_U0_indices_01_read;
wire    tdf3_readInputs_U0_indices_12_read;
wire   [4:0] tdf3_readInputs_U0_ifmap_vec_0_0_address0;
wire    tdf3_readInputs_U0_ifmap_vec_0_0_ce0;
wire    tdf3_readInputs_U0_ifmap_vec_0_0_we0;
wire   [15:0] tdf3_readInputs_U0_ifmap_vec_0_0_d0;
wire   [4:0] tdf3_readInputs_U0_ifmap_vec_0_0_address1;
wire    tdf3_readInputs_U0_ifmap_vec_0_0_ce1;
wire    tdf3_readInputs_U0_ifmap_vec_0_0_we1;
wire   [15:0] tdf3_readInputs_U0_ifmap_vec_0_0_d1;
wire   [5:0] tdf3_readInputs_U0_indices_01_out_din;
wire    tdf3_readInputs_U0_indices_01_out_write;
wire   [11:0] tdf3_readInputs_U0_indices_12_out_din;
wire    tdf3_readInputs_U0_indices_12_out_write;
wire    tdf3_readInputs_U0_in_data_full_n;
wire    tdf3_readInputs_U0_in_data_write;
wire    ap_channel_done_ifmap_vec_0_0;
wire    tdf3_readInputs_U0_ifmap_vec_0_0_full_n;
wire    tdf3_readFilters30_U0_ap_start;
wire    tdf3_readFilters30_U0_ap_done;
wire    tdf3_readFilters30_U0_ap_continue;
wire    tdf3_readFilters30_U0_ap_idle;
wire    tdf3_readFilters30_U0_ap_ready;
wire   [8:0] tdf3_readFilters30_U0_filter_data_address0;
wire    tdf3_readFilters30_U0_filter_data_ce0;
wire    tdf3_readFilters30_U0_indices_23_read;
wire   [4:0] tdf3_readFilters30_U0_weight_vecs_0_0_0_address0;
wire    tdf3_readFilters30_U0_weight_vecs_0_0_0_ce0;
wire    tdf3_readFilters30_U0_weight_vecs_0_0_0_we0;
wire   [15:0] tdf3_readFilters30_U0_weight_vecs_0_0_0_d0;
wire    ap_channel_done_weight_vecs_0_0_0;
wire    tdf3_readFilters30_U0_weight_vecs_0_0_0_full_n;
wire    tdf3_dot_product_U0_ap_start;
wire    tdf3_dot_product_U0_ap_done;
wire    tdf3_dot_product_U0_ap_continue;
wire    tdf3_dot_product_U0_ap_idle;
wire    tdf3_dot_product_U0_ap_ready;
wire   [4:0] tdf3_dot_product_U0_ifmap_vec_0_0_address0;
wire    tdf3_dot_product_U0_ifmap_vec_0_0_ce0;
wire   [4:0] tdf3_dot_product_U0_weight_vecs_0_0_0_address0;
wire    tdf3_dot_product_U0_weight_vecs_0_0_0_ce0;
wire   [4:0] tdf3_dot_product_U0_products_0_address0;
wire    tdf3_dot_product_U0_products_0_ce0;
wire    tdf3_dot_product_U0_products_0_we0;
wire   [15:0] tdf3_dot_product_U0_products_0_d0;
wire    ap_channel_done_products_0;
wire    tdf3_dot_product_U0_products_0_full_n;
wire    tdf3_accum_1_U0_ap_start;
wire    tdf3_accum_1_U0_ap_done;
wire    tdf3_accum_1_U0_ap_continue;
wire    tdf3_accum_1_U0_ap_idle;
wire    tdf3_accum_1_U0_ap_ready;
wire   [4:0] tdf3_accum_1_U0_accum_in_0_address0;
wire    tdf3_accum_1_U0_accum_in_0_ce0;
wire   [4:0] tdf3_accum_1_U0_accum_in_0_address1;
wire    tdf3_accum_1_U0_accum_in_0_ce1;
wire   [2:0] tdf3_accum_1_U0_accum_out_address0;
wire    tdf3_accum_1_U0_accum_out_ce0;
wire    tdf3_accum_1_U0_accum_out_we0;
wire   [15:0] tdf3_accum_1_U0_accum_out_d0;
wire   [2:0] tdf3_accum_1_U0_accum_out_address1;
wire    tdf3_accum_1_U0_accum_out_ce1;
wire    tdf3_accum_1_U0_accum_out_we1;
wire   [15:0] tdf3_accum_1_U0_accum_out_d1;
wire    ap_channel_done_accum1_out_0;
wire    tdf3_accum_1_U0_accum_out_full_n;
wire    tdf3_accum_2_U0_ap_start;
wire    tdf3_accum_2_U0_ap_done;
wire    tdf3_accum_2_U0_ap_continue;
wire    tdf3_accum_2_U0_ap_idle;
wire    tdf3_accum_2_U0_ap_ready;
wire   [15:0] tdf3_accum_2_U0_accum_in_14;
wire    tdf3_accum_2_U0_accum_in_14_ap_vld;
wire   [2:0] tdf3_accum_2_U0_accum_in_address0;
wire    tdf3_accum_2_U0_accum_in_ce0;
wire    ap_channel_done_tmp_channel;
wire    tmp_channel_full_n;
wire    Block_entry_proc_proc397_U0_ap_start;
wire    Block_entry_proc_proc397_U0_ap_done;
wire    Block_entry_proc_proc397_U0_ap_continue;
wire    Block_entry_proc_proc397_U0_ap_idle;
wire    Block_entry_proc_proc397_U0_ap_ready;
wire   [15:0] Block_entry_proc_proc397_U0_ap_return;
wire    ap_channel_done_sums_0;
wire    sums_0_full_n;
wire    tdf3_adjust_U0_ap_start;
wire    tdf3_adjust_U0_ap_done;
wire    tdf3_adjust_U0_ap_continue;
wire    tdf3_adjust_U0_ap_idle;
wire    tdf3_adjust_U0_ap_ready;
wire   [3:0] tdf3_adjust_U0_adjustments_address0;
wire    tdf3_adjust_U0_adjustments_ce0;
wire    tdf3_adjust_U0_indices_23_read;
wire   [15:0] tdf3_adjust_U0_ap_return;
wire    ap_channel_done_outputs_0;
wire    outputs_0_full_n;
wire    tdf3_writeOutputs_unaligned_U0_ap_start;
wire    tdf3_writeOutputs_unaligned_U0_ap_done;
wire    tdf3_writeOutputs_unaligned_U0_ap_continue;
wire    tdf3_writeOutputs_unaligned_U0_ap_idle;
wire    tdf3_writeOutputs_unaligned_U0_ap_ready;
wire    tdf3_writeOutputs_unaligned_U0_indices_01_read;
wire    tdf3_writeOutputs_unaligned_U0_indices_12_read;
wire   [13:0] tdf3_writeOutputs_unaligned_U0_out_data_address1;
wire    tdf3_writeOutputs_unaligned_U0_out_data_ce1;
wire    tdf3_writeOutputs_unaligned_U0_out_data_we1;
wire   [63:0] tdf3_writeOutputs_unaligned_U0_out_data_d1;
wire    tdf3_writeOutputs_unaligned_U0_out_data_full_n;
wire    tdf3_writeOutputs_unaligned_U0_out_data_write;
wire    ap_sync_continue;
wire    ifmap_vec_0_0_i_full_n;
wire    ifmap_vec_0_0_t_empty_n;
wire    weight_vecs_0_0_0_i_full_n;
wire    weight_vecs_0_0_0_t_empty_n;
wire    products_0_i_full_n;
wire    products_0_t_empty_n;
wire   [15:0] products_0_t_d1;
wire    products_0_t_we1;
wire    accum1_out_0_i_full_n;
wire    accum1_out_0_t_empty_n;
wire    indices_01_c_full_n;
wire   [15:0] indices_01_c_dout;
wire    indices_01_c_empty_n;
wire    indices_12_c_full_n;
wire   [15:0] indices_12_c_dout;
wire    indices_12_c_empty_n;
wire    indices_23_c_full_n;
wire   [3:0] indices_23_c_dout;
wire    indices_23_c_empty_n;
wire    indices_23_c1_full_n;
wire   [3:0] indices_23_c1_dout;
wire    indices_23_c1_empty_n;
wire    indices_01_c2_full_n;
wire   [5:0] indices_01_c2_dout;
wire    indices_01_c2_empty_n;
wire    indices_12_c3_full_n;
wire   [11:0] indices_12_c3_dout;
wire    indices_12_c3_empty_n;
wire   [15:0] tmp_channel_dout;
wire    tmp_channel_empty_n;
wire   [15:0] sums_0_dout;
wire    sums_0_empty_n;
wire   [15:0] outputs_0_dout;
wire    outputs_0_empty_n;
wire    ap_sync_done;
wire    ap_sync_ready;
reg    ap_sync_reg_tdf3_get_next_ijk_U0_ap_ready;
wire    ap_sync_tdf3_get_next_ijk_U0_ap_ready;
reg    ap_sync_reg_tdf3_readInputs_U0_ap_ready;
wire    ap_sync_tdf3_readInputs_U0_ap_ready;
wire   [0:0] start_for_tdf3_readFilters30_U0_din;
wire    start_for_tdf3_readFilters30_U0_full_n;
wire   [0:0] start_for_tdf3_readFilters30_U0_dout;
wire    start_for_tdf3_readFilters30_U0_empty_n;
wire    tdf3_readInputs_U0_start_full_n;
wire    tdf3_readInputs_U0_start_write;
wire    tdf3_readFilters30_U0_start_full_n;
wire    tdf3_readFilters30_U0_start_write;
wire    tdf3_dot_product_U0_start_full_n;
wire    tdf3_dot_product_U0_start_write;
wire    tdf3_accum_1_U0_start_full_n;
wire    tdf3_accum_1_U0_start_write;
wire    tdf3_accum_2_U0_start_full_n;
wire    tdf3_accum_2_U0_start_write;
wire    Block_entry_proc_proc397_U0_start_full_n;
wire    Block_entry_proc_proc397_U0_start_write;
wire    tdf3_adjust_U0_start_full_n;
wire    tdf3_adjust_U0_start_write;
wire    tdf3_writeOutputs_unaligned_U0_start_full_n;
wire    tdf3_writeOutputs_unaligned_U0_start_write;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_sync_reg_tdf3_get_next_ijk_U0_ap_ready = 1'b0;
#0 ap_sync_reg_tdf3_readInputs_U0_ap_ready = 1'b0;
end

td_fused_top_dataflow_in_loop_TOP_LOOP37928_ifmap_vec_0_0 #(
    .DataWidth( 16 ),
    .AddressRange( 32 ),
    .AddressWidth( 5 ))
ifmap_vec_0_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf3_readInputs_U0_ap_done),
    .i_full_n(ifmap_vec_0_0_i_full_n),
    .i_ce0(tdf3_readInputs_U0_ifmap_vec_0_0_ce0),
    .i_we0(tdf3_readInputs_U0_ifmap_vec_0_0_we0),
    .i_address0(tdf3_readInputs_U0_ifmap_vec_0_0_address0),
    .i_d0(tdf3_readInputs_U0_ifmap_vec_0_0_d0),
    .i_q0(ifmap_vec_0_0_i_q0),
    .i_ce1(tdf3_readInputs_U0_ifmap_vec_0_0_ce1),
    .i_we1(tdf3_readInputs_U0_ifmap_vec_0_0_we1),
    .i_address1(tdf3_readInputs_U0_ifmap_vec_0_0_address1),
    .i_d1(tdf3_readInputs_U0_ifmap_vec_0_0_d1),
    .t_ce(1'b1),
    .t_read(tdf3_dot_product_U0_ap_ready),
    .t_empty_n(ifmap_vec_0_0_t_empty_n),
    .t_ce0(tdf3_dot_product_U0_ifmap_vec_0_0_ce0),
    .t_we0(1'b0),
    .t_address0(tdf3_dot_product_U0_ifmap_vec_0_0_address0),
    .t_d0(16'd0),
    .t_q0(ifmap_vec_0_0_t_q0),
    .t_ce1(1'b0),
    .t_we1(1'b0),
    .t_address1(5'd0),
    .t_d1(16'd0)
);

td_fused_top_dataflow_in_loop_TOP_LOOP37928_weight_vecs_0_0_0 #(
    .DataWidth( 16 ),
    .AddressRange( 32 ),
    .AddressWidth( 5 ))
weight_vecs_0_0_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf3_readFilters30_U0_ap_done),
    .i_full_n(weight_vecs_0_0_0_i_full_n),
    .i_ce0(tdf3_readFilters30_U0_weight_vecs_0_0_0_ce0),
    .i_we0(tdf3_readFilters30_U0_weight_vecs_0_0_0_we0),
    .i_address0(tdf3_readFilters30_U0_weight_vecs_0_0_0_address0),
    .i_d0(tdf3_readFilters30_U0_weight_vecs_0_0_0_d0),
    .i_q0(weight_vecs_0_0_0_i_q0),
    .t_ce(1'b1),
    .t_read(tdf3_dot_product_U0_ap_ready),
    .t_empty_n(weight_vecs_0_0_0_t_empty_n),
    .t_ce0(tdf3_dot_product_U0_weight_vecs_0_0_0_ce0),
    .t_we0(1'b0),
    .t_address0(tdf3_dot_product_U0_weight_vecs_0_0_0_address0),
    .t_d0(16'd0),
    .t_q0(weight_vecs_0_0_0_t_q0)
);

td_fused_top_dataflow_in_loop_TOP_LOOP37928_products_0 #(
    .DataWidth( 16 ),
    .AddressRange( 32 ),
    .AddressWidth( 5 ))
products_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf3_dot_product_U0_ap_done),
    .i_full_n(products_0_i_full_n),
    .i_ce0(tdf3_dot_product_U0_products_0_ce0),
    .i_we0(tdf3_dot_product_U0_products_0_we0),
    .i_address0(tdf3_dot_product_U0_products_0_address0),
    .i_d0(tdf3_dot_product_U0_products_0_d0),
    .i_q0(products_0_i_q0),
    .i_ce1(1'b0),
    .i_address1(5'd0),
    .i_q1(products_0_i_q1),
    .t_ce(1'b1),
    .t_read(tdf3_accum_1_U0_ap_ready),
    .t_empty_n(products_0_t_empty_n),
    .t_ce0(tdf3_accum_1_U0_accum_in_0_ce0),
    .t_we0(1'b0),
    .t_address0(tdf3_accum_1_U0_accum_in_0_address0),
    .t_d0(16'd0),
    .t_q0(products_0_t_q0),
    .t_ce1(tdf3_accum_1_U0_accum_in_0_ce1),
    .t_address1(tdf3_accum_1_U0_accum_in_0_address1),
    .t_q1(products_0_t_q1)
);

td_fused_top_dataflow_in_loop_TOP_LOOP37928_accum1_out_0 #(
    .DataWidth( 16 ),
    .AddressRange( 8 ),
    .AddressWidth( 3 ))
accum1_out_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf3_accum_1_U0_ap_done),
    .i_full_n(accum1_out_0_i_full_n),
    .i_ce0(tdf3_accum_1_U0_accum_out_ce0),
    .i_we0(tdf3_accum_1_U0_accum_out_we0),
    .i_address0(tdf3_accum_1_U0_accum_out_address0),
    .i_d0(tdf3_accum_1_U0_accum_out_d0),
    .i_q0(accum1_out_0_i_q0),
    .i_ce1(tdf3_accum_1_U0_accum_out_ce1),
    .i_we1(tdf3_accum_1_U0_accum_out_we1),
    .i_address1(tdf3_accum_1_U0_accum_out_address1),
    .i_d1(tdf3_accum_1_U0_accum_out_d1),
    .t_ce(1'b1),
    .t_read(tdf3_accum_2_U0_ap_ready),
    .t_empty_n(accum1_out_0_t_empty_n),
    .t_ce0(tdf3_accum_2_U0_accum_in_ce0),
    .t_we0(1'b0),
    .t_address0(tdf3_accum_2_U0_accum_in_address0),
    .t_d0(16'd0),
    .t_q0(accum1_out_0_t_q0),
    .t_ce1(1'b0),
    .t_we1(1'b0),
    .t_address1(3'd0),
    .t_d1(16'd0)
);

td_fused_top_tdf3_get_next_ijk tdf3_get_next_ijk_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf3_get_next_ijk_U0_ap_start),
    .start_full_n(start_for_tdf3_readFilters30_U0_full_n),
    .ap_done(tdf3_get_next_ijk_U0_ap_done),
    .ap_continue(tdf3_get_next_ijk_U0_ap_continue),
    .ap_idle(tdf3_get_next_ijk_U0_ap_idle),
    .ap_ready(tdf3_get_next_ijk_U0_ap_ready),
    .start_out(tdf3_get_next_ijk_U0_start_out),
    .start_write(tdf3_get_next_ijk_U0_start_write),
    .indices_0_din(tdf3_get_next_ijk_U0_indices_0_din),
    .indices_0_full_n(indices_01_c_full_n),
    .indices_0_write(tdf3_get_next_ijk_U0_indices_0_write),
    .indices_1_din(tdf3_get_next_ijk_U0_indices_1_din),
    .indices_1_full_n(indices_12_c_full_n),
    .indices_1_write(tdf3_get_next_ijk_U0_indices_1_write),
    .indices_2_out_din(tdf3_get_next_ijk_U0_indices_2_out_din),
    .indices_2_out_full_n(indices_23_c_full_n),
    .indices_2_out_write(tdf3_get_next_ijk_U0_indices_2_out_write),
    .indices_2_out1_din(tdf3_get_next_ijk_U0_indices_2_out1_din),
    .indices_2_out1_full_n(indices_23_c1_full_n),
    .indices_2_out1_write(tdf3_get_next_ijk_U0_indices_2_out1_write)
);

td_fused_top_tdf3_readInputs tdf3_readInputs_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf3_readInputs_U0_ap_start),
    .ap_done(tdf3_readInputs_U0_ap_done),
    .ap_continue(tdf3_readInputs_U0_ap_continue),
    .ap_idle(tdf3_readInputs_U0_ap_idle),
    .ap_ready(tdf3_readInputs_U0_ap_ready),
    .in_data_address0(tdf3_readInputs_U0_in_data_address0),
    .in_data_ce0(tdf3_readInputs_U0_in_data_ce0),
    .in_data_q0(in_data_q0),
    .indices_01_dout(indices_01_c_dout),
    .indices_01_empty_n(indices_01_c_empty_n),
    .indices_01_read(tdf3_readInputs_U0_indices_01_read),
    .indices_12_dout(indices_12_c_dout),
    .indices_12_empty_n(indices_12_c_empty_n),
    .indices_12_read(tdf3_readInputs_U0_indices_12_read),
    .ifmap_vec_0_0_address0(tdf3_readInputs_U0_ifmap_vec_0_0_address0),
    .ifmap_vec_0_0_ce0(tdf3_readInputs_U0_ifmap_vec_0_0_ce0),
    .ifmap_vec_0_0_we0(tdf3_readInputs_U0_ifmap_vec_0_0_we0),
    .ifmap_vec_0_0_d0(tdf3_readInputs_U0_ifmap_vec_0_0_d0),
    .ifmap_vec_0_0_address1(tdf3_readInputs_U0_ifmap_vec_0_0_address1),
    .ifmap_vec_0_0_ce1(tdf3_readInputs_U0_ifmap_vec_0_0_ce1),
    .ifmap_vec_0_0_we1(tdf3_readInputs_U0_ifmap_vec_0_0_we1),
    .ifmap_vec_0_0_d1(tdf3_readInputs_U0_ifmap_vec_0_0_d1),
    .indices_01_out_din(tdf3_readInputs_U0_indices_01_out_din),
    .indices_01_out_full_n(indices_01_c2_full_n),
    .indices_01_out_write(tdf3_readInputs_U0_indices_01_out_write),
    .indices_12_out_din(tdf3_readInputs_U0_indices_12_out_din),
    .indices_12_out_full_n(indices_12_c3_full_n),
    .indices_12_out_write(tdf3_readInputs_U0_indices_12_out_write)
);

td_fused_top_tdf3_readFilters30 tdf3_readFilters30_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf3_readFilters30_U0_ap_start),
    .ap_done(tdf3_readFilters30_U0_ap_done),
    .ap_continue(tdf3_readFilters30_U0_ap_continue),
    .ap_idle(tdf3_readFilters30_U0_ap_idle),
    .ap_ready(tdf3_readFilters30_U0_ap_ready),
    .filter_data_address0(tdf3_readFilters30_U0_filter_data_address0),
    .filter_data_ce0(tdf3_readFilters30_U0_filter_data_ce0),
    .filter_data_q0(filter_data_q0),
    .indices_23_dout(indices_23_c_dout),
    .indices_23_empty_n(indices_23_c_empty_n),
    .indices_23_read(tdf3_readFilters30_U0_indices_23_read),
    .weight_vecs_0_0_0_address0(tdf3_readFilters30_U0_weight_vecs_0_0_0_address0),
    .weight_vecs_0_0_0_ce0(tdf3_readFilters30_U0_weight_vecs_0_0_0_ce0),
    .weight_vecs_0_0_0_we0(tdf3_readFilters30_U0_weight_vecs_0_0_0_we0),
    .weight_vecs_0_0_0_d0(tdf3_readFilters30_U0_weight_vecs_0_0_0_d0)
);

td_fused_top_tdf3_dot_product tdf3_dot_product_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf3_dot_product_U0_ap_start),
    .ap_done(tdf3_dot_product_U0_ap_done),
    .ap_continue(tdf3_dot_product_U0_ap_continue),
    .ap_idle(tdf3_dot_product_U0_ap_idle),
    .ap_ready(tdf3_dot_product_U0_ap_ready),
    .ifmap_vec_0_0_address0(tdf3_dot_product_U0_ifmap_vec_0_0_address0),
    .ifmap_vec_0_0_ce0(tdf3_dot_product_U0_ifmap_vec_0_0_ce0),
    .ifmap_vec_0_0_q0(ifmap_vec_0_0_t_q0),
    .weight_vecs_0_0_0_address0(tdf3_dot_product_U0_weight_vecs_0_0_0_address0),
    .weight_vecs_0_0_0_ce0(tdf3_dot_product_U0_weight_vecs_0_0_0_ce0),
    .weight_vecs_0_0_0_q0(weight_vecs_0_0_0_t_q0),
    .products_0_address0(tdf3_dot_product_U0_products_0_address0),
    .products_0_ce0(tdf3_dot_product_U0_products_0_ce0),
    .products_0_we0(tdf3_dot_product_U0_products_0_we0),
    .products_0_d0(tdf3_dot_product_U0_products_0_d0)
);

td_fused_top_tdf3_accum_1 tdf3_accum_1_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf3_accum_1_U0_ap_start),
    .ap_done(tdf3_accum_1_U0_ap_done),
    .ap_continue(tdf3_accum_1_U0_ap_continue),
    .ap_idle(tdf3_accum_1_U0_ap_idle),
    .ap_ready(tdf3_accum_1_U0_ap_ready),
    .accum_in_0_address0(tdf3_accum_1_U0_accum_in_0_address0),
    .accum_in_0_ce0(tdf3_accum_1_U0_accum_in_0_ce0),
    .accum_in_0_q0(products_0_t_q0),
    .accum_in_0_address1(tdf3_accum_1_U0_accum_in_0_address1),
    .accum_in_0_ce1(tdf3_accum_1_U0_accum_in_0_ce1),
    .accum_in_0_q1(products_0_t_q1),
    .accum_out_address0(tdf3_accum_1_U0_accum_out_address0),
    .accum_out_ce0(tdf3_accum_1_U0_accum_out_ce0),
    .accum_out_we0(tdf3_accum_1_U0_accum_out_we0),
    .accum_out_d0(tdf3_accum_1_U0_accum_out_d0),
    .accum_out_address1(tdf3_accum_1_U0_accum_out_address1),
    .accum_out_ce1(tdf3_accum_1_U0_accum_out_ce1),
    .accum_out_we1(tdf3_accum_1_U0_accum_out_we1),
    .accum_out_d1(tdf3_accum_1_U0_accum_out_d1)
);

td_fused_top_tdf3_accum_2 tdf3_accum_2_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf3_accum_2_U0_ap_start),
    .ap_done(tdf3_accum_2_U0_ap_done),
    .ap_continue(tdf3_accum_2_U0_ap_continue),
    .ap_idle(tdf3_accum_2_U0_ap_idle),
    .ap_ready(tdf3_accum_2_U0_ap_ready),
    .accum_in_14(tdf3_accum_2_U0_accum_in_14),
    .accum_in_14_ap_vld(tdf3_accum_2_U0_accum_in_14_ap_vld),
    .accum_in_address0(tdf3_accum_2_U0_accum_in_address0),
    .accum_in_ce0(tdf3_accum_2_U0_accum_in_ce0),
    .accum_in_q0(accum1_out_0_t_q0)
);

td_fused_top_Block_entry_proc_proc397 Block_entry_proc_proc397_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(Block_entry_proc_proc397_U0_ap_start),
    .ap_done(Block_entry_proc_proc397_U0_ap_done),
    .ap_continue(Block_entry_proc_proc397_U0_ap_continue),
    .ap_idle(Block_entry_proc_proc397_U0_ap_idle),
    .ap_ready(Block_entry_proc_proc397_U0_ap_ready),
    .tmp(tmp_channel_dout),
    .ap_return(Block_entry_proc_proc397_U0_ap_return)
);

td_fused_top_tdf3_adjust tdf3_adjust_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf3_adjust_U0_ap_start),
    .ap_done(tdf3_adjust_U0_ap_done),
    .ap_continue(tdf3_adjust_U0_ap_continue),
    .ap_idle(tdf3_adjust_U0_ap_idle),
    .ap_ready(tdf3_adjust_U0_ap_ready),
    .sums_read(sums_0_dout),
    .adjustments_address0(tdf3_adjust_U0_adjustments_address0),
    .adjustments_ce0(tdf3_adjust_U0_adjustments_ce0),
    .adjustments_q0(adjustments_q0),
    .indices_23_dout(indices_23_c1_dout),
    .indices_23_empty_n(indices_23_c1_empty_n),
    .indices_23_read(tdf3_adjust_U0_indices_23_read),
    .ap_return(tdf3_adjust_U0_ap_return)
);

td_fused_top_tdf3_writeOutputs_unaligned tdf3_writeOutputs_unaligned_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf3_writeOutputs_unaligned_U0_ap_start),
    .ap_done(tdf3_writeOutputs_unaligned_U0_ap_done),
    .ap_continue(tdf3_writeOutputs_unaligned_U0_ap_continue),
    .ap_idle(tdf3_writeOutputs_unaligned_U0_ap_idle),
    .ap_ready(tdf3_writeOutputs_unaligned_U0_ap_ready),
    .indices_01_dout(indices_01_c2_dout),
    .indices_01_empty_n(indices_01_c2_empty_n),
    .indices_01_read(tdf3_writeOutputs_unaligned_U0_indices_01_read),
    .indices_12_dout(indices_12_c3_dout),
    .indices_12_empty_n(indices_12_c3_empty_n),
    .indices_12_read(tdf3_writeOutputs_unaligned_U0_indices_12_read),
    .p_read(outputs_0_dout),
    .out_data_address1(tdf3_writeOutputs_unaligned_U0_out_data_address1),
    .out_data_ce1(tdf3_writeOutputs_unaligned_U0_out_data_ce1),
    .out_data_we1(tdf3_writeOutputs_unaligned_U0_out_data_we1),
    .out_data_d1(tdf3_writeOutputs_unaligned_U0_out_data_d1)
);

td_fused_top_fifo_w16_d2_S_x0 indices_01_c_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(indices_01_c_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf3_readInputs_U0_indices_01_read),
    .if_dout(indices_01_c_dout),
    .if_full_n(indices_01_c_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf3_get_next_ijk_U0_indices_0_write),
    .if_din(tdf3_get_next_ijk_U0_indices_0_din)
);

td_fused_top_fifo_w16_d2_S_x0 indices_12_c_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(indices_12_c_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf3_readInputs_U0_indices_12_read),
    .if_dout(indices_12_c_dout),
    .if_full_n(indices_12_c_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf3_get_next_ijk_U0_indices_1_write),
    .if_din(tdf3_get_next_ijk_U0_indices_1_din)
);

td_fused_top_fifo_w4_d2_S_x indices_23_c_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(indices_23_c_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf3_readFilters30_U0_indices_23_read),
    .if_dout(indices_23_c_dout),
    .if_full_n(indices_23_c_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf3_get_next_ijk_U0_indices_2_out_write),
    .if_din(tdf3_get_next_ijk_U0_indices_2_out_din)
);

td_fused_top_fifo_w4_d7_S indices_23_c1_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(indices_23_c1_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf3_adjust_U0_indices_23_read),
    .if_dout(indices_23_c1_dout),
    .if_full_n(indices_23_c1_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf3_get_next_ijk_U0_indices_2_out1_write),
    .if_din(tdf3_get_next_ijk_U0_indices_2_out1_din)
);

td_fused_top_fifo_w6_d7_S indices_01_c2_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(indices_01_c2_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf3_writeOutputs_unaligned_U0_indices_01_read),
    .if_dout(indices_01_c2_dout),
    .if_full_n(indices_01_c2_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf3_readInputs_U0_indices_01_out_write),
    .if_din(tdf3_readInputs_U0_indices_01_out_din)
);

td_fused_top_fifo_w12_d7_S indices_12_c3_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(indices_12_c3_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf3_writeOutputs_unaligned_U0_indices_12_read),
    .if_dout(indices_12_c3_dout),
    .if_full_n(indices_12_c3_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf3_readInputs_U0_indices_12_out_write),
    .if_din(tdf3_readInputs_U0_indices_12_out_din)
);

td_fused_top_fifo_w16_d2_S_x0 tmp_channel_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(tmp_channel_empty_n),
    .if_read_ce(1'b1),
    .if_read(Block_entry_proc_proc397_U0_ap_ready),
    .if_dout(tmp_channel_dout),
    .if_full_n(tmp_channel_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf3_accum_2_U0_ap_done),
    .if_din(tdf3_accum_2_U0_accum_in_14)
);

td_fused_top_fifo_w16_d2_S_x0 sums_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(sums_0_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf3_adjust_U0_ap_ready),
    .if_dout(sums_0_dout),
    .if_full_n(sums_0_full_n),
    .if_write_ce(1'b1),
    .if_write(Block_entry_proc_proc397_U0_ap_done),
    .if_din(Block_entry_proc_proc397_U0_ap_return)
);

td_fused_top_fifo_w16_d2_S_x0 outputs_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(outputs_0_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf3_writeOutputs_unaligned_U0_ap_ready),
    .if_dout(outputs_0_dout),
    .if_full_n(outputs_0_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf3_adjust_U0_ap_done),
    .if_din(tdf3_adjust_U0_ap_return)
);

td_fused_top_start_for_tdf3_readFilters30_U0 start_for_tdf3_readFilters30_U0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(start_for_tdf3_readFilters30_U0_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf3_readFilters30_U0_ap_ready),
    .if_dout(start_for_tdf3_readFilters30_U0_dout),
    .if_full_n(start_for_tdf3_readFilters30_U0_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf3_get_next_ijk_U0_start_write),
    .if_din(start_for_tdf3_readFilters30_U0_din)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_sync_reg_tdf3_get_next_ijk_U0_ap_ready <= 1'b0;
    end else begin
        if (((ap_sync_ready & ap_start) == 1'b1)) begin
            ap_sync_reg_tdf3_get_next_ijk_U0_ap_ready <= 1'b0;
        end else begin
            ap_sync_reg_tdf3_get_next_ijk_U0_ap_ready <= ap_sync_tdf3_get_next_ijk_U0_ap_ready;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_sync_reg_tdf3_readInputs_U0_ap_ready <= 1'b0;
    end else begin
        if (((ap_sync_ready & ap_start) == 1'b1)) begin
            ap_sync_reg_tdf3_readInputs_U0_ap_ready <= 1'b0;
        end else begin
            ap_sync_reg_tdf3_readInputs_U0_ap_ready <= ap_sync_tdf3_readInputs_U0_ap_ready;
        end
    end
end

assign Block_entry_proc_proc397_U0_ap_continue = sums_0_full_n;

assign Block_entry_proc_proc397_U0_ap_start = tmp_channel_empty_n;

assign Block_entry_proc_proc397_U0_start_full_n = 1'b1;

assign Block_entry_proc_proc397_U0_start_write = 1'b0;

assign adjustments_address0 = tdf3_adjust_U0_adjustments_address0;

assign adjustments_address1 = 4'd0;

assign adjustments_ce0 = tdf3_adjust_U0_adjustments_ce0;

assign adjustments_ce1 = 1'b0;

assign adjustments_d0 = 48'd0;

assign adjustments_d1 = 48'd0;

assign adjustments_we0 = 1'b0;

assign adjustments_we1 = 1'b0;

assign ap_channel_done_accum1_out_0 = tdf3_accum_1_U0_ap_done;

assign ap_channel_done_ifmap_vec_0_0 = tdf3_readInputs_U0_ap_done;

assign ap_channel_done_outputs_0 = tdf3_adjust_U0_ap_done;

assign ap_channel_done_products_0 = tdf3_dot_product_U0_ap_done;

assign ap_channel_done_sums_0 = Block_entry_proc_proc397_U0_ap_done;

assign ap_channel_done_tmp_channel = tdf3_accum_2_U0_ap_done;

assign ap_channel_done_weight_vecs_0_0_0 = tdf3_readFilters30_U0_ap_done;

assign ap_done = tdf3_writeOutputs_unaligned_U0_ap_done;

assign ap_idle = (tdf3_writeOutputs_unaligned_U0_ap_idle & tdf3_readInputs_U0_ap_idle & tdf3_readFilters30_U0_ap_idle & tdf3_get_next_ijk_U0_ap_idle & tdf3_dot_product_U0_ap_idle & tdf3_adjust_U0_ap_idle & tdf3_accum_2_U0_ap_idle & tdf3_accum_1_U0_ap_idle & (outputs_0_empty_n ^ 1'b1) & (sums_0_empty_n ^ 1'b1) & (tmp_channel_empty_n ^ 1'b1) & (products_0_t_empty_n ^ 1'b1) & (weight_vecs_0_0_0_t_empty_n ^ 1'b1) & (ifmap_vec_0_0_t_empty_n ^ 1'b1) & (1'b1 ^ accum1_out_0_t_empty_n) & Block_entry_proc_proc397_U0_ap_idle);

assign ap_ready = ap_sync_ready;

assign ap_sync_continue = ap_continue;

assign ap_sync_done = tdf3_writeOutputs_unaligned_U0_ap_done;

assign ap_sync_ready = (ap_sync_tdf3_readInputs_U0_ap_ready & ap_sync_tdf3_get_next_ijk_U0_ap_ready);

assign ap_sync_tdf3_get_next_ijk_U0_ap_ready = (tdf3_get_next_ijk_U0_ap_ready | ap_sync_reg_tdf3_get_next_ijk_U0_ap_ready);

assign ap_sync_tdf3_readInputs_U0_ap_ready = (tdf3_readInputs_U0_ap_ready | ap_sync_reg_tdf3_readInputs_U0_ap_ready);

assign filter_data_address0 = tdf3_readFilters30_U0_filter_data_address0;

assign filter_data_address1 = 9'd0;

assign filter_data_ce0 = tdf3_readFilters30_U0_filter_data_ce0;

assign filter_data_ce1 = 1'b0;

assign filter_data_d0 = 16'd0;

assign filter_data_d1 = 16'd0;

assign filter_data_we0 = 1'b0;

assign filter_data_we1 = 1'b0;

assign in_data_address0 = tdf3_readInputs_U0_in_data_address0;

assign in_data_address1 = 15'd0;

assign in_data_ce0 = tdf3_readInputs_U0_in_data_ce0;

assign in_data_ce1 = 1'b0;

assign in_data_d0 = 64'd0;

assign in_data_d1 = 64'd0;

assign in_data_read = tdf3_readInputs_U0_in_data_write;

assign in_data_we0 = 1'b0;

assign in_data_we1 = 1'b0;

assign out_data_address0 = 14'd0;

assign out_data_address1 = tdf3_writeOutputs_unaligned_U0_out_data_address1;

assign out_data_ce0 = 1'b0;

assign out_data_ce1 = tdf3_writeOutputs_unaligned_U0_out_data_ce1;

assign out_data_d0 = 64'd0;

assign out_data_d1 = tdf3_writeOutputs_unaligned_U0_out_data_d1;

assign out_data_we0 = 1'b0;

assign out_data_we1 = tdf3_writeOutputs_unaligned_U0_out_data_we1;

assign out_data_write = tdf3_writeOutputs_unaligned_U0_out_data_write;

assign products_0_t_d1 = 16'd0;

assign products_0_t_we1 = 1'b0;

assign start_for_tdf3_readFilters30_U0_din = 1'b1;

assign tdf3_accum_1_U0_accum_out_full_n = accum1_out_0_i_full_n;

assign tdf3_accum_1_U0_ap_continue = accum1_out_0_i_full_n;

assign tdf3_accum_1_U0_ap_start = products_0_t_empty_n;

assign tdf3_accum_1_U0_start_full_n = 1'b1;

assign tdf3_accum_1_U0_start_write = 1'b0;

assign tdf3_accum_2_U0_ap_continue = tmp_channel_full_n;

assign tdf3_accum_2_U0_ap_start = accum1_out_0_t_empty_n;

assign tdf3_accum_2_U0_start_full_n = 1'b1;

assign tdf3_accum_2_U0_start_write = 1'b0;

assign tdf3_adjust_U0_ap_continue = outputs_0_full_n;

assign tdf3_adjust_U0_ap_start = sums_0_empty_n;

assign tdf3_adjust_U0_start_full_n = 1'b1;

assign tdf3_adjust_U0_start_write = 1'b0;

assign tdf3_dot_product_U0_ap_continue = products_0_i_full_n;

assign tdf3_dot_product_U0_ap_start = (weight_vecs_0_0_0_t_empty_n & ifmap_vec_0_0_t_empty_n);

assign tdf3_dot_product_U0_products_0_full_n = products_0_i_full_n;

assign tdf3_dot_product_U0_start_full_n = 1'b1;

assign tdf3_dot_product_U0_start_write = 1'b0;

assign tdf3_get_next_ijk_U0_ap_continue = 1'b1;

assign tdf3_get_next_ijk_U0_ap_start = ((ap_sync_reg_tdf3_get_next_ijk_U0_ap_ready ^ 1'b1) & ap_start);

assign tdf3_readFilters30_U0_ap_continue = weight_vecs_0_0_0_i_full_n;

assign tdf3_readFilters30_U0_ap_start = start_for_tdf3_readFilters30_U0_empty_n;

assign tdf3_readFilters30_U0_start_full_n = 1'b1;

assign tdf3_readFilters30_U0_start_write = 1'b0;

assign tdf3_readFilters30_U0_weight_vecs_0_0_0_full_n = weight_vecs_0_0_0_i_full_n;

assign tdf3_readInputs_U0_ap_continue = ifmap_vec_0_0_i_full_n;

assign tdf3_readInputs_U0_ap_start = ((ap_sync_reg_tdf3_readInputs_U0_ap_ready ^ 1'b1) & ap_start);

assign tdf3_readInputs_U0_ifmap_vec_0_0_full_n = ifmap_vec_0_0_i_full_n;

assign tdf3_readInputs_U0_in_data_full_n = in_data_empty_n;

assign tdf3_readInputs_U0_in_data_write = 1'b0;

assign tdf3_readInputs_U0_start_full_n = 1'b1;

assign tdf3_readInputs_U0_start_write = 1'b0;

assign tdf3_writeOutputs_unaligned_U0_ap_continue = ap_continue;

assign tdf3_writeOutputs_unaligned_U0_ap_start = outputs_0_empty_n;

assign tdf3_writeOutputs_unaligned_U0_out_data_full_n = out_data_full_n;

assign tdf3_writeOutputs_unaligned_U0_out_data_write = 1'b0;

assign tdf3_writeOutputs_unaligned_U0_start_full_n = 1'b1;

assign tdf3_writeOutputs_unaligned_U0_start_write = 1'b0;

endmodule //td_fused_top_dataflow_in_loop_TOP_LOOP37928
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37928_weight_vecs_0_0_0_memcore_ram (addr0, ce0, d0, we0, q0, addr1, ce1, d1, we1, q1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
output reg[DWIDTH-1:0] q1;
input clk;

reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];




always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1) 
            ram[addr1] <= d1; 
        q1 <= ram[addr1];
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP37928_weight_vecs_0_0_0_memcore(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    q0,
    address1,
    ce1,
    we1,
    d1,
    q1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;
output[DataWidth - 1:0] q1;



td_fused_top_dataflow_in_loop_TOP_LOOP37928_weight_vecs_0_0_0_memcore_ram td_fused_top_dataflow_in_loop_TOP_LOOP37928_weight_vecs_0_0_0_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 ),
    .q1( q1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_dataflow_in_loop_TOP_LOOP37928_weight_vecs_0_0_0
#(parameter
    DataWidth    = 16,
    AddressRange = 32,
    AddressWidth = 5,
    BufferCount  = 2,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire                    i_we0,
    input  wire [AddressWidth-1:0] i_address0,
    input  wire [DataWidth-1:0]    i_d0,
    output wire [DataWidth-1:0]    i_q0,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire                    t_we0,
    input  wire [AddressWidth-1:0] t_address0,
    input  wire [DataWidth-1:0]    t_d0,
    output wire [DataWidth-1:0]    t_q0
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
wire [AddressWidth+IndexWidth-1:0]   memcore_iaddr;
wire [AddressWidth+IndexWidth-1:0]   memcore_taddr;

//------------------------Instantiation------------------
assign memcore_iaddr = {i_address0, iptr};
assign memcore_taddr = {t_address0, tptr};
td_fused_top_dataflow_in_loop_TOP_LOOP37928_weight_vecs_0_0_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP37928_weight_vecs_0_0_0_memcore_U (
    .reset    ( reset ),
    .clk      ( clk ),
    .address0 ( memcore_iaddr ),
    .ce0      ( i_ce0 ),
    .we0      ( i_we0),
    .d0       ( i_d0 ),
    .q0       ( i_q0 ),
    .address1 ( memcore_taddr ),
    .ce1      ( t_ce0 ),
    .we1      ( t_we0),
    .d1       ( t_d0 ),
    .q1       ( t_q0 )

);

//------------------------Body---------------------------

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP38022_accum1_out_0_memcore_ram (addr0, ce0, d0, we0, q0, addr1, ce1, d1, we1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 3;
parameter MEM_SIZE = 8;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
input clk;

reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];




always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1) 
            ram[addr1] <= d1; 
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP38022_accum1_out_0_memcore(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    q0,
    address1,
    ce1,
    we1,
    d1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd8;
parameter AddressWidth = 32'd3;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;



td_fused_top_dataflow_in_loop_TOP_LOOP38022_accum1_out_0_memcore_ram td_fused_top_dataflow_in_loop_TOP_LOOP38022_accum1_out_0_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_dataflow_in_loop_TOP_LOOP38022_accum1_out_0
#(parameter
    DataWidth    = 16,
    AddressRange = 32,
    AddressWidth = 3,
    BufferCount  = 2,
    MemLatency   = 1,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire                    i_we0,
    input  wire [AddressWidth-1:0] i_address0,
    input  wire [DataWidth-1:0]    i_d0,
    output wire [DataWidth-1:0]    i_q0,
    input  wire                    i_ce1,
    input  wire                    i_we1,
    input  wire [AddressWidth-1:0] i_address1,
    input  wire [DataWidth-1:0]    i_d1,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire                    t_we0,
    input  wire [AddressWidth-1:0] t_address0,
    input  wire [DataWidth-1:0]    t_d0,
    output wire [DataWidth-1:0]    t_q0,
    input  wire                    t_ce1,
    input  wire                    t_we1,
    input  wire [AddressWidth-1:0] t_address1,
    input  wire [DataWidth-1:0]    t_d1
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth-1:0]   prev_iptr    = 1'b0; // previous initiator index
reg  [IndexWidth-1:0]   prev_tptr    = 1'b0; // previous target index
reg  [DataWidth-1:0]    reg_q0      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid0    = 1'b0; // buffer has valid data
reg  [DataWidth-1:0]    reg_q1      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid1    = 1'b0; // buffer has valid data
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
// buffer signals
wire [BufferCount-1:0] buf_ce0;
wire [BufferCount-1:0] buf_we0;
wire [AddressWidth-1:0] buf_a0_0, buf_a0_1;
wire [DataWidth-1:0] buf_d0_0, buf_d0_1;
wire [DataWidth-1:0] buf_q0_0, buf_q0_1;
wire [BufferCount-1:0] buf_ce1;
wire [BufferCount-1:0] buf_we1;
wire [AddressWidth-1:0] buf_a1_0, buf_a1_1;
wire [DataWidth-1:0] buf_d1_0, buf_d1_1;
//------------------------Instantiation------------------
//genvar i;
        td_fused_top_dataflow_in_loop_TOP_LOOP38022_accum1_out_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP38022_accum1_out_0_memcore_U_0 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_0 ),
            .ce0      ( buf_ce0[ 0 ] ),
            .we0      ( buf_we0[ 0 ] ),
            .d0       ( buf_d0_0 ),
            .q0       ( buf_q0_0 ),
            .address1 ( buf_a1_0 ),
            .ce1      ( buf_ce1[ 0 ] ),
            .we1      ( buf_we1[ 0 ] ),
            .d1       ( buf_d1_0 )
        );
        td_fused_top_dataflow_in_loop_TOP_LOOP38022_accum1_out_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP38022_accum1_out_0_memcore_U_1 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_1 ),
            .ce0      ( buf_ce0[ 1 ] ),
            .we0      ( buf_we0[ 1 ] ),
            .d0       ( buf_d0_1 ),
            .q0       ( buf_q0_1 ),
            .address1 ( buf_a1_1 ),
            .ce1      ( buf_ce1[ 1 ] ),
            .we1      ( buf_we1[ 1 ] ),
            .d1       ( buf_d1_1 )
        );

//++++++++++++++++++++++++buffer signals+++++++++++++++++
        assign buf_ce0[ 0 ] = (tptr ==  0  && empty_n) ? t_ce0
                             : (iptr ==  0 ) ? i_ce0 : 1'b0;
        assign buf_a0_0  = (tptr ==  0  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 0 ] = (tptr ==  0  && empty_n)  ? t_we0
                             : (iptr ==  0 ) ? i_we0 : 1'b0;
        assign buf_d0_0  = (tptr ==  0  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 0 ] = (tptr ==  0  && empty_n) ? t_ce1
                             : (iptr ==  0 ) ? i_ce1 : 1'b0;
        assign buf_a1_0  = (tptr ==  0  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 0 ] = (tptr ==  0  && empty_n)  ? t_we1
                             : (iptr ==  0 ) ? i_we1 : 1'b0;
        assign buf_d1_0  = (tptr ==  0  && empty_n) ? t_d1       : i_d1;
        assign buf_ce0[ 1 ] = (tptr ==  1  && empty_n) ? t_ce0
                             : (iptr ==  1 ) ? i_ce0 : 1'b0;
        assign buf_a0_1  = (tptr ==  1  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 1 ] = (tptr ==  1  && empty_n)  ? t_we0
                             : (iptr ==  1 ) ? i_we0 : 1'b0;
        assign buf_d0_1  = (tptr ==  1  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 1 ] = (tptr ==  1  && empty_n) ? t_ce1
                             : (iptr ==  1 ) ? i_ce1 : 1'b0;
        assign buf_a1_1  = (tptr ==  1  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 1 ] = (tptr ==  1  && empty_n)  ? t_we1
                             : (iptr ==  1 ) ? i_we1 : 1'b0;
        assign buf_d1_1  = (tptr ==  1  && empty_n) ? t_d1       : i_d1;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//------------------------Body---------------------------
assign i_q0      = (prev_iptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign t_q0      = reg_valid0 ? reg_q0 : (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// prev_iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_iptr <= 1'b0;
    else begin
        prev_iptr <= iptr;
    end
end

// prev_tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_tptr <= 1'b0;
    else begin
        prev_tptr <= tptr;
    end
end

// reg_q0 and reg_valid0
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q0     <= 1'b0;
        reg_valid0 <= 1'b0;
    end else if (!t_ce0 && !reg_valid0) begin
        reg_q0     <= (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
        reg_valid0 <= 1'b1;
    end else if (t_ce0) begin
        reg_valid0 <= 1'b0;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP38022_ifmap_vec_memcore_ram (addr0, ce0, d0, we0, q0, addr1, ce1, d1, we1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 8;
parameter MEM_SIZE = 144;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
input clk;

reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];




always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1) 
            ram[addr1] <= d1; 
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP38022_ifmap_vec_memcore(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    q0,
    address1,
    ce1,
    we1,
    d1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd144;
parameter AddressWidth = 32'd8;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;



td_fused_top_dataflow_in_loop_TOP_LOOP38022_ifmap_vec_memcore_ram td_fused_top_dataflow_in_loop_TOP_LOOP38022_ifmap_vec_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_dataflow_in_loop_TOP_LOOP38022_ifmap_vec
#(parameter
    DataWidth    = 16,
    AddressRange = 32,
    AddressWidth = 8,
    BufferCount  = 2,
    MemLatency   = 1,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire                    i_we0,
    input  wire [AddressWidth-1:0] i_address0,
    input  wire [DataWidth-1:0]    i_d0,
    output wire [DataWidth-1:0]    i_q0,
    input  wire                    i_ce1,
    input  wire                    i_we1,
    input  wire [AddressWidth-1:0] i_address1,
    input  wire [DataWidth-1:0]    i_d1,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire                    t_we0,
    input  wire [AddressWidth-1:0] t_address0,
    input  wire [DataWidth-1:0]    t_d0,
    output wire [DataWidth-1:0]    t_q0,
    input  wire                    t_ce1,
    input  wire                    t_we1,
    input  wire [AddressWidth-1:0] t_address1,
    input  wire [DataWidth-1:0]    t_d1
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth-1:0]   prev_iptr    = 1'b0; // previous initiator index
reg  [IndexWidth-1:0]   prev_tptr    = 1'b0; // previous target index
reg  [DataWidth-1:0]    reg_q0      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid0    = 1'b0; // buffer has valid data
reg  [DataWidth-1:0]    reg_q1      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid1    = 1'b0; // buffer has valid data
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
// buffer signals
wire [BufferCount-1:0] buf_ce0;
wire [BufferCount-1:0] buf_we0;
wire [AddressWidth-1:0] buf_a0_0, buf_a0_1;
wire [DataWidth-1:0] buf_d0_0, buf_d0_1;
wire [DataWidth-1:0] buf_q0_0, buf_q0_1;
wire [BufferCount-1:0] buf_ce1;
wire [BufferCount-1:0] buf_we1;
wire [AddressWidth-1:0] buf_a1_0, buf_a1_1;
wire [DataWidth-1:0] buf_d1_0, buf_d1_1;
//------------------------Instantiation------------------
//genvar i;
        td_fused_top_dataflow_in_loop_TOP_LOOP38022_ifmap_vec_memcore td_fused_top_dataflow_in_loop_TOP_LOOP38022_ifmap_vec_memcore_U_0 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_0 ),
            .ce0      ( buf_ce0[ 0 ] ),
            .we0      ( buf_we0[ 0 ] ),
            .d0       ( buf_d0_0 ),
            .q0       ( buf_q0_0 ),
            .address1 ( buf_a1_0 ),
            .ce1      ( buf_ce1[ 0 ] ),
            .we1      ( buf_we1[ 0 ] ),
            .d1       ( buf_d1_0 )
        );
        td_fused_top_dataflow_in_loop_TOP_LOOP38022_ifmap_vec_memcore td_fused_top_dataflow_in_loop_TOP_LOOP38022_ifmap_vec_memcore_U_1 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_1 ),
            .ce0      ( buf_ce0[ 1 ] ),
            .we0      ( buf_we0[ 1 ] ),
            .d0       ( buf_d0_1 ),
            .q0       ( buf_q0_1 ),
            .address1 ( buf_a1_1 ),
            .ce1      ( buf_ce1[ 1 ] ),
            .we1      ( buf_we1[ 1 ] ),
            .d1       ( buf_d1_1 )
        );

//++++++++++++++++++++++++buffer signals+++++++++++++++++
        assign buf_ce0[ 0 ] = (tptr ==  0  && empty_n) ? t_ce0
                             : (iptr ==  0 ) ? i_ce0 : 1'b0;
        assign buf_a0_0  = (tptr ==  0  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 0 ] = (tptr ==  0  && empty_n)  ? t_we0
                             : (iptr ==  0 ) ? i_we0 : 1'b0;
        assign buf_d0_0  = (tptr ==  0  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 0 ] = (tptr ==  0  && empty_n) ? t_ce1
                             : (iptr ==  0 ) ? i_ce1 : 1'b0;
        assign buf_a1_0  = (tptr ==  0  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 0 ] = (tptr ==  0  && empty_n)  ? t_we1
                             : (iptr ==  0 ) ? i_we1 : 1'b0;
        assign buf_d1_0  = (tptr ==  0  && empty_n) ? t_d1       : i_d1;
        assign buf_ce0[ 1 ] = (tptr ==  1  && empty_n) ? t_ce0
                             : (iptr ==  1 ) ? i_ce0 : 1'b0;
        assign buf_a0_1  = (tptr ==  1  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 1 ] = (tptr ==  1  && empty_n)  ? t_we0
                             : (iptr ==  1 ) ? i_we0 : 1'b0;
        assign buf_d0_1  = (tptr ==  1  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 1 ] = (tptr ==  1  && empty_n) ? t_ce1
                             : (iptr ==  1 ) ? i_ce1 : 1'b0;
        assign buf_a1_1  = (tptr ==  1  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 1 ] = (tptr ==  1  && empty_n)  ? t_we1
                             : (iptr ==  1 ) ? i_we1 : 1'b0;
        assign buf_d1_1  = (tptr ==  1  && empty_n) ? t_d1       : i_d1;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//------------------------Body---------------------------
assign i_q0      = (prev_iptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign t_q0      = reg_valid0 ? reg_q0 : (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// prev_iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_iptr <= 1'b0;
    else begin
        prev_iptr <= iptr;
    end
end

// prev_tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_tptr <= 1'b0;
    else begin
        prev_tptr <= tptr;
    end
end

// reg_q0 and reg_valid0
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q0     <= 1'b0;
        reg_valid0 <= 1'b0;
    end else if (!t_ce0 && !reg_valid0) begin
        reg_q0     <= (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
        reg_valid0 <= 1'b1;
    end else if (t_ce0) begin
        reg_valid0 <= 1'b0;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP38022_products_0_memcore_ram (addr0, ce0, d0, we0, q0, addr1, ce1, q1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 8;
parameter MEM_SIZE = 144;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
output reg[DWIDTH-1:0] q1;
input clk;

reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];




always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        q1 <= ram[addr1];
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP38022_products_0_memcore(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    q0,
    address1,
    ce1,
    q1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd144;
parameter AddressWidth = 32'd8;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
output[DataWidth - 1:0] q1;



td_fused_top_dataflow_in_loop_TOP_LOOP38022_products_0_memcore_ram td_fused_top_dataflow_in_loop_TOP_LOOP38022_products_0_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .q1( q1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_dataflow_in_loop_TOP_LOOP38022_products_0
#(parameter
    DataWidth    = 16,
    AddressRange = 32,
    AddressWidth = 8,
    BufferCount  = 2,
    MemLatency   = 1,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire                    i_we0,
    input  wire [AddressWidth-1:0] i_address0,
    input  wire [DataWidth-1:0]    i_d0,
    output wire [DataWidth-1:0]    i_q0,
    input  wire                    i_ce1,
    input  wire [AddressWidth-1:0] i_address1,
    output wire [DataWidth-1:0]    i_q1,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire                    t_we0,
    input  wire [AddressWidth-1:0] t_address0,
    input  wire [DataWidth-1:0]    t_d0,
    output wire [DataWidth-1:0]    t_q0,
    input  wire                    t_ce1,
    input  wire [AddressWidth-1:0] t_address1,
    output wire [DataWidth-1:0]    t_q1
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth-1:0]   prev_iptr    = 1'b0; // previous initiator index
reg  [IndexWidth-1:0]   prev_tptr    = 1'b0; // previous target index
reg  [DataWidth-1:0]    reg_q0      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid0    = 1'b0; // buffer has valid data
reg  [DataWidth-1:0]    reg_q1      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid1    = 1'b0; // buffer has valid data
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
// buffer signals
wire [BufferCount-1:0] buf_ce0;
wire [BufferCount-1:0] buf_we0;
wire [AddressWidth-1:0] buf_a0_0, buf_a0_1;
wire [DataWidth-1:0] buf_d0_0, buf_d0_1;
wire [DataWidth-1:0] buf_q0_0, buf_q0_1;
wire [BufferCount-1:0] buf_ce1;
wire [AddressWidth-1:0] buf_a1_0, buf_a1_1;
wire [DataWidth-1:0] buf_q1_0, buf_q1_1;
//------------------------Instantiation------------------
//genvar i;
        td_fused_top_dataflow_in_loop_TOP_LOOP38022_products_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP38022_products_0_memcore_U_0 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_0 ),
            .ce0      ( buf_ce0[ 0 ] ),
            .we0      ( buf_we0[ 0 ] ),
            .d0       ( buf_d0_0 ),
            .q0       ( buf_q0_0 ),
            .address1 ( buf_a1_0 ),
            .ce1      ( buf_ce1[ 0 ] ),
            .q1       ( buf_q1_0 )
        );
        td_fused_top_dataflow_in_loop_TOP_LOOP38022_products_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP38022_products_0_memcore_U_1 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_1 ),
            .ce0      ( buf_ce0[ 1 ] ),
            .we0      ( buf_we0[ 1 ] ),
            .d0       ( buf_d0_1 ),
            .q0       ( buf_q0_1 ),
            .address1 ( buf_a1_1 ),
            .ce1      ( buf_ce1[ 1 ] ),
            .q1       ( buf_q1_1 )
        );

//++++++++++++++++++++++++buffer signals+++++++++++++++++
        assign buf_ce0[ 0 ] = (tptr ==  0  && empty_n) ? t_ce0
                             : (iptr ==  0 ) ? i_ce0 : 1'b0;
        assign buf_a0_0  = (tptr ==  0  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 0 ] = (tptr ==  0  && empty_n)  ? t_we0
                             : (iptr ==  0 ) ? i_we0 : 1'b0;
        assign buf_d0_0  = (tptr ==  0  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 0 ] = (tptr ==  0  && empty_n) ? t_ce1
                             : (iptr ==  0 ) ? i_ce1 : 1'b0;
        assign buf_a1_0  = (tptr ==  0  && empty_n) ?  t_address1 : i_address1;
        assign buf_ce0[ 1 ] = (tptr ==  1  && empty_n) ? t_ce0
                             : (iptr ==  1 ) ? i_ce0 : 1'b0;
        assign buf_a0_1  = (tptr ==  1  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 1 ] = (tptr ==  1  && empty_n)  ? t_we0
                             : (iptr ==  1 ) ? i_we0 : 1'b0;
        assign buf_d0_1  = (tptr ==  1  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 1 ] = (tptr ==  1  && empty_n) ? t_ce1
                             : (iptr ==  1 ) ? i_ce1 : 1'b0;
        assign buf_a1_1  = (tptr ==  1  && empty_n) ?  t_address1 : i_address1;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//------------------------Body---------------------------
assign i_q0      = (prev_iptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign t_q0      = reg_valid0 ? reg_q0 : (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign i_q1      = (prev_iptr == 1'b1 ? buf_q1_1 : buf_q1_0);
assign t_q1      = reg_valid1 ? reg_q1 : (prev_tptr == 1'b1 ? buf_q1_1 : buf_q1_0);

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// prev_iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_iptr <= 1'b0;
    else begin
        prev_iptr <= iptr;
    end
end

// prev_tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_tptr <= 1'b0;
    else begin
        prev_tptr <= tptr;
    end
end

// reg_q0 and reg_valid0
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q0     <= 1'b0;
        reg_valid0 <= 1'b0;
    end else if (!t_ce0 && !reg_valid0) begin
        reg_q0     <= (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
        reg_valid0 <= 1'b1;
    end else if (t_ce0) begin
        reg_valid0 <= 1'b0;
    end
end

// reg_q1 and reg_valid1
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q1     <= 1'b0;
        reg_valid1 <= 1'b0;
    end else if (!t_ce1 && !reg_valid1) begin
        reg_q1     <= (prev_tptr == 1'b1 ? buf_q1_1 : buf_q1_0);
        reg_valid1 <= 1'b1;
    end else if (t_ce1) begin
        reg_valid1 <= 1'b0;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_dataflow_in_loop_TOP_LOOP38022 (
        ap_clk,
        ap_rst,
        in_data_address0,
        in_data_ce0,
        in_data_d0,
        in_data_q0,
        in_data_we0,
        in_data_address1,
        in_data_ce1,
        in_data_d1,
        in_data_q1,
        in_data_we1,
        filter_data_address0,
        filter_data_ce0,
        filter_data_d0,
        filter_data_q0,
        filter_data_we0,
        filter_data_address1,
        filter_data_ce1,
        filter_data_d1,
        filter_data_q1,
        filter_data_we1,
        adjustments_address0,
        adjustments_ce0,
        adjustments_d0,
        adjustments_q0,
        adjustments_we0,
        adjustments_address1,
        adjustments_ce1,
        adjustments_d1,
        adjustments_q1,
        adjustments_we1,
        out_data_address0,
        out_data_ce0,
        out_data_d0,
        out_data_q0,
        out_data_we0,
        out_data_address1,
        out_data_ce1,
        out_data_d1,
        out_data_q1,
        out_data_we1,
        ap_start,
        in_data_empty_n,
        in_data_read,
        out_data_full_n,
        out_data_write,
        ap_done,
        ap_ready,
        ap_idle,
        ap_continue
);


input   ap_clk;
input   ap_rst;
output  [15:0] in_data_address0;
output   in_data_ce0;
output  [63:0] in_data_d0;
input  [63:0] in_data_q0;
output   in_data_we0;
output  [15:0] in_data_address1;
output   in_data_ce1;
output  [63:0] in_data_d1;
input  [63:0] in_data_q1;
output   in_data_we1;
output  [12:0] filter_data_address0;
output   filter_data_ce0;
output  [15:0] filter_data_d0;
input  [15:0] filter_data_q0;
output   filter_data_we0;
output  [12:0] filter_data_address1;
output   filter_data_ce1;
output  [15:0] filter_data_d1;
input  [15:0] filter_data_q1;
output   filter_data_we1;
output  [4:0] adjustments_address0;
output   adjustments_ce0;
output  [47:0] adjustments_d0;
input  [47:0] adjustments_q0;
output   adjustments_we0;
output  [4:0] adjustments_address1;
output   adjustments_ce1;
output  [47:0] adjustments_d1;
input  [47:0] adjustments_q1;
output   adjustments_we1;
output  [14:0] out_data_address0;
output   out_data_ce0;
output  [63:0] out_data_d0;
input  [63:0] out_data_q0;
output   out_data_we0;
output  [14:0] out_data_address1;
output   out_data_ce1;
output  [63:0] out_data_d1;
input  [63:0] out_data_q1;
output   out_data_we1;
input   ap_start;
input   in_data_empty_n;
output   in_data_read;
input   out_data_full_n;
output   out_data_write;
output   ap_done;
output   ap_ready;
output   ap_idle;
input   ap_continue;

wire   [15:0] ifmap_vec_i_q0;
wire   [15:0] ifmap_vec_t_q0;
wire   [15:0] weight_vecs_0_i_q0;
wire   [15:0] weight_vecs_0_t_q0;
wire   [15:0] products_0_i_q0;
wire   [15:0] products_0_i_q1;
wire   [15:0] products_0_t_q0;
wire   [15:0] products_0_t_q1;
wire   [15:0] accum1_out_0_i_q0;
wire   [15:0] accum1_out_0_t_q0;
wire    tdf2_get_next_ijk_U0_ap_start;
wire    tdf2_get_next_ijk_U0_ap_done;
wire    tdf2_get_next_ijk_U0_ap_continue;
wire    tdf2_get_next_ijk_U0_ap_idle;
wire    tdf2_get_next_ijk_U0_ap_ready;
wire    tdf2_get_next_ijk_U0_start_out;
wire    tdf2_get_next_ijk_U0_start_write;
wire   [4:0] tdf2_get_next_ijk_U0_input_indices_2_out_din;
wire    tdf2_get_next_ijk_U0_input_indices_2_out_write;
wire   [4:0] tdf2_get_next_ijk_U0_input_indices_2_out1_din;
wire    tdf2_get_next_ijk_U0_input_indices_2_out1_write;
wire   [5:0] tdf2_get_next_ijk_U0_output_indices_0_din;
wire    tdf2_get_next_ijk_U0_output_indices_0_write;
wire   [11:0] tdf2_get_next_ijk_U0_output_indices_1_din;
wire    tdf2_get_next_ijk_U0_output_indices_1_write;
wire    tdf2_get_next_ijk_U0_resetMaximum_din;
wire    tdf2_get_next_ijk_U0_resetMaximum_write;
wire    tdf2_get_next_ijk_U0_storeOutput_din;
wire    tdf2_get_next_ijk_U0_storeOutput_write;
wire   [15:0] tdf2_get_next_ijk_U0_ap_return_0;
wire   [15:0] tdf2_get_next_ijk_U0_ap_return_1;
wire    ap_channel_done_input_indices_1;
wire    input_indices_1_full_n;
reg    ap_sync_reg_channel_write_input_indices_1;
wire    ap_sync_channel_write_input_indices_1;
wire    ap_channel_done_input_indices_0;
wire    input_indices_0_full_n;
reg    ap_sync_reg_channel_write_input_indices_0;
wire    ap_sync_channel_write_input_indices_0;
wire    tdf2_readInputs25_U0_ap_start;
wire    tdf2_readInputs25_U0_ap_done;
wire    tdf2_readInputs25_U0_ap_continue;
wire    tdf2_readInputs25_U0_ap_idle;
wire    tdf2_readInputs25_U0_ap_ready;
wire   [15:0] tdf2_readInputs25_U0_in_data_address0;
wire    tdf2_readInputs25_U0_in_data_ce0;
wire   [7:0] tdf2_readInputs25_U0_ifmap_vec_address0;
wire    tdf2_readInputs25_U0_ifmap_vec_ce0;
wire    tdf2_readInputs25_U0_ifmap_vec_we0;
wire   [15:0] tdf2_readInputs25_U0_ifmap_vec_d0;
wire   [7:0] tdf2_readInputs25_U0_ifmap_vec_address1;
wire    tdf2_readInputs25_U0_ifmap_vec_ce1;
wire    tdf2_readInputs25_U0_ifmap_vec_we1;
wire   [15:0] tdf2_readInputs25_U0_ifmap_vec_d1;
wire    tdf2_readInputs25_U0_in_data_full_n;
wire    tdf2_readInputs25_U0_in_data_write;
wire    ap_channel_done_ifmap_vec;
wire    tdf2_readInputs25_U0_ifmap_vec_full_n;
wire    tdf2_readFilters24_U0_ap_start;
wire    tdf2_readFilters24_U0_ap_done;
wire    tdf2_readFilters24_U0_ap_continue;
wire    tdf2_readFilters24_U0_ap_idle;
wire    tdf2_readFilters24_U0_ap_ready;
wire   [12:0] tdf2_readFilters24_U0_filter_data_address0;
wire    tdf2_readFilters24_U0_filter_data_ce0;
wire    tdf2_readFilters24_U0_input_indices_23_read;
wire   [7:0] tdf2_readFilters24_U0_weight_vecs_0_address0;
wire    tdf2_readFilters24_U0_weight_vecs_0_ce0;
wire    tdf2_readFilters24_U0_weight_vecs_0_we0;
wire   [15:0] tdf2_readFilters24_U0_weight_vecs_0_d0;
wire    ap_channel_done_weight_vecs_0;
wire    tdf2_readFilters24_U0_weight_vecs_0_full_n;
wire    tdf2_dot_product_U0_ap_start;
wire    tdf2_dot_product_U0_ap_done;
wire    tdf2_dot_product_U0_ap_continue;
wire    tdf2_dot_product_U0_ap_idle;
wire    tdf2_dot_product_U0_ap_ready;
wire   [7:0] tdf2_dot_product_U0_ifmap_vec_address0;
wire    tdf2_dot_product_U0_ifmap_vec_ce0;
wire   [7:0] tdf2_dot_product_U0_weight_vecs_0_address0;
wire    tdf2_dot_product_U0_weight_vecs_0_ce0;
wire   [7:0] tdf2_dot_product_U0_products_0_address0;
wire    tdf2_dot_product_U0_products_0_ce0;
wire    tdf2_dot_product_U0_products_0_we0;
wire   [15:0] tdf2_dot_product_U0_products_0_d0;
wire    ap_channel_done_products_0;
wire    tdf2_dot_product_U0_products_0_full_n;
wire    tdf2_accum_1_U0_ap_start;
wire    tdf2_accum_1_U0_ap_done;
wire    tdf2_accum_1_U0_ap_continue;
wire    tdf2_accum_1_U0_ap_idle;
wire    tdf2_accum_1_U0_ap_ready;
wire   [7:0] tdf2_accum_1_U0_accum_in_0_address0;
wire    tdf2_accum_1_U0_accum_in_0_ce0;
wire   [7:0] tdf2_accum_1_U0_accum_in_0_address1;
wire    tdf2_accum_1_U0_accum_in_0_ce1;
wire   [2:0] tdf2_accum_1_U0_accum_out_address0;
wire    tdf2_accum_1_U0_accum_out_ce0;
wire    tdf2_accum_1_U0_accum_out_we0;
wire   [15:0] tdf2_accum_1_U0_accum_out_d0;
wire   [2:0] tdf2_accum_1_U0_accum_out_address1;
wire    tdf2_accum_1_U0_accum_out_ce1;
wire    tdf2_accum_1_U0_accum_out_we1;
wire   [15:0] tdf2_accum_1_U0_accum_out_d1;
wire    ap_channel_done_accum1_out_0;
wire    tdf2_accum_1_U0_accum_out_full_n;
wire    tdf2_accum_2_U0_ap_start;
wire    tdf2_accum_2_U0_ap_done;
wire    tdf2_accum_2_U0_ap_continue;
wire    tdf2_accum_2_U0_ap_idle;
wire    tdf2_accum_2_U0_ap_ready;
wire   [15:0] tdf2_accum_2_U0_accum_in_16;
wire    tdf2_accum_2_U0_accum_in_16_ap_vld;
wire   [2:0] tdf2_accum_2_U0_accum_in_address0;
wire    tdf2_accum_2_U0_accum_in_ce0;
wire    ap_channel_done_tmp_channel;
wire    tmp_channel_full_n;
wire    Block_entry_proc_proc392_U0_ap_start;
wire    Block_entry_proc_proc392_U0_ap_done;
wire    Block_entry_proc_proc392_U0_ap_continue;
wire    Block_entry_proc_proc392_U0_ap_idle;
wire    Block_entry_proc_proc392_U0_ap_ready;
wire   [15:0] Block_entry_proc_proc392_U0_ap_return;
wire    ap_channel_done_sums_0;
wire    sums_0_full_n;
wire    tdf2_adjust_U0_ap_start;
wire    tdf2_adjust_U0_ap_done;
wire    tdf2_adjust_U0_ap_continue;
wire    tdf2_adjust_U0_ap_idle;
wire    tdf2_adjust_U0_ap_ready;
wire   [4:0] tdf2_adjust_U0_adjustments_address0;
wire    tdf2_adjust_U0_adjustments_ce0;
wire    tdf2_adjust_U0_input_indices_23_read;
wire   [15:0] tdf2_adjust_U0_ap_return;
wire    ap_channel_done_outputs_0;
wire    outputs_0_full_n;
wire    tdf2_poolOutputs_U0_ap_start;
wire    tdf2_poolOutputs_U0_ap_done;
wire    tdf2_poolOutputs_U0_ap_continue;
wire    tdf2_poolOutputs_U0_ap_idle;
wire    tdf2_poolOutputs_U0_ap_ready;
wire    tdf2_poolOutputs_U0_output_indices_04_read;
wire    tdf2_poolOutputs_U0_output_indices_15_read;
wire    tdf2_poolOutputs_U0_resetMaximum6_read;
wire    tdf2_poolOutputs_U0_storeOutput7_read;
wire   [14:0] tdf2_poolOutputs_U0_out_data_address1;
wire    tdf2_poolOutputs_U0_out_data_ce1;
wire    tdf2_poolOutputs_U0_out_data_we1;
wire   [63:0] tdf2_poolOutputs_U0_out_data_d1;
wire    tdf2_poolOutputs_U0_out_data_full_n;
wire    tdf2_poolOutputs_U0_out_data_write;
wire    ap_sync_continue;
wire    ifmap_vec_i_full_n;
wire    ifmap_vec_t_empty_n;
wire    weight_vecs_0_i_full_n;
wire    weight_vecs_0_t_empty_n;
wire    products_0_i_full_n;
wire    products_0_t_empty_n;
wire   [15:0] products_0_t_d1;
wire    products_0_t_we1;
wire    accum1_out_0_i_full_n;
wire    accum1_out_0_t_empty_n;
wire    input_indices_23_c_full_n;
wire   [4:0] input_indices_23_c_dout;
wire    input_indices_23_c_empty_n;
wire    input_indices_23_c1_full_n;
wire   [4:0] input_indices_23_c1_dout;
wire    input_indices_23_c1_empty_n;
wire    output_indices_04_c_full_n;
wire   [5:0] output_indices_04_c_dout;
wire    output_indices_04_c_empty_n;
wire    output_indices_15_c_full_n;
wire   [11:0] output_indices_15_c_dout;
wire    output_indices_15_c_empty_n;
wire   [0:0] resetMaximum6_c_din;
wire    resetMaximum6_c_full_n;
wire   [0:0] resetMaximum6_c_dout;
wire    resetMaximum6_c_empty_n;
wire   [0:0] storeOutput7_c_din;
wire    storeOutput7_c_full_n;
wire   [0:0] storeOutput7_c_dout;
wire    storeOutput7_c_empty_n;
wire   [15:0] input_indices_0_dout;
wire    input_indices_0_empty_n;
wire   [15:0] input_indices_1_dout;
wire    input_indices_1_empty_n;
wire   [15:0] tmp_channel_dout;
wire    tmp_channel_empty_n;
wire   [15:0] sums_0_dout;
wire    sums_0_empty_n;
wire   [15:0] outputs_0_dout;
wire    outputs_0_empty_n;
wire    ap_sync_done;
wire    ap_sync_ready;
reg    ap_sync_reg_tdf2_get_next_ijk_U0_ap_ready;
wire    ap_sync_tdf2_get_next_ijk_U0_ap_ready;
reg    ap_sync_reg_tdf2_readInputs25_U0_ap_ready;
wire    ap_sync_tdf2_readInputs25_U0_ap_ready;
wire   [0:0] start_for_tdf2_readFilters24_U0_din;
wire    start_for_tdf2_readFilters24_U0_full_n;
wire   [0:0] start_for_tdf2_readFilters24_U0_dout;
wire    start_for_tdf2_readFilters24_U0_empty_n;
wire    tdf2_readInputs25_U0_start_full_n;
wire    tdf2_readInputs25_U0_start_write;
wire    tdf2_readFilters24_U0_start_full_n;
wire    tdf2_readFilters24_U0_start_write;
wire    tdf2_dot_product_U0_start_full_n;
wire    tdf2_dot_product_U0_start_write;
wire    tdf2_accum_1_U0_start_full_n;
wire    tdf2_accum_1_U0_start_write;
wire    tdf2_accum_2_U0_start_full_n;
wire    tdf2_accum_2_U0_start_write;
wire    Block_entry_proc_proc392_U0_start_full_n;
wire    Block_entry_proc_proc392_U0_start_write;
wire    tdf2_adjust_U0_start_full_n;
wire    tdf2_adjust_U0_start_write;
wire    tdf2_poolOutputs_U0_start_full_n;
wire    tdf2_poolOutputs_U0_start_write;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_sync_reg_channel_write_input_indices_1 = 1'b0;
#0 ap_sync_reg_channel_write_input_indices_0 = 1'b0;
#0 ap_sync_reg_tdf2_get_next_ijk_U0_ap_ready = 1'b0;
#0 ap_sync_reg_tdf2_readInputs25_U0_ap_ready = 1'b0;
end

td_fused_top_dataflow_in_loop_TOP_LOOP38022_ifmap_vec #(
    .DataWidth( 16 ),
    .AddressRange( 144 ),
    .AddressWidth( 8 ))
ifmap_vec_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf2_readInputs25_U0_ap_done),
    .i_full_n(ifmap_vec_i_full_n),
    .i_ce0(tdf2_readInputs25_U0_ifmap_vec_ce0),
    .i_we0(tdf2_readInputs25_U0_ifmap_vec_we0),
    .i_address0(tdf2_readInputs25_U0_ifmap_vec_address0),
    .i_d0(tdf2_readInputs25_U0_ifmap_vec_d0),
    .i_q0(ifmap_vec_i_q0),
    .i_ce1(tdf2_readInputs25_U0_ifmap_vec_ce1),
    .i_we1(tdf2_readInputs25_U0_ifmap_vec_we1),
    .i_address1(tdf2_readInputs25_U0_ifmap_vec_address1),
    .i_d1(tdf2_readInputs25_U0_ifmap_vec_d1),
    .t_ce(1'b1),
    .t_read(tdf2_dot_product_U0_ap_ready),
    .t_empty_n(ifmap_vec_t_empty_n),
    .t_ce0(tdf2_dot_product_U0_ifmap_vec_ce0),
    .t_we0(1'b0),
    .t_address0(tdf2_dot_product_U0_ifmap_vec_address0),
    .t_d0(16'd0),
    .t_q0(ifmap_vec_t_q0),
    .t_ce1(1'b0),
    .t_we1(1'b0),
    .t_address1(8'd0),
    .t_d1(16'd0)
);

td_fused_top_dataflow_in_loop_TOP_LOOP38022_weight_vecs_0 #(
    .DataWidth( 16 ),
    .AddressRange( 144 ),
    .AddressWidth( 8 ))
weight_vecs_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf2_readFilters24_U0_ap_done),
    .i_full_n(weight_vecs_0_i_full_n),
    .i_ce0(tdf2_readFilters24_U0_weight_vecs_0_ce0),
    .i_we0(tdf2_readFilters24_U0_weight_vecs_0_we0),
    .i_address0(tdf2_readFilters24_U0_weight_vecs_0_address0),
    .i_d0(tdf2_readFilters24_U0_weight_vecs_0_d0),
    .i_q0(weight_vecs_0_i_q0),
    .t_ce(1'b1),
    .t_read(tdf2_dot_product_U0_ap_ready),
    .t_empty_n(weight_vecs_0_t_empty_n),
    .t_ce0(tdf2_dot_product_U0_weight_vecs_0_ce0),
    .t_we0(1'b0),
    .t_address0(tdf2_dot_product_U0_weight_vecs_0_address0),
    .t_d0(16'd0),
    .t_q0(weight_vecs_0_t_q0)
);

td_fused_top_dataflow_in_loop_TOP_LOOP38022_products_0 #(
    .DataWidth( 16 ),
    .AddressRange( 144 ),
    .AddressWidth( 8 ))
products_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf2_dot_product_U0_ap_done),
    .i_full_n(products_0_i_full_n),
    .i_ce0(tdf2_dot_product_U0_products_0_ce0),
    .i_we0(tdf2_dot_product_U0_products_0_we0),
    .i_address0(tdf2_dot_product_U0_products_0_address0),
    .i_d0(tdf2_dot_product_U0_products_0_d0),
    .i_q0(products_0_i_q0),
    .i_ce1(1'b0),
    .i_address1(8'd0),
    .i_q1(products_0_i_q1),
    .t_ce(1'b1),
    .t_read(tdf2_accum_1_U0_ap_ready),
    .t_empty_n(products_0_t_empty_n),
    .t_ce0(tdf2_accum_1_U0_accum_in_0_ce0),
    .t_we0(1'b0),
    .t_address0(tdf2_accum_1_U0_accum_in_0_address0),
    .t_d0(16'd0),
    .t_q0(products_0_t_q0),
    .t_ce1(tdf2_accum_1_U0_accum_in_0_ce1),
    .t_address1(tdf2_accum_1_U0_accum_in_0_address1),
    .t_q1(products_0_t_q1)
);

td_fused_top_dataflow_in_loop_TOP_LOOP38022_accum1_out_0 #(
    .DataWidth( 16 ),
    .AddressRange( 8 ),
    .AddressWidth( 3 ))
accum1_out_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf2_accum_1_U0_ap_done),
    .i_full_n(accum1_out_0_i_full_n),
    .i_ce0(tdf2_accum_1_U0_accum_out_ce0),
    .i_we0(tdf2_accum_1_U0_accum_out_we0),
    .i_address0(tdf2_accum_1_U0_accum_out_address0),
    .i_d0(tdf2_accum_1_U0_accum_out_d0),
    .i_q0(accum1_out_0_i_q0),
    .i_ce1(tdf2_accum_1_U0_accum_out_ce1),
    .i_we1(tdf2_accum_1_U0_accum_out_we1),
    .i_address1(tdf2_accum_1_U0_accum_out_address1),
    .i_d1(tdf2_accum_1_U0_accum_out_d1),
    .t_ce(1'b1),
    .t_read(tdf2_accum_2_U0_ap_ready),
    .t_empty_n(accum1_out_0_t_empty_n),
    .t_ce0(tdf2_accum_2_U0_accum_in_ce0),
    .t_we0(1'b0),
    .t_address0(tdf2_accum_2_U0_accum_in_address0),
    .t_d0(16'd0),
    .t_q0(accum1_out_0_t_q0),
    .t_ce1(1'b0),
    .t_we1(1'b0),
    .t_address1(3'd0),
    .t_d1(16'd0)
);

td_fused_top_tdf2_get_next_ijk tdf2_get_next_ijk_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf2_get_next_ijk_U0_ap_start),
    .start_full_n(start_for_tdf2_readFilters24_U0_full_n),
    .ap_done(tdf2_get_next_ijk_U0_ap_done),
    .ap_continue(tdf2_get_next_ijk_U0_ap_continue),
    .ap_idle(tdf2_get_next_ijk_U0_ap_idle),
    .ap_ready(tdf2_get_next_ijk_U0_ap_ready),
    .start_out(tdf2_get_next_ijk_U0_start_out),
    .start_write(tdf2_get_next_ijk_U0_start_write),
    .input_indices_2_out_din(tdf2_get_next_ijk_U0_input_indices_2_out_din),
    .input_indices_2_out_full_n(input_indices_23_c_full_n),
    .input_indices_2_out_write(tdf2_get_next_ijk_U0_input_indices_2_out_write),
    .input_indices_2_out1_din(tdf2_get_next_ijk_U0_input_indices_2_out1_din),
    .input_indices_2_out1_full_n(input_indices_23_c1_full_n),
    .input_indices_2_out1_write(tdf2_get_next_ijk_U0_input_indices_2_out1_write),
    .output_indices_0_din(tdf2_get_next_ijk_U0_output_indices_0_din),
    .output_indices_0_full_n(output_indices_04_c_full_n),
    .output_indices_0_write(tdf2_get_next_ijk_U0_output_indices_0_write),
    .output_indices_1_din(tdf2_get_next_ijk_U0_output_indices_1_din),
    .output_indices_1_full_n(output_indices_15_c_full_n),
    .output_indices_1_write(tdf2_get_next_ijk_U0_output_indices_1_write),
    .resetMaximum_din(tdf2_get_next_ijk_U0_resetMaximum_din),
    .resetMaximum_full_n(resetMaximum6_c_full_n),
    .resetMaximum_write(tdf2_get_next_ijk_U0_resetMaximum_write),
    .storeOutput_din(tdf2_get_next_ijk_U0_storeOutput_din),
    .storeOutput_full_n(storeOutput7_c_full_n),
    .storeOutput_write(tdf2_get_next_ijk_U0_storeOutput_write),
    .ap_return_0(tdf2_get_next_ijk_U0_ap_return_0),
    .ap_return_1(tdf2_get_next_ijk_U0_ap_return_1)
);

td_fused_top_tdf2_readInputs25 tdf2_readInputs25_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf2_readInputs25_U0_ap_start),
    .ap_done(tdf2_readInputs25_U0_ap_done),
    .ap_continue(tdf2_readInputs25_U0_ap_continue),
    .ap_idle(tdf2_readInputs25_U0_ap_idle),
    .ap_ready(tdf2_readInputs25_U0_ap_ready),
    .in_data_address0(tdf2_readInputs25_U0_in_data_address0),
    .in_data_ce0(tdf2_readInputs25_U0_in_data_ce0),
    .in_data_q0(in_data_q0),
    .i_17(input_indices_0_dout),
    .j_17(input_indices_1_dout),
    .ifmap_vec_address0(tdf2_readInputs25_U0_ifmap_vec_address0),
    .ifmap_vec_ce0(tdf2_readInputs25_U0_ifmap_vec_ce0),
    .ifmap_vec_we0(tdf2_readInputs25_U0_ifmap_vec_we0),
    .ifmap_vec_d0(tdf2_readInputs25_U0_ifmap_vec_d0),
    .ifmap_vec_address1(tdf2_readInputs25_U0_ifmap_vec_address1),
    .ifmap_vec_ce1(tdf2_readInputs25_U0_ifmap_vec_ce1),
    .ifmap_vec_we1(tdf2_readInputs25_U0_ifmap_vec_we1),
    .ifmap_vec_d1(tdf2_readInputs25_U0_ifmap_vec_d1)
);

td_fused_top_tdf2_readFilters24 tdf2_readFilters24_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf2_readFilters24_U0_ap_start),
    .ap_done(tdf2_readFilters24_U0_ap_done),
    .ap_continue(tdf2_readFilters24_U0_ap_continue),
    .ap_idle(tdf2_readFilters24_U0_ap_idle),
    .ap_ready(tdf2_readFilters24_U0_ap_ready),
    .filter_data_address0(tdf2_readFilters24_U0_filter_data_address0),
    .filter_data_ce0(tdf2_readFilters24_U0_filter_data_ce0),
    .filter_data_q0(filter_data_q0),
    .input_indices_23_dout(input_indices_23_c_dout),
    .input_indices_23_empty_n(input_indices_23_c_empty_n),
    .input_indices_23_read(tdf2_readFilters24_U0_input_indices_23_read),
    .weight_vecs_0_address0(tdf2_readFilters24_U0_weight_vecs_0_address0),
    .weight_vecs_0_ce0(tdf2_readFilters24_U0_weight_vecs_0_ce0),
    .weight_vecs_0_we0(tdf2_readFilters24_U0_weight_vecs_0_we0),
    .weight_vecs_0_d0(tdf2_readFilters24_U0_weight_vecs_0_d0)
);

td_fused_top_tdf2_dot_product tdf2_dot_product_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf2_dot_product_U0_ap_start),
    .ap_done(tdf2_dot_product_U0_ap_done),
    .ap_continue(tdf2_dot_product_U0_ap_continue),
    .ap_idle(tdf2_dot_product_U0_ap_idle),
    .ap_ready(tdf2_dot_product_U0_ap_ready),
    .ifmap_vec_address0(tdf2_dot_product_U0_ifmap_vec_address0),
    .ifmap_vec_ce0(tdf2_dot_product_U0_ifmap_vec_ce0),
    .ifmap_vec_q0(ifmap_vec_t_q0),
    .weight_vecs_0_address0(tdf2_dot_product_U0_weight_vecs_0_address0),
    .weight_vecs_0_ce0(tdf2_dot_product_U0_weight_vecs_0_ce0),
    .weight_vecs_0_q0(weight_vecs_0_t_q0),
    .products_0_address0(tdf2_dot_product_U0_products_0_address0),
    .products_0_ce0(tdf2_dot_product_U0_products_0_ce0),
    .products_0_we0(tdf2_dot_product_U0_products_0_we0),
    .products_0_d0(tdf2_dot_product_U0_products_0_d0)
);

td_fused_top_tdf2_accum_1 tdf2_accum_1_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf2_accum_1_U0_ap_start),
    .ap_done(tdf2_accum_1_U0_ap_done),
    .ap_continue(tdf2_accum_1_U0_ap_continue),
    .ap_idle(tdf2_accum_1_U0_ap_idle),
    .ap_ready(tdf2_accum_1_U0_ap_ready),
    .accum_in_0_address0(tdf2_accum_1_U0_accum_in_0_address0),
    .accum_in_0_ce0(tdf2_accum_1_U0_accum_in_0_ce0),
    .accum_in_0_q0(products_0_t_q0),
    .accum_in_0_address1(tdf2_accum_1_U0_accum_in_0_address1),
    .accum_in_0_ce1(tdf2_accum_1_U0_accum_in_0_ce1),
    .accum_in_0_q1(products_0_t_q1),
    .accum_out_address0(tdf2_accum_1_U0_accum_out_address0),
    .accum_out_ce0(tdf2_accum_1_U0_accum_out_ce0),
    .accum_out_we0(tdf2_accum_1_U0_accum_out_we0),
    .accum_out_d0(tdf2_accum_1_U0_accum_out_d0),
    .accum_out_address1(tdf2_accum_1_U0_accum_out_address1),
    .accum_out_ce1(tdf2_accum_1_U0_accum_out_ce1),
    .accum_out_we1(tdf2_accum_1_U0_accum_out_we1),
    .accum_out_d1(tdf2_accum_1_U0_accum_out_d1)
);

td_fused_top_tdf2_accum_2 tdf2_accum_2_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf2_accum_2_U0_ap_start),
    .ap_done(tdf2_accum_2_U0_ap_done),
    .ap_continue(tdf2_accum_2_U0_ap_continue),
    .ap_idle(tdf2_accum_2_U0_ap_idle),
    .ap_ready(tdf2_accum_2_U0_ap_ready),
    .accum_in_16(tdf2_accum_2_U0_accum_in_16),
    .accum_in_16_ap_vld(tdf2_accum_2_U0_accum_in_16_ap_vld),
    .accum_in_address0(tdf2_accum_2_U0_accum_in_address0),
    .accum_in_ce0(tdf2_accum_2_U0_accum_in_ce0),
    .accum_in_q0(accum1_out_0_t_q0)
);

td_fused_top_Block_entry_proc_proc392 Block_entry_proc_proc392_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(Block_entry_proc_proc392_U0_ap_start),
    .ap_done(Block_entry_proc_proc392_U0_ap_done),
    .ap_continue(Block_entry_proc_proc392_U0_ap_continue),
    .ap_idle(Block_entry_proc_proc392_U0_ap_idle),
    .ap_ready(Block_entry_proc_proc392_U0_ap_ready),
    .tmp(tmp_channel_dout),
    .ap_return(Block_entry_proc_proc392_U0_ap_return)
);

td_fused_top_tdf2_adjust tdf2_adjust_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf2_adjust_U0_ap_start),
    .ap_done(tdf2_adjust_U0_ap_done),
    .ap_continue(tdf2_adjust_U0_ap_continue),
    .ap_idle(tdf2_adjust_U0_ap_idle),
    .ap_ready(tdf2_adjust_U0_ap_ready),
    .sums_read(sums_0_dout),
    .adjustments_address0(tdf2_adjust_U0_adjustments_address0),
    .adjustments_ce0(tdf2_adjust_U0_adjustments_ce0),
    .adjustments_q0(adjustments_q0),
    .input_indices_23_dout(input_indices_23_c1_dout),
    .input_indices_23_empty_n(input_indices_23_c1_empty_n),
    .input_indices_23_read(tdf2_adjust_U0_input_indices_23_read),
    .ap_return(tdf2_adjust_U0_ap_return)
);

td_fused_top_tdf2_poolOutputs tdf2_poolOutputs_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf2_poolOutputs_U0_ap_start),
    .ap_done(tdf2_poolOutputs_U0_ap_done),
    .ap_continue(tdf2_poolOutputs_U0_ap_continue),
    .ap_idle(tdf2_poolOutputs_U0_ap_idle),
    .ap_ready(tdf2_poolOutputs_U0_ap_ready),
    .output_indices_04_dout(output_indices_04_c_dout),
    .output_indices_04_empty_n(output_indices_04_c_empty_n),
    .output_indices_04_read(tdf2_poolOutputs_U0_output_indices_04_read),
    .output_indices_15_dout(output_indices_15_c_dout),
    .output_indices_15_empty_n(output_indices_15_c_empty_n),
    .output_indices_15_read(tdf2_poolOutputs_U0_output_indices_15_read),
    .resetMaximum6_dout(resetMaximum6_c_dout),
    .resetMaximum6_empty_n(resetMaximum6_c_empty_n),
    .resetMaximum6_read(tdf2_poolOutputs_U0_resetMaximum6_read),
    .storeOutput7_dout(storeOutput7_c_dout),
    .storeOutput7_empty_n(storeOutput7_c_empty_n),
    .storeOutput7_read(tdf2_poolOutputs_U0_storeOutput7_read),
    .p_read(outputs_0_dout),
    .out_data_address1(tdf2_poolOutputs_U0_out_data_address1),
    .out_data_ce1(tdf2_poolOutputs_U0_out_data_ce1),
    .out_data_we1(tdf2_poolOutputs_U0_out_data_we1),
    .out_data_d1(tdf2_poolOutputs_U0_out_data_d1)
);

td_fused_top_fifo_w5_d2_S input_indices_23_c_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(input_indices_23_c_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf2_readFilters24_U0_input_indices_23_read),
    .if_dout(input_indices_23_c_dout),
    .if_full_n(input_indices_23_c_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf2_get_next_ijk_U0_input_indices_2_out_write),
    .if_din(tdf2_get_next_ijk_U0_input_indices_2_out_din)
);

td_fused_top_fifo_w5_d7_S input_indices_23_c1_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(input_indices_23_c1_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf2_adjust_U0_input_indices_23_read),
    .if_dout(input_indices_23_c1_dout),
    .if_full_n(input_indices_23_c1_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf2_get_next_ijk_U0_input_indices_2_out1_write),
    .if_din(tdf2_get_next_ijk_U0_input_indices_2_out1_din)
);

td_fused_top_fifo_w6_d8_S output_indices_04_c_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(output_indices_04_c_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf2_poolOutputs_U0_output_indices_04_read),
    .if_dout(output_indices_04_c_dout),
    .if_full_n(output_indices_04_c_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf2_get_next_ijk_U0_output_indices_0_write),
    .if_din(tdf2_get_next_ijk_U0_output_indices_0_din)
);

td_fused_top_fifo_w12_d8_S output_indices_15_c_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(output_indices_15_c_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf2_poolOutputs_U0_output_indices_15_read),
    .if_dout(output_indices_15_c_dout),
    .if_full_n(output_indices_15_c_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf2_get_next_ijk_U0_output_indices_1_write),
    .if_din(tdf2_get_next_ijk_U0_output_indices_1_din)
);

td_fused_top_fifo_w1_d8_S resetMaximum6_c_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(resetMaximum6_c_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf2_poolOutputs_U0_resetMaximum6_read),
    .if_dout(resetMaximum6_c_dout),
    .if_full_n(resetMaximum6_c_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf2_get_next_ijk_U0_resetMaximum_write),
    .if_din(resetMaximum6_c_din)
);

td_fused_top_fifo_w1_d8_S storeOutput7_c_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(storeOutput7_c_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf2_poolOutputs_U0_storeOutput7_read),
    .if_dout(storeOutput7_c_dout),
    .if_full_n(storeOutput7_c_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf2_get_next_ijk_U0_storeOutput_write),
    .if_din(storeOutput7_c_din)
);

td_fused_top_fifo_w16_d2_S_x input_indices_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(input_indices_0_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf2_readInputs25_U0_ap_ready),
    .if_dout(input_indices_0_dout),
    .if_full_n(input_indices_0_full_n),
    .if_write_ce(1'b1),
    .if_write(ap_channel_done_input_indices_0),
    .if_din(tdf2_get_next_ijk_U0_ap_return_0)
);

td_fused_top_fifo_w16_d2_S_x input_indices_1_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(input_indices_1_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf2_readInputs25_U0_ap_ready),
    .if_dout(input_indices_1_dout),
    .if_full_n(input_indices_1_full_n),
    .if_write_ce(1'b1),
    .if_write(ap_channel_done_input_indices_1),
    .if_din(tdf2_get_next_ijk_U0_ap_return_1)
);

td_fused_top_fifo_w16_d2_S_x tmp_channel_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(tmp_channel_empty_n),
    .if_read_ce(1'b1),
    .if_read(Block_entry_proc_proc392_U0_ap_ready),
    .if_dout(tmp_channel_dout),
    .if_full_n(tmp_channel_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf2_accum_2_U0_ap_done),
    .if_din(tdf2_accum_2_U0_accum_in_16)
);

td_fused_top_fifo_w16_d2_S_x sums_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(sums_0_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf2_adjust_U0_ap_ready),
    .if_dout(sums_0_dout),
    .if_full_n(sums_0_full_n),
    .if_write_ce(1'b1),
    .if_write(Block_entry_proc_proc392_U0_ap_done),
    .if_din(Block_entry_proc_proc392_U0_ap_return)
);

td_fused_top_fifo_w16_d2_S_x outputs_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(outputs_0_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf2_poolOutputs_U0_ap_ready),
    .if_dout(outputs_0_dout),
    .if_full_n(outputs_0_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf2_adjust_U0_ap_done),
    .if_din(tdf2_adjust_U0_ap_return)
);

td_fused_top_start_for_tdf2_readFilters24_U0 start_for_tdf2_readFilters24_U0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(start_for_tdf2_readFilters24_U0_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf2_readFilters24_U0_ap_ready),
    .if_dout(start_for_tdf2_readFilters24_U0_dout),
    .if_full_n(start_for_tdf2_readFilters24_U0_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf2_get_next_ijk_U0_start_write),
    .if_din(start_for_tdf2_readFilters24_U0_din)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_sync_reg_channel_write_input_indices_0 <= 1'b0;
    end else begin
        if (((tdf2_get_next_ijk_U0_ap_done & tdf2_get_next_ijk_U0_ap_continue) == 1'b1)) begin
            ap_sync_reg_channel_write_input_indices_0 <= 1'b0;
        end else begin
            ap_sync_reg_channel_write_input_indices_0 <= ap_sync_channel_write_input_indices_0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_sync_reg_channel_write_input_indices_1 <= 1'b0;
    end else begin
        if (((tdf2_get_next_ijk_U0_ap_done & tdf2_get_next_ijk_U0_ap_continue) == 1'b1)) begin
            ap_sync_reg_channel_write_input_indices_1 <= 1'b0;
        end else begin
            ap_sync_reg_channel_write_input_indices_1 <= ap_sync_channel_write_input_indices_1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_sync_reg_tdf2_get_next_ijk_U0_ap_ready <= 1'b0;
    end else begin
        if (((ap_sync_ready & ap_start) == 1'b1)) begin
            ap_sync_reg_tdf2_get_next_ijk_U0_ap_ready <= 1'b0;
        end else begin
            ap_sync_reg_tdf2_get_next_ijk_U0_ap_ready <= ap_sync_tdf2_get_next_ijk_U0_ap_ready;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_sync_reg_tdf2_readInputs25_U0_ap_ready <= 1'b0;
    end else begin
        if (((ap_sync_ready & ap_start) == 1'b1)) begin
            ap_sync_reg_tdf2_readInputs25_U0_ap_ready <= 1'b0;
        end else begin
            ap_sync_reg_tdf2_readInputs25_U0_ap_ready <= ap_sync_tdf2_readInputs25_U0_ap_ready;
        end
    end
end

assign Block_entry_proc_proc392_U0_ap_continue = sums_0_full_n;

assign Block_entry_proc_proc392_U0_ap_start = tmp_channel_empty_n;

assign Block_entry_proc_proc392_U0_start_full_n = 1'b1;

assign Block_entry_proc_proc392_U0_start_write = 1'b0;

assign adjustments_address0 = tdf2_adjust_U0_adjustments_address0;

assign adjustments_address1 = 5'd0;

assign adjustments_ce0 = tdf2_adjust_U0_adjustments_ce0;

assign adjustments_ce1 = 1'b0;

assign adjustments_d0 = 48'd0;

assign adjustments_d1 = 48'd0;

assign adjustments_we0 = 1'b0;

assign adjustments_we1 = 1'b0;

assign ap_channel_done_accum1_out_0 = tdf2_accum_1_U0_ap_done;

assign ap_channel_done_ifmap_vec = tdf2_readInputs25_U0_ap_done;

assign ap_channel_done_input_indices_0 = (tdf2_get_next_ijk_U0_ap_done & (ap_sync_reg_channel_write_input_indices_0 ^ 1'b1));

assign ap_channel_done_input_indices_1 = (tdf2_get_next_ijk_U0_ap_done & (ap_sync_reg_channel_write_input_indices_1 ^ 1'b1));

assign ap_channel_done_outputs_0 = tdf2_adjust_U0_ap_done;

assign ap_channel_done_products_0 = tdf2_dot_product_U0_ap_done;

assign ap_channel_done_sums_0 = Block_entry_proc_proc392_U0_ap_done;

assign ap_channel_done_tmp_channel = tdf2_accum_2_U0_ap_done;

assign ap_channel_done_weight_vecs_0 = tdf2_readFilters24_U0_ap_done;

assign ap_done = tdf2_poolOutputs_U0_ap_done;

assign ap_idle = (tdf2_readInputs25_U0_ap_idle & tdf2_readFilters24_U0_ap_idle & tdf2_poolOutputs_U0_ap_idle & tdf2_get_next_ijk_U0_ap_idle & tdf2_dot_product_U0_ap_idle & tdf2_adjust_U0_ap_idle & tdf2_accum_2_U0_ap_idle & tdf2_accum_1_U0_ap_idle & (outputs_0_empty_n ^ 1'b1) & (sums_0_empty_n ^ 1'b1) & (tmp_channel_empty_n ^ 1'b1) & (input_indices_1_empty_n ^ 1'b1) & (input_indices_0_empty_n ^ 1'b1) & (products_0_t_empty_n ^ 1'b1) & (weight_vecs_0_t_empty_n ^ 1'b1) & (ifmap_vec_t_empty_n ^ 1'b1) & (1'b1 ^ accum1_out_0_t_empty_n) & Block_entry_proc_proc392_U0_ap_idle);

assign ap_ready = ap_sync_ready;

assign ap_sync_channel_write_input_indices_0 = ((input_indices_0_full_n & ap_channel_done_input_indices_0) | ap_sync_reg_channel_write_input_indices_0);

assign ap_sync_channel_write_input_indices_1 = ((input_indices_1_full_n & ap_channel_done_input_indices_1) | ap_sync_reg_channel_write_input_indices_1);

assign ap_sync_continue = ap_continue;

assign ap_sync_done = tdf2_poolOutputs_U0_ap_done;

assign ap_sync_ready = (ap_sync_tdf2_readInputs25_U0_ap_ready & ap_sync_tdf2_get_next_ijk_U0_ap_ready);

assign ap_sync_tdf2_get_next_ijk_U0_ap_ready = (tdf2_get_next_ijk_U0_ap_ready | ap_sync_reg_tdf2_get_next_ijk_U0_ap_ready);

assign ap_sync_tdf2_readInputs25_U0_ap_ready = (tdf2_readInputs25_U0_ap_ready | ap_sync_reg_tdf2_readInputs25_U0_ap_ready);

assign filter_data_address0 = tdf2_readFilters24_U0_filter_data_address0;

assign filter_data_address1 = 13'd0;

assign filter_data_ce0 = tdf2_readFilters24_U0_filter_data_ce0;

assign filter_data_ce1 = 1'b0;

assign filter_data_d0 = 16'd0;

assign filter_data_d1 = 16'd0;

assign filter_data_we0 = 1'b0;

assign filter_data_we1 = 1'b0;

assign in_data_address0 = tdf2_readInputs25_U0_in_data_address0;

assign in_data_address1 = 16'd0;

assign in_data_ce0 = tdf2_readInputs25_U0_in_data_ce0;

assign in_data_ce1 = 1'b0;

assign in_data_d0 = 64'd0;

assign in_data_d1 = 64'd0;

assign in_data_read = tdf2_readInputs25_U0_in_data_write;

assign in_data_we0 = 1'b0;

assign in_data_we1 = 1'b0;

assign out_data_address0 = 15'd0;

assign out_data_address1 = tdf2_poolOutputs_U0_out_data_address1;

assign out_data_ce0 = 1'b0;

assign out_data_ce1 = tdf2_poolOutputs_U0_out_data_ce1;

assign out_data_d0 = 64'd0;

assign out_data_d1 = tdf2_poolOutputs_U0_out_data_d1;

assign out_data_we0 = 1'b0;

assign out_data_we1 = tdf2_poolOutputs_U0_out_data_we1;

assign out_data_write = tdf2_poolOutputs_U0_out_data_write;

assign products_0_t_d1 = 16'd0;

assign products_0_t_we1 = 1'b0;

assign resetMaximum6_c_din = tdf2_get_next_ijk_U0_resetMaximum_din;

assign start_for_tdf2_readFilters24_U0_din = 1'b1;

assign storeOutput7_c_din = tdf2_get_next_ijk_U0_storeOutput_din;

assign tdf2_accum_1_U0_accum_out_full_n = accum1_out_0_i_full_n;

assign tdf2_accum_1_U0_ap_continue = accum1_out_0_i_full_n;

assign tdf2_accum_1_U0_ap_start = products_0_t_empty_n;

assign tdf2_accum_1_U0_start_full_n = 1'b1;

assign tdf2_accum_1_U0_start_write = 1'b0;

assign tdf2_accum_2_U0_ap_continue = tmp_channel_full_n;

assign tdf2_accum_2_U0_ap_start = accum1_out_0_t_empty_n;

assign tdf2_accum_2_U0_start_full_n = 1'b1;

assign tdf2_accum_2_U0_start_write = 1'b0;

assign tdf2_adjust_U0_ap_continue = outputs_0_full_n;

assign tdf2_adjust_U0_ap_start = sums_0_empty_n;

assign tdf2_adjust_U0_start_full_n = 1'b1;

assign tdf2_adjust_U0_start_write = 1'b0;

assign tdf2_dot_product_U0_ap_continue = products_0_i_full_n;

assign tdf2_dot_product_U0_ap_start = (weight_vecs_0_t_empty_n & ifmap_vec_t_empty_n);

assign tdf2_dot_product_U0_products_0_full_n = products_0_i_full_n;

assign tdf2_dot_product_U0_start_full_n = 1'b1;

assign tdf2_dot_product_U0_start_write = 1'b0;

assign tdf2_get_next_ijk_U0_ap_continue = (ap_sync_channel_write_input_indices_1 & ap_sync_channel_write_input_indices_0);

assign tdf2_get_next_ijk_U0_ap_start = ((ap_sync_reg_tdf2_get_next_ijk_U0_ap_ready ^ 1'b1) & ap_start);

assign tdf2_poolOutputs_U0_ap_continue = ap_continue;

assign tdf2_poolOutputs_U0_ap_start = outputs_0_empty_n;

assign tdf2_poolOutputs_U0_out_data_full_n = out_data_full_n;

assign tdf2_poolOutputs_U0_out_data_write = 1'b0;

assign tdf2_poolOutputs_U0_start_full_n = 1'b1;

assign tdf2_poolOutputs_U0_start_write = 1'b0;

assign tdf2_readFilters24_U0_ap_continue = weight_vecs_0_i_full_n;

assign tdf2_readFilters24_U0_ap_start = start_for_tdf2_readFilters24_U0_empty_n;

assign tdf2_readFilters24_U0_start_full_n = 1'b1;

assign tdf2_readFilters24_U0_start_write = 1'b0;

assign tdf2_readFilters24_U0_weight_vecs_0_full_n = weight_vecs_0_i_full_n;

assign tdf2_readInputs25_U0_ap_continue = ifmap_vec_i_full_n;

assign tdf2_readInputs25_U0_ap_start = (input_indices_1_empty_n & input_indices_0_empty_n & (ap_sync_reg_tdf2_readInputs25_U0_ap_ready ^ 1'b1) & ap_start);

assign tdf2_readInputs25_U0_ifmap_vec_full_n = ifmap_vec_i_full_n;

assign tdf2_readInputs25_U0_in_data_full_n = in_data_empty_n;

assign tdf2_readInputs25_U0_in_data_write = 1'b0;

assign tdf2_readInputs25_U0_start_full_n = 1'b1;

assign tdf2_readInputs25_U0_start_write = 1'b0;

endmodule //td_fused_top_dataflow_in_loop_TOP_LOOP38022
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP38022_weight_vecs_0_memcore_ram (addr0, ce0, d0, we0, q0, addr1, ce1, d1, we1, q1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 9;
parameter MEM_SIZE = 288;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
output reg[DWIDTH-1:0] q1;
input clk;

reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];




always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1) 
            ram[addr1] <= d1; 
        q1 <= ram[addr1];
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP38022_weight_vecs_0_memcore(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    q0,
    address1,
    ce1,
    we1,
    d1,
    q1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd288;
parameter AddressWidth = 32'd9;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;
output[DataWidth - 1:0] q1;



td_fused_top_dataflow_in_loop_TOP_LOOP38022_weight_vecs_0_memcore_ram td_fused_top_dataflow_in_loop_TOP_LOOP38022_weight_vecs_0_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 ),
    .q1( q1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_dataflow_in_loop_TOP_LOOP38022_weight_vecs_0
#(parameter
    DataWidth    = 16,
    AddressRange = 32,
    AddressWidth = 8,
    BufferCount  = 2,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire                    i_we0,
    input  wire [AddressWidth-1:0] i_address0,
    input  wire [DataWidth-1:0]    i_d0,
    output wire [DataWidth-1:0]    i_q0,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire                    t_we0,
    input  wire [AddressWidth-1:0] t_address0,
    input  wire [DataWidth-1:0]    t_d0,
    output wire [DataWidth-1:0]    t_q0
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
wire [AddressWidth+IndexWidth-1:0]   memcore_iaddr;
wire [AddressWidth+IndexWidth-1:0]   memcore_taddr;

//------------------------Instantiation------------------
assign memcore_iaddr = {i_address0, iptr};
assign memcore_taddr = {t_address0, tptr};
td_fused_top_dataflow_in_loop_TOP_LOOP38022_weight_vecs_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP38022_weight_vecs_0_memcore_U (
    .reset    ( reset ),
    .clk      ( clk ),
    .address0 ( memcore_iaddr ),
    .ce0      ( i_ce0 ),
    .we0      ( i_we0),
    .d0       ( i_d0 ),
    .q0       ( i_q0 ),
    .address1 ( memcore_taddr ),
    .ce1      ( t_ce0 ),
    .we1      ( t_we0),
    .d1       ( t_d0 ),
    .q1       ( t_q0 )

);

//------------------------Body---------------------------

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP38116_accum1_out_0_memcore_ram (addr0, ce0, d0, we0, q0, addr1, ce1, q1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 14;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
output reg[DWIDTH-1:0] q1;
input clk;

reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];




always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        q1 <= ram[addr1];
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP38116_accum1_out_0_memcore(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    q0,
    address1,
    ce1,
    q1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd14;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
output[DataWidth - 1:0] q1;



td_fused_top_dataflow_in_loop_TOP_LOOP38116_accum1_out_0_memcore_ram td_fused_top_dataflow_in_loop_TOP_LOOP38116_accum1_out_0_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .q1( q1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_dataflow_in_loop_TOP_LOOP38116_accum1_out_0
#(parameter
    DataWidth    = 16,
    AddressRange = 32,
    AddressWidth = 4,
    BufferCount  = 2,
    MemLatency   = 1,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire                    i_we0,
    input  wire [AddressWidth-1:0] i_address0,
    input  wire [DataWidth-1:0]    i_d0,
    output wire [DataWidth-1:0]    i_q0,
    input  wire                    i_ce1,
    input  wire [AddressWidth-1:0] i_address1,
    output wire [DataWidth-1:0]    i_q1,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire                    t_we0,
    input  wire [AddressWidth-1:0] t_address0,
    input  wire [DataWidth-1:0]    t_d0,
    output wire [DataWidth-1:0]    t_q0,
    input  wire                    t_ce1,
    input  wire [AddressWidth-1:0] t_address1,
    output wire [DataWidth-1:0]    t_q1
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth-1:0]   prev_iptr    = 1'b0; // previous initiator index
reg  [IndexWidth-1:0]   prev_tptr    = 1'b0; // previous target index
reg  [DataWidth-1:0]    reg_q0      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid0    = 1'b0; // buffer has valid data
reg  [DataWidth-1:0]    reg_q1      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid1    = 1'b0; // buffer has valid data
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
// buffer signals
wire [BufferCount-1:0] buf_ce0;
wire [BufferCount-1:0] buf_we0;
wire [AddressWidth-1:0] buf_a0_0, buf_a0_1;
wire [DataWidth-1:0] buf_d0_0, buf_d0_1;
wire [DataWidth-1:0] buf_q0_0, buf_q0_1;
wire [BufferCount-1:0] buf_ce1;
wire [AddressWidth-1:0] buf_a1_0, buf_a1_1;
wire [DataWidth-1:0] buf_q1_0, buf_q1_1;
//------------------------Instantiation------------------
//genvar i;
        td_fused_top_dataflow_in_loop_TOP_LOOP38116_accum1_out_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP38116_accum1_out_0_memcore_U_0 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_0 ),
            .ce0      ( buf_ce0[ 0 ] ),
            .we0      ( buf_we0[ 0 ] ),
            .d0       ( buf_d0_0 ),
            .q0       ( buf_q0_0 ),
            .address1 ( buf_a1_0 ),
            .ce1      ( buf_ce1[ 0 ] ),
            .q1       ( buf_q1_0 )
        );
        td_fused_top_dataflow_in_loop_TOP_LOOP38116_accum1_out_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP38116_accum1_out_0_memcore_U_1 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_1 ),
            .ce0      ( buf_ce0[ 1 ] ),
            .we0      ( buf_we0[ 1 ] ),
            .d0       ( buf_d0_1 ),
            .q0       ( buf_q0_1 ),
            .address1 ( buf_a1_1 ),
            .ce1      ( buf_ce1[ 1 ] ),
            .q1       ( buf_q1_1 )
        );

//++++++++++++++++++++++++buffer signals+++++++++++++++++
        assign buf_ce0[ 0 ] = (tptr ==  0  && empty_n) ? t_ce0
                             : (iptr ==  0 ) ? i_ce0 : 1'b0;
        assign buf_a0_0  = (tptr ==  0  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 0 ] = (tptr ==  0  && empty_n)  ? t_we0
                             : (iptr ==  0 ) ? i_we0 : 1'b0;
        assign buf_d0_0  = (tptr ==  0  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 0 ] = (tptr ==  0  && empty_n) ? t_ce1
                             : (iptr ==  0 ) ? i_ce1 : 1'b0;
        assign buf_a1_0  = (tptr ==  0  && empty_n) ?  t_address1 : i_address1;
        assign buf_ce0[ 1 ] = (tptr ==  1  && empty_n) ? t_ce0
                             : (iptr ==  1 ) ? i_ce0 : 1'b0;
        assign buf_a0_1  = (tptr ==  1  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 1 ] = (tptr ==  1  && empty_n)  ? t_we0
                             : (iptr ==  1 ) ? i_we0 : 1'b0;
        assign buf_d0_1  = (tptr ==  1  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 1 ] = (tptr ==  1  && empty_n) ? t_ce1
                             : (iptr ==  1 ) ? i_ce1 : 1'b0;
        assign buf_a1_1  = (tptr ==  1  && empty_n) ?  t_address1 : i_address1;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//------------------------Body---------------------------
assign i_q0      = (prev_iptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign t_q0      = reg_valid0 ? reg_q0 : (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign i_q1      = (prev_iptr == 1'b1 ? buf_q1_1 : buf_q1_0);
assign t_q1      = reg_valid1 ? reg_q1 : (prev_tptr == 1'b1 ? buf_q1_1 : buf_q1_0);

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// prev_iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_iptr <= 1'b0;
    else begin
        prev_iptr <= iptr;
    end
end

// prev_tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_tptr <= 1'b0;
    else begin
        prev_tptr <= tptr;
    end
end

// reg_q0 and reg_valid0
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q0     <= 1'b0;
        reg_valid0 <= 1'b0;
    end else if (!t_ce0 && !reg_valid0) begin
        reg_q0     <= (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
        reg_valid0 <= 1'b1;
    end else if (t_ce0) begin
        reg_valid0 <= 1'b0;
    end
end

// reg_q1 and reg_valid1
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q1     <= 1'b0;
        reg_valid1 <= 1'b0;
    end else if (!t_ce1 && !reg_valid1) begin
        reg_q1     <= (prev_tptr == 1'b1 ? buf_q1_1 : buf_q1_0);
        reg_valid1 <= 1'b1;
    end else if (t_ce1) begin
        reg_valid1 <= 1'b0;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP38116_accum2_out_0_memcore_ram (addr0, ce0, d0, we0, q0, addr1, ce1, d1, we1, q1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 14;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
output reg[DWIDTH-1:0] q1;
input clk;

reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];




always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1) 
            ram[addr1] <= d1; 
        q1 <= ram[addr1];
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP38116_accum2_out_0_memcore(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    q0,
    address1,
    ce1,
    we1,
    d1,
    q1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd14;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;
output[DataWidth - 1:0] q1;



td_fused_top_dataflow_in_loop_TOP_LOOP38116_accum2_out_0_memcore_ram td_fused_top_dataflow_in_loop_TOP_LOOP38116_accum2_out_0_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 ),
    .q1( q1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_dataflow_in_loop_TOP_LOOP38116_accum2_out_0
#(parameter
    DataWidth    = 16,
    AddressRange = 32,
    AddressWidth = 3,
    BufferCount  = 2,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire                    i_we0,
    input  wire [AddressWidth-1:0] i_address0,
    input  wire [DataWidth-1:0]    i_d0,
    output wire [DataWidth-1:0]    i_q0,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire                    t_we0,
    input  wire [AddressWidth-1:0] t_address0,
    input  wire [DataWidth-1:0]    t_d0,
    output wire [DataWidth-1:0]    t_q0
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
wire [AddressWidth+IndexWidth-1:0]   memcore_iaddr;
wire [AddressWidth+IndexWidth-1:0]   memcore_taddr;

//------------------------Instantiation------------------
assign memcore_iaddr = {i_address0, iptr};
assign memcore_taddr = {t_address0, tptr};
td_fused_top_dataflow_in_loop_TOP_LOOP38116_accum2_out_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP38116_accum2_out_0_memcore_U (
    .reset    ( reset ),
    .clk      ( clk ),
    .address0 ( memcore_iaddr ),
    .ce0      ( i_ce0 ),
    .we0      ( i_we0),
    .d0       ( i_d0 ),
    .q0       ( i_q0 ),
    .address1 ( memcore_taddr ),
    .ce1      ( t_ce0 ),
    .we1      ( t_we0),
    .d1       ( t_d0 ),
    .q1       ( t_q0 )

);

//------------------------Body---------------------------

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP38116_ifmap_vec_memcore_ram (addr0, ce0, d0, we0, q0, addr1, ce1, d1, we1, q1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 6;
parameter MEM_SIZE = 54;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
output reg[DWIDTH-1:0] q1;
input clk;

reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];




always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1) 
            ram[addr1] <= d1; 
        q1 <= ram[addr1];
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP38116_ifmap_vec_memcore(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    q0,
    address1,
    ce1,
    we1,
    d1,
    q1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd54;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;
output[DataWidth - 1:0] q1;



td_fused_top_dataflow_in_loop_TOP_LOOP38116_ifmap_vec_memcore_ram td_fused_top_dataflow_in_loop_TOP_LOOP38116_ifmap_vec_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 ),
    .q1( q1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_dataflow_in_loop_TOP_LOOP38116_ifmap_vec
#(parameter
    DataWidth    = 16,
    AddressRange = 32,
    AddressWidth = 5,
    BufferCount  = 2,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire                    i_we0,
    input  wire [AddressWidth-1:0] i_address0,
    input  wire [DataWidth-1:0]    i_d0,
    output wire [DataWidth-1:0]    i_q0,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire                    t_we0,
    input  wire [AddressWidth-1:0] t_address0,
    input  wire [DataWidth-1:0]    t_d0,
    output wire [DataWidth-1:0]    t_q0
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
wire [AddressWidth+IndexWidth-1:0]   memcore_iaddr;
wire [AddressWidth+IndexWidth-1:0]   memcore_taddr;

//------------------------Instantiation------------------
assign memcore_iaddr = {i_address0, iptr};
assign memcore_taddr = {t_address0, tptr};
td_fused_top_dataflow_in_loop_TOP_LOOP38116_ifmap_vec_memcore td_fused_top_dataflow_in_loop_TOP_LOOP38116_ifmap_vec_memcore_U (
    .reset    ( reset ),
    .clk      ( clk ),
    .address0 ( memcore_iaddr ),
    .ce0      ( i_ce0 ),
    .we0      ( i_we0),
    .d0       ( i_d0 ),
    .q0       ( i_q0 ),
    .address1 ( memcore_taddr ),
    .ce1      ( t_ce0 ),
    .we1      ( t_we0),
    .d1       ( t_d0 ),
    .q1       ( t_q0 )

);

//------------------------Body---------------------------

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP38116_products_0_memcore_ram (addr0, ce0, d0, we0, q0, addr1, ce1, q1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 5;
parameter MEM_SIZE = 27;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
output reg[DWIDTH-1:0] q1;
input clk;

reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];




always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        q1 <= ram[addr1];
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP38116_products_0_memcore(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    q0,
    address1,
    ce1,
    q1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd27;
parameter AddressWidth = 32'd5;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
output[DataWidth - 1:0] q1;



td_fused_top_dataflow_in_loop_TOP_LOOP38116_products_0_memcore_ram td_fused_top_dataflow_in_loop_TOP_LOOP38116_products_0_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .q1( q1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_dataflow_in_loop_TOP_LOOP38116_products_0
#(parameter
    DataWidth    = 16,
    AddressRange = 32,
    AddressWidth = 5,
    BufferCount  = 2,
    MemLatency   = 1,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire                    i_we0,
    input  wire [AddressWidth-1:0] i_address0,
    input  wire [DataWidth-1:0]    i_d0,
    output wire [DataWidth-1:0]    i_q0,
    input  wire                    i_ce1,
    input  wire [AddressWidth-1:0] i_address1,
    output wire [DataWidth-1:0]    i_q1,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire                    t_we0,
    input  wire [AddressWidth-1:0] t_address0,
    input  wire [DataWidth-1:0]    t_d0,
    output wire [DataWidth-1:0]    t_q0,
    input  wire                    t_ce1,
    input  wire [AddressWidth-1:0] t_address1,
    output wire [DataWidth-1:0]    t_q1
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth-1:0]   prev_iptr    = 1'b0; // previous initiator index
reg  [IndexWidth-1:0]   prev_tptr    = 1'b0; // previous target index
reg  [DataWidth-1:0]    reg_q0      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid0    = 1'b0; // buffer has valid data
reg  [DataWidth-1:0]    reg_q1      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid1    = 1'b0; // buffer has valid data
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
// buffer signals
wire [BufferCount-1:0] buf_ce0;
wire [BufferCount-1:0] buf_we0;
wire [AddressWidth-1:0] buf_a0_0, buf_a0_1;
wire [DataWidth-1:0] buf_d0_0, buf_d0_1;
wire [DataWidth-1:0] buf_q0_0, buf_q0_1;
wire [BufferCount-1:0] buf_ce1;
wire [AddressWidth-1:0] buf_a1_0, buf_a1_1;
wire [DataWidth-1:0] buf_q1_0, buf_q1_1;
//------------------------Instantiation------------------
//genvar i;
        td_fused_top_dataflow_in_loop_TOP_LOOP38116_products_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP38116_products_0_memcore_U_0 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_0 ),
            .ce0      ( buf_ce0[ 0 ] ),
            .we0      ( buf_we0[ 0 ] ),
            .d0       ( buf_d0_0 ),
            .q0       ( buf_q0_0 ),
            .address1 ( buf_a1_0 ),
            .ce1      ( buf_ce1[ 0 ] ),
            .q1       ( buf_q1_0 )
        );
        td_fused_top_dataflow_in_loop_TOP_LOOP38116_products_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP38116_products_0_memcore_U_1 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_1 ),
            .ce0      ( buf_ce0[ 1 ] ),
            .we0      ( buf_we0[ 1 ] ),
            .d0       ( buf_d0_1 ),
            .q0       ( buf_q0_1 ),
            .address1 ( buf_a1_1 ),
            .ce1      ( buf_ce1[ 1 ] ),
            .q1       ( buf_q1_1 )
        );

//++++++++++++++++++++++++buffer signals+++++++++++++++++
        assign buf_ce0[ 0 ] = (tptr ==  0  && empty_n) ? t_ce0
                             : (iptr ==  0 ) ? i_ce0 : 1'b0;
        assign buf_a0_0  = (tptr ==  0  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 0 ] = (tptr ==  0  && empty_n)  ? t_we0
                             : (iptr ==  0 ) ? i_we0 : 1'b0;
        assign buf_d0_0  = (tptr ==  0  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 0 ] = (tptr ==  0  && empty_n) ? t_ce1
                             : (iptr ==  0 ) ? i_ce1 : 1'b0;
        assign buf_a1_0  = (tptr ==  0  && empty_n) ?  t_address1 : i_address1;
        assign buf_ce0[ 1 ] = (tptr ==  1  && empty_n) ? t_ce0
                             : (iptr ==  1 ) ? i_ce0 : 1'b0;
        assign buf_a0_1  = (tptr ==  1  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 1 ] = (tptr ==  1  && empty_n)  ? t_we0
                             : (iptr ==  1 ) ? i_we0 : 1'b0;
        assign buf_d0_1  = (tptr ==  1  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 1 ] = (tptr ==  1  && empty_n) ? t_ce1
                             : (iptr ==  1 ) ? i_ce1 : 1'b0;
        assign buf_a1_1  = (tptr ==  1  && empty_n) ?  t_address1 : i_address1;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//------------------------Body---------------------------
assign i_q0      = (prev_iptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign t_q0      = reg_valid0 ? reg_q0 : (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign i_q1      = (prev_iptr == 1'b1 ? buf_q1_1 : buf_q1_0);
assign t_q1      = reg_valid1 ? reg_q1 : (prev_tptr == 1'b1 ? buf_q1_1 : buf_q1_0);

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// prev_iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_iptr <= 1'b0;
    else begin
        prev_iptr <= iptr;
    end
end

// prev_tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_tptr <= 1'b0;
    else begin
        prev_tptr <= tptr;
    end
end

// reg_q0 and reg_valid0
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q0     <= 1'b0;
        reg_valid0 <= 1'b0;
    end else if (!t_ce0 && !reg_valid0) begin
        reg_q0     <= (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
        reg_valid0 <= 1'b1;
    end else if (t_ce0) begin
        reg_valid0 <= 1'b0;
    end
end

// reg_q1 and reg_valid1
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q1     <= 1'b0;
        reg_valid1 <= 1'b0;
    end else if (!t_ce1 && !reg_valid1) begin
        reg_q1     <= (prev_tptr == 1'b1 ? buf_q1_1 : buf_q1_0);
        reg_valid1 <= 1'b1;
    end else if (t_ce1) begin
        reg_valid1 <= 1'b0;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_dataflow_in_loop_TOP_LOOP38116 (
        ap_clk,
        ap_rst,
        in_data_address0,
        in_data_ce0,
        in_data_d0,
        in_data_q0,
        in_data_we0,
        in_data_address1,
        in_data_ce1,
        in_data_d1,
        in_data_q1,
        in_data_we1,
        filter_data_address0,
        filter_data_ce0,
        filter_data_d0,
        filter_data_q0,
        filter_data_we0,
        filter_data_address1,
        filter_data_ce1,
        filter_data_d1,
        filter_data_q1,
        filter_data_we1,
        adjustments_address0,
        adjustments_ce0,
        adjustments_d0,
        adjustments_q0,
        adjustments_we0,
        adjustments_address1,
        adjustments_ce1,
        adjustments_d1,
        adjustments_q1,
        adjustments_we1,
        out_data_address0,
        out_data_ce0,
        out_data_d0,
        out_data_q0,
        out_data_we0,
        out_data_address1,
        out_data_ce1,
        out_data_d1,
        out_data_q1,
        out_data_we1,
        ap_start,
        in_data_empty_n,
        in_data_read,
        out_data_full_n,
        out_data_write,
        ap_done,
        ap_ready,
        ap_idle,
        ap_continue
);


input   ap_clk;
input   ap_rst;
output  [15:0] in_data_address0;
output   in_data_ce0;
output  [63:0] in_data_d0;
input  [63:0] in_data_q0;
output   in_data_we0;
output  [15:0] in_data_address1;
output   in_data_ce1;
output  [63:0] in_data_d1;
input  [63:0] in_data_q1;
output   in_data_we1;
output  [8:0] filter_data_address0;
output   filter_data_ce0;
output  [15:0] filter_data_d0;
input  [15:0] filter_data_q0;
output   filter_data_we0;
output  [8:0] filter_data_address1;
output   filter_data_ce1;
output  [15:0] filter_data_d1;
input  [15:0] filter_data_q1;
output   filter_data_we1;
output  [3:0] adjustments_address0;
output   adjustments_ce0;
output  [47:0] adjustments_d0;
input  [47:0] adjustments_q0;
output   adjustments_we0;
output  [3:0] adjustments_address1;
output   adjustments_ce1;
output  [47:0] adjustments_d1;
input  [47:0] adjustments_q1;
output   adjustments_we1;
output  [15:0] out_data_address0;
output   out_data_ce0;
output  [63:0] out_data_d0;
input  [63:0] out_data_q0;
output   out_data_we0;
output  [15:0] out_data_address1;
output   out_data_ce1;
output  [63:0] out_data_d1;
input  [63:0] out_data_q1;
output   out_data_we1;
input   ap_start;
input   in_data_empty_n;
output   in_data_read;
input   out_data_full_n;
output   out_data_write;
output   ap_done;
output   ap_ready;
output   ap_idle;
input   ap_continue;

wire   [15:0] ifmap_vec_i_q0;
wire   [15:0] ifmap_vec_t_q0;
wire   [15:0] weight_vecs_0_i_q0;
wire   [15:0] weight_vecs_0_t_q0;
wire   [15:0] products_0_i_q0;
wire   [15:0] products_0_i_q1;
wire   [15:0] products_0_t_q0;
wire   [15:0] products_0_t_q1;
wire   [15:0] accum1_out_0_i_q0;
wire   [15:0] accum1_out_0_i_q1;
wire   [15:0] accum1_out_0_t_q0;
wire   [15:0] accum1_out_0_t_q1;
wire   [15:0] accum2_out_0_i_q0;
wire   [15:0] accum2_out_0_t_q0;
wire    tdf1_get_next_ijk_U0_ap_start;
wire    tdf1_get_next_ijk_U0_ap_done;
wire    tdf1_get_next_ijk_U0_ap_continue;
wire    tdf1_get_next_ijk_U0_ap_idle;
wire    tdf1_get_next_ijk_U0_ap_ready;
wire    tdf1_get_next_ijk_U0_start_out;
wire    tdf1_get_next_ijk_U0_start_write;
wire   [3:0] tdf1_get_next_ijk_U0_input_indices_2_out_din;
wire    tdf1_get_next_ijk_U0_input_indices_2_out_write;
wire   [3:0] tdf1_get_next_ijk_U0_input_indices_2_out1_din;
wire    tdf1_get_next_ijk_U0_input_indices_2_out1_write;
wire   [6:0] tdf1_get_next_ijk_U0_output_indices_0_din;
wire    tdf1_get_next_ijk_U0_output_indices_0_write;
wire   [13:0] tdf1_get_next_ijk_U0_output_indices_1_din;
wire    tdf1_get_next_ijk_U0_output_indices_1_write;
wire    tdf1_get_next_ijk_U0_resetMaximum_din;
wire    tdf1_get_next_ijk_U0_resetMaximum_write;
wire    tdf1_get_next_ijk_U0_storeOutput_din;
wire    tdf1_get_next_ijk_U0_storeOutput_write;
wire   [15:0] tdf1_get_next_ijk_U0_ap_return_0;
wire   [15:0] tdf1_get_next_ijk_U0_ap_return_1;
wire    ap_channel_done_input_indices_1;
wire    input_indices_1_full_n;
reg    ap_sync_reg_channel_write_input_indices_1;
wire    ap_sync_channel_write_input_indices_1;
wire    ap_channel_done_input_indices_0;
wire    input_indices_0_full_n;
reg    ap_sync_reg_channel_write_input_indices_0;
wire    ap_sync_channel_write_input_indices_0;
wire    tdf1_readInputs19_U0_ap_start;
wire    tdf1_readInputs19_U0_ap_done;
wire    tdf1_readInputs19_U0_ap_continue;
wire    tdf1_readInputs19_U0_ap_idle;
wire    tdf1_readInputs19_U0_ap_ready;
wire   [15:0] tdf1_readInputs19_U0_in_data_address0;
wire    tdf1_readInputs19_U0_in_data_ce0;
wire   [4:0] tdf1_readInputs19_U0_ifmap_vec_address0;
wire    tdf1_readInputs19_U0_ifmap_vec_ce0;
wire    tdf1_readInputs19_U0_ifmap_vec_we0;
wire   [15:0] tdf1_readInputs19_U0_ifmap_vec_d0;
wire    tdf1_readInputs19_U0_in_data_full_n;
wire    tdf1_readInputs19_U0_in_data_write;
wire    ap_channel_done_ifmap_vec;
wire    tdf1_readInputs19_U0_ifmap_vec_full_n;
wire    tdf1_readFilters18_U0_ap_start;
wire    tdf1_readFilters18_U0_ap_done;
wire    tdf1_readFilters18_U0_ap_continue;
wire    tdf1_readFilters18_U0_ap_idle;
wire    tdf1_readFilters18_U0_ap_ready;
wire   [8:0] tdf1_readFilters18_U0_filter_data_address0;
wire    tdf1_readFilters18_U0_filter_data_ce0;
wire    tdf1_readFilters18_U0_input_indices_23_read;
wire   [4:0] tdf1_readFilters18_U0_weight_vecs_0_address0;
wire    tdf1_readFilters18_U0_weight_vecs_0_ce0;
wire    tdf1_readFilters18_U0_weight_vecs_0_we0;
wire   [15:0] tdf1_readFilters18_U0_weight_vecs_0_d0;
wire    ap_channel_done_weight_vecs_0;
wire    tdf1_readFilters18_U0_weight_vecs_0_full_n;
wire    tdf1_dot_product_U0_ap_start;
wire    tdf1_dot_product_U0_ap_done;
wire    tdf1_dot_product_U0_ap_continue;
wire    tdf1_dot_product_U0_ap_idle;
wire    tdf1_dot_product_U0_ap_ready;
wire   [4:0] tdf1_dot_product_U0_ifmap_vec_address0;
wire    tdf1_dot_product_U0_ifmap_vec_ce0;
wire   [4:0] tdf1_dot_product_U0_weight_vecs_0_address0;
wire    tdf1_dot_product_U0_weight_vecs_0_ce0;
wire   [4:0] tdf1_dot_product_U0_products_0_address0;
wire    tdf1_dot_product_U0_products_0_ce0;
wire    tdf1_dot_product_U0_products_0_we0;
wire   [15:0] tdf1_dot_product_U0_products_0_d0;
wire    ap_channel_done_products_0;
wire    tdf1_dot_product_U0_products_0_full_n;
wire    tdf1_accum_1_U0_ap_start;
wire    tdf1_accum_1_U0_ap_done;
wire    tdf1_accum_1_U0_ap_continue;
wire    tdf1_accum_1_U0_ap_idle;
wire    tdf1_accum_1_U0_ap_ready;
wire   [4:0] tdf1_accum_1_U0_accum_in_0_address0;
wire    tdf1_accum_1_U0_accum_in_0_ce0;
wire   [4:0] tdf1_accum_1_U0_accum_in_0_address1;
wire    tdf1_accum_1_U0_accum_in_0_ce1;
wire   [3:0] tdf1_accum_1_U0_accum_out_address0;
wire    tdf1_accum_1_U0_accum_out_ce0;
wire    tdf1_accum_1_U0_accum_out_we0;
wire   [15:0] tdf1_accum_1_U0_accum_out_d0;
wire    ap_channel_done_accum1_out_0;
wire    tdf1_accum_1_U0_accum_out_full_n;
wire    tdf1_accum_2_U0_ap_start;
wire    tdf1_accum_2_U0_ap_done;
wire    tdf1_accum_2_U0_ap_continue;
wire    tdf1_accum_2_U0_ap_idle;
wire    tdf1_accum_2_U0_ap_ready;
wire   [3:0] tdf1_accum_2_U0_accum_in_address0;
wire    tdf1_accum_2_U0_accum_in_ce0;
wire   [3:0] tdf1_accum_2_U0_accum_in_address1;
wire    tdf1_accum_2_U0_accum_in_ce1;
wire   [2:0] tdf1_accum_2_U0_accum_out_address0;
wire    tdf1_accum_2_U0_accum_out_ce0;
wire    tdf1_accum_2_U0_accum_out_we0;
wire   [15:0] tdf1_accum_2_U0_accum_out_d0;
wire    ap_channel_done_accum2_out_0;
wire    tdf1_accum_2_U0_accum_out_full_n;
wire    tdf1_accum_3_U0_ap_start;
wire    tdf1_accum_3_U0_ap_done;
wire    tdf1_accum_3_U0_ap_continue;
wire    tdf1_accum_3_U0_ap_idle;
wire    tdf1_accum_3_U0_ap_ready;
wire   [15:0] tdf1_accum_3_U0_accum_in_18;
wire    tdf1_accum_3_U0_accum_in_18_ap_vld;
wire   [2:0] tdf1_accum_3_U0_accum_in_address0;
wire    tdf1_accum_3_U0_accum_in_ce0;
wire    ap_channel_done_tmp_channel;
wire    tmp_channel_full_n;
wire    Block_entry_proc_proc_U0_ap_start;
wire    Block_entry_proc_proc_U0_ap_done;
wire    Block_entry_proc_proc_U0_ap_continue;
wire    Block_entry_proc_proc_U0_ap_idle;
wire    Block_entry_proc_proc_U0_ap_ready;
wire   [15:0] Block_entry_proc_proc_U0_ap_return;
wire    ap_channel_done_sums_0;
wire    sums_0_full_n;
wire    tdf1_adjust_U0_ap_start;
wire    tdf1_adjust_U0_ap_done;
wire    tdf1_adjust_U0_ap_continue;
wire    tdf1_adjust_U0_ap_idle;
wire    tdf1_adjust_U0_ap_ready;
wire   [3:0] tdf1_adjust_U0_adjustments_address0;
wire    tdf1_adjust_U0_adjustments_ce0;
wire    tdf1_adjust_U0_input_indices_23_read;
wire   [15:0] tdf1_adjust_U0_ap_return;
wire    ap_channel_done_outputs_0;
wire    outputs_0_full_n;
wire    tdf1_poolOutputs_U0_ap_start;
wire    tdf1_poolOutputs_U0_ap_done;
wire    tdf1_poolOutputs_U0_ap_continue;
wire    tdf1_poolOutputs_U0_ap_idle;
wire    tdf1_poolOutputs_U0_ap_ready;
wire    tdf1_poolOutputs_U0_output_indices_04_read;
wire    tdf1_poolOutputs_U0_output_indices_15_read;
wire    tdf1_poolOutputs_U0_resetMaximum6_read;
wire    tdf1_poolOutputs_U0_storeOutput7_read;
wire   [15:0] tdf1_poolOutputs_U0_out_data_address1;
wire    tdf1_poolOutputs_U0_out_data_ce1;
wire    tdf1_poolOutputs_U0_out_data_we1;
wire   [63:0] tdf1_poolOutputs_U0_out_data_d1;
wire    tdf1_poolOutputs_U0_out_data_full_n;
wire    tdf1_poolOutputs_U0_out_data_write;
wire    ap_sync_continue;
wire    ifmap_vec_i_full_n;
wire    ifmap_vec_t_empty_n;
wire    weight_vecs_0_i_full_n;
wire    weight_vecs_0_t_empty_n;
wire    products_0_i_full_n;
wire    products_0_t_empty_n;
wire   [15:0] products_0_t_d1;
wire    products_0_t_we1;
wire    accum1_out_0_i_full_n;
wire    accum1_out_0_t_empty_n;
wire   [15:0] accum1_out_0_t_d1;
wire    accum1_out_0_t_we1;
wire    accum2_out_0_i_full_n;
wire    accum2_out_0_t_empty_n;
wire    input_indices_23_c_full_n;
wire   [3:0] input_indices_23_c_dout;
wire    input_indices_23_c_empty_n;
wire    input_indices_23_c1_full_n;
wire   [3:0] input_indices_23_c1_dout;
wire    input_indices_23_c1_empty_n;
wire    output_indices_04_c_full_n;
wire   [6:0] output_indices_04_c_dout;
wire    output_indices_04_c_empty_n;
wire    output_indices_15_c_full_n;
wire   [13:0] output_indices_15_c_dout;
wire    output_indices_15_c_empty_n;
wire   [0:0] resetMaximum6_c_din;
wire    resetMaximum6_c_full_n;
wire   [0:0] resetMaximum6_c_dout;
wire    resetMaximum6_c_empty_n;
wire   [0:0] storeOutput7_c_din;
wire    storeOutput7_c_full_n;
wire   [0:0] storeOutput7_c_dout;
wire    storeOutput7_c_empty_n;
wire   [15:0] input_indices_0_dout;
wire    input_indices_0_empty_n;
wire   [15:0] input_indices_1_dout;
wire    input_indices_1_empty_n;
wire   [15:0] tmp_channel_dout;
wire    tmp_channel_empty_n;
wire   [15:0] sums_0_dout;
wire    sums_0_empty_n;
wire   [15:0] outputs_0_dout;
wire    outputs_0_empty_n;
wire    ap_sync_done;
wire    ap_sync_ready;
reg    ap_sync_reg_tdf1_get_next_ijk_U0_ap_ready;
wire    ap_sync_tdf1_get_next_ijk_U0_ap_ready;
reg    ap_sync_reg_tdf1_readInputs19_U0_ap_ready;
wire    ap_sync_tdf1_readInputs19_U0_ap_ready;
wire   [0:0] start_for_tdf1_readFilters18_U0_din;
wire    start_for_tdf1_readFilters18_U0_full_n;
wire   [0:0] start_for_tdf1_readFilters18_U0_dout;
wire    start_for_tdf1_readFilters18_U0_empty_n;
wire    tdf1_readInputs19_U0_start_full_n;
wire    tdf1_readInputs19_U0_start_write;
wire    tdf1_readFilters18_U0_start_full_n;
wire    tdf1_readFilters18_U0_start_write;
wire    tdf1_dot_product_U0_start_full_n;
wire    tdf1_dot_product_U0_start_write;
wire    tdf1_accum_1_U0_start_full_n;
wire    tdf1_accum_1_U0_start_write;
wire    tdf1_accum_2_U0_start_full_n;
wire    tdf1_accum_2_U0_start_write;
wire    tdf1_accum_3_U0_start_full_n;
wire    tdf1_accum_3_U0_start_write;
wire    Block_entry_proc_proc_U0_start_full_n;
wire    Block_entry_proc_proc_U0_start_write;
wire    tdf1_adjust_U0_start_full_n;
wire    tdf1_adjust_U0_start_write;
wire    tdf1_poolOutputs_U0_start_full_n;
wire    tdf1_poolOutputs_U0_start_write;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_sync_reg_channel_write_input_indices_1 = 1'b0;
#0 ap_sync_reg_channel_write_input_indices_0 = 1'b0;
#0 ap_sync_reg_tdf1_get_next_ijk_U0_ap_ready = 1'b0;
#0 ap_sync_reg_tdf1_readInputs19_U0_ap_ready = 1'b0;
end

td_fused_top_dataflow_in_loop_TOP_LOOP38116_ifmap_vec #(
    .DataWidth( 16 ),
    .AddressRange( 27 ),
    .AddressWidth( 5 ))
ifmap_vec_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf1_readInputs19_U0_ap_done),
    .i_full_n(ifmap_vec_i_full_n),
    .i_ce0(tdf1_readInputs19_U0_ifmap_vec_ce0),
    .i_we0(tdf1_readInputs19_U0_ifmap_vec_we0),
    .i_address0(tdf1_readInputs19_U0_ifmap_vec_address0),
    .i_d0(tdf1_readInputs19_U0_ifmap_vec_d0),
    .i_q0(ifmap_vec_i_q0),
    .t_ce(1'b1),
    .t_read(tdf1_dot_product_U0_ap_ready),
    .t_empty_n(ifmap_vec_t_empty_n),
    .t_ce0(tdf1_dot_product_U0_ifmap_vec_ce0),
    .t_we0(1'b0),
    .t_address0(tdf1_dot_product_U0_ifmap_vec_address0),
    .t_d0(16'd0),
    .t_q0(ifmap_vec_t_q0)
);

td_fused_top_dataflow_in_loop_TOP_LOOP38116_ifmap_vec #(
    .DataWidth( 16 ),
    .AddressRange( 27 ),
    .AddressWidth( 5 ))
weight_vecs_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf1_readFilters18_U0_ap_done),
    .i_full_n(weight_vecs_0_i_full_n),
    .i_ce0(tdf1_readFilters18_U0_weight_vecs_0_ce0),
    .i_we0(tdf1_readFilters18_U0_weight_vecs_0_we0),
    .i_address0(tdf1_readFilters18_U0_weight_vecs_0_address0),
    .i_d0(tdf1_readFilters18_U0_weight_vecs_0_d0),
    .i_q0(weight_vecs_0_i_q0),
    .t_ce(1'b1),
    .t_read(tdf1_dot_product_U0_ap_ready),
    .t_empty_n(weight_vecs_0_t_empty_n),
    .t_ce0(tdf1_dot_product_U0_weight_vecs_0_ce0),
    .t_we0(1'b0),
    .t_address0(tdf1_dot_product_U0_weight_vecs_0_address0),
    .t_d0(16'd0),
    .t_q0(weight_vecs_0_t_q0)
);

td_fused_top_dataflow_in_loop_TOP_LOOP38116_products_0 #(
    .DataWidth( 16 ),
    .AddressRange( 27 ),
    .AddressWidth( 5 ))
products_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf1_dot_product_U0_ap_done),
    .i_full_n(products_0_i_full_n),
    .i_ce0(tdf1_dot_product_U0_products_0_ce0),
    .i_we0(tdf1_dot_product_U0_products_0_we0),
    .i_address0(tdf1_dot_product_U0_products_0_address0),
    .i_d0(tdf1_dot_product_U0_products_0_d0),
    .i_q0(products_0_i_q0),
    .i_ce1(1'b0),
    .i_address1(5'd0),
    .i_q1(products_0_i_q1),
    .t_ce(1'b1),
    .t_read(tdf1_accum_1_U0_ap_ready),
    .t_empty_n(products_0_t_empty_n),
    .t_ce0(tdf1_accum_1_U0_accum_in_0_ce0),
    .t_we0(1'b0),
    .t_address0(tdf1_accum_1_U0_accum_in_0_address0),
    .t_d0(16'd0),
    .t_q0(products_0_t_q0),
    .t_ce1(tdf1_accum_1_U0_accum_in_0_ce1),
    .t_address1(tdf1_accum_1_U0_accum_in_0_address1),
    .t_q1(products_0_t_q1)
);

td_fused_top_dataflow_in_loop_TOP_LOOP38116_accum1_out_0 #(
    .DataWidth( 16 ),
    .AddressRange( 14 ),
    .AddressWidth( 4 ))
accum1_out_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf1_accum_1_U0_ap_done),
    .i_full_n(accum1_out_0_i_full_n),
    .i_ce0(tdf1_accum_1_U0_accum_out_ce0),
    .i_we0(tdf1_accum_1_U0_accum_out_we0),
    .i_address0(tdf1_accum_1_U0_accum_out_address0),
    .i_d0(tdf1_accum_1_U0_accum_out_d0),
    .i_q0(accum1_out_0_i_q0),
    .i_ce1(1'b0),
    .i_address1(4'd0),
    .i_q1(accum1_out_0_i_q1),
    .t_ce(1'b1),
    .t_read(tdf1_accum_2_U0_ap_ready),
    .t_empty_n(accum1_out_0_t_empty_n),
    .t_ce0(tdf1_accum_2_U0_accum_in_ce0),
    .t_we0(1'b0),
    .t_address0(tdf1_accum_2_U0_accum_in_address0),
    .t_d0(16'd0),
    .t_q0(accum1_out_0_t_q0),
    .t_ce1(tdf1_accum_2_U0_accum_in_ce1),
    .t_address1(tdf1_accum_2_U0_accum_in_address1),
    .t_q1(accum1_out_0_t_q1)
);

td_fused_top_dataflow_in_loop_TOP_LOOP38116_accum2_out_0 #(
    .DataWidth( 16 ),
    .AddressRange( 7 ),
    .AddressWidth( 3 ))
accum2_out_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf1_accum_2_U0_ap_done),
    .i_full_n(accum2_out_0_i_full_n),
    .i_ce0(tdf1_accum_2_U0_accum_out_ce0),
    .i_we0(tdf1_accum_2_U0_accum_out_we0),
    .i_address0(tdf1_accum_2_U0_accum_out_address0),
    .i_d0(tdf1_accum_2_U0_accum_out_d0),
    .i_q0(accum2_out_0_i_q0),
    .t_ce(1'b1),
    .t_read(tdf1_accum_3_U0_ap_ready),
    .t_empty_n(accum2_out_0_t_empty_n),
    .t_ce0(tdf1_accum_3_U0_accum_in_ce0),
    .t_we0(1'b0),
    .t_address0(tdf1_accum_3_U0_accum_in_address0),
    .t_d0(16'd0),
    .t_q0(accum2_out_0_t_q0)
);

td_fused_top_tdf1_get_next_ijk tdf1_get_next_ijk_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf1_get_next_ijk_U0_ap_start),
    .start_full_n(start_for_tdf1_readFilters18_U0_full_n),
    .ap_done(tdf1_get_next_ijk_U0_ap_done),
    .ap_continue(tdf1_get_next_ijk_U0_ap_continue),
    .ap_idle(tdf1_get_next_ijk_U0_ap_idle),
    .ap_ready(tdf1_get_next_ijk_U0_ap_ready),
    .start_out(tdf1_get_next_ijk_U0_start_out),
    .start_write(tdf1_get_next_ijk_U0_start_write),
    .input_indices_2_out_din(tdf1_get_next_ijk_U0_input_indices_2_out_din),
    .input_indices_2_out_full_n(input_indices_23_c_full_n),
    .input_indices_2_out_write(tdf1_get_next_ijk_U0_input_indices_2_out_write),
    .input_indices_2_out1_din(tdf1_get_next_ijk_U0_input_indices_2_out1_din),
    .input_indices_2_out1_full_n(input_indices_23_c1_full_n),
    .input_indices_2_out1_write(tdf1_get_next_ijk_U0_input_indices_2_out1_write),
    .output_indices_0_din(tdf1_get_next_ijk_U0_output_indices_0_din),
    .output_indices_0_full_n(output_indices_04_c_full_n),
    .output_indices_0_write(tdf1_get_next_ijk_U0_output_indices_0_write),
    .output_indices_1_din(tdf1_get_next_ijk_U0_output_indices_1_din),
    .output_indices_1_full_n(output_indices_15_c_full_n),
    .output_indices_1_write(tdf1_get_next_ijk_U0_output_indices_1_write),
    .resetMaximum_din(tdf1_get_next_ijk_U0_resetMaximum_din),
    .resetMaximum_full_n(resetMaximum6_c_full_n),
    .resetMaximum_write(tdf1_get_next_ijk_U0_resetMaximum_write),
    .storeOutput_din(tdf1_get_next_ijk_U0_storeOutput_din),
    .storeOutput_full_n(storeOutput7_c_full_n),
    .storeOutput_write(tdf1_get_next_ijk_U0_storeOutput_write),
    .ap_return_0(tdf1_get_next_ijk_U0_ap_return_0),
    .ap_return_1(tdf1_get_next_ijk_U0_ap_return_1)
);

td_fused_top_tdf1_readInputs19 tdf1_readInputs19_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf1_readInputs19_U0_ap_start),
    .ap_done(tdf1_readInputs19_U0_ap_done),
    .ap_continue(tdf1_readInputs19_U0_ap_continue),
    .ap_idle(tdf1_readInputs19_U0_ap_idle),
    .ap_ready(tdf1_readInputs19_U0_ap_ready),
    .in_data_address0(tdf1_readInputs19_U0_in_data_address0),
    .in_data_ce0(tdf1_readInputs19_U0_in_data_ce0),
    .in_data_q0(in_data_q0),
    .i_19(input_indices_0_dout),
    .j_19(input_indices_1_dout),
    .ifmap_vec_address0(tdf1_readInputs19_U0_ifmap_vec_address0),
    .ifmap_vec_ce0(tdf1_readInputs19_U0_ifmap_vec_ce0),
    .ifmap_vec_we0(tdf1_readInputs19_U0_ifmap_vec_we0),
    .ifmap_vec_d0(tdf1_readInputs19_U0_ifmap_vec_d0)
);

td_fused_top_tdf1_readFilters18 tdf1_readFilters18_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf1_readFilters18_U0_ap_start),
    .ap_done(tdf1_readFilters18_U0_ap_done),
    .ap_continue(tdf1_readFilters18_U0_ap_continue),
    .ap_idle(tdf1_readFilters18_U0_ap_idle),
    .ap_ready(tdf1_readFilters18_U0_ap_ready),
    .filter_data_address0(tdf1_readFilters18_U0_filter_data_address0),
    .filter_data_ce0(tdf1_readFilters18_U0_filter_data_ce0),
    .filter_data_q0(filter_data_q0),
    .input_indices_23_dout(input_indices_23_c_dout),
    .input_indices_23_empty_n(input_indices_23_c_empty_n),
    .input_indices_23_read(tdf1_readFilters18_U0_input_indices_23_read),
    .weight_vecs_0_address0(tdf1_readFilters18_U0_weight_vecs_0_address0),
    .weight_vecs_0_ce0(tdf1_readFilters18_U0_weight_vecs_0_ce0),
    .weight_vecs_0_we0(tdf1_readFilters18_U0_weight_vecs_0_we0),
    .weight_vecs_0_d0(tdf1_readFilters18_U0_weight_vecs_0_d0)
);

td_fused_top_tdf1_dot_product tdf1_dot_product_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf1_dot_product_U0_ap_start),
    .ap_done(tdf1_dot_product_U0_ap_done),
    .ap_continue(tdf1_dot_product_U0_ap_continue),
    .ap_idle(tdf1_dot_product_U0_ap_idle),
    .ap_ready(tdf1_dot_product_U0_ap_ready),
    .ifmap_vec_address0(tdf1_dot_product_U0_ifmap_vec_address0),
    .ifmap_vec_ce0(tdf1_dot_product_U0_ifmap_vec_ce0),
    .ifmap_vec_q0(ifmap_vec_t_q0),
    .weight_vecs_0_address0(tdf1_dot_product_U0_weight_vecs_0_address0),
    .weight_vecs_0_ce0(tdf1_dot_product_U0_weight_vecs_0_ce0),
    .weight_vecs_0_q0(weight_vecs_0_t_q0),
    .products_0_address0(tdf1_dot_product_U0_products_0_address0),
    .products_0_ce0(tdf1_dot_product_U0_products_0_ce0),
    .products_0_we0(tdf1_dot_product_U0_products_0_we0),
    .products_0_d0(tdf1_dot_product_U0_products_0_d0)
);

td_fused_top_tdf1_accum_1 tdf1_accum_1_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf1_accum_1_U0_ap_start),
    .ap_done(tdf1_accum_1_U0_ap_done),
    .ap_continue(tdf1_accum_1_U0_ap_continue),
    .ap_idle(tdf1_accum_1_U0_ap_idle),
    .ap_ready(tdf1_accum_1_U0_ap_ready),
    .accum_in_0_address0(tdf1_accum_1_U0_accum_in_0_address0),
    .accum_in_0_ce0(tdf1_accum_1_U0_accum_in_0_ce0),
    .accum_in_0_q0(products_0_t_q0),
    .accum_in_0_address1(tdf1_accum_1_U0_accum_in_0_address1),
    .accum_in_0_ce1(tdf1_accum_1_U0_accum_in_0_ce1),
    .accum_in_0_q1(products_0_t_q1),
    .accum_out_address0(tdf1_accum_1_U0_accum_out_address0),
    .accum_out_ce0(tdf1_accum_1_U0_accum_out_ce0),
    .accum_out_we0(tdf1_accum_1_U0_accum_out_we0),
    .accum_out_d0(tdf1_accum_1_U0_accum_out_d0)
);

td_fused_top_tdf1_accum_2 tdf1_accum_2_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf1_accum_2_U0_ap_start),
    .ap_done(tdf1_accum_2_U0_ap_done),
    .ap_continue(tdf1_accum_2_U0_ap_continue),
    .ap_idle(tdf1_accum_2_U0_ap_idle),
    .ap_ready(tdf1_accum_2_U0_ap_ready),
    .accum_in_address0(tdf1_accum_2_U0_accum_in_address0),
    .accum_in_ce0(tdf1_accum_2_U0_accum_in_ce0),
    .accum_in_q0(accum1_out_0_t_q0),
    .accum_in_address1(tdf1_accum_2_U0_accum_in_address1),
    .accum_in_ce1(tdf1_accum_2_U0_accum_in_ce1),
    .accum_in_q1(accum1_out_0_t_q1),
    .accum_out_address0(tdf1_accum_2_U0_accum_out_address0),
    .accum_out_ce0(tdf1_accum_2_U0_accum_out_ce0),
    .accum_out_we0(tdf1_accum_2_U0_accum_out_we0),
    .accum_out_d0(tdf1_accum_2_U0_accum_out_d0)
);

td_fused_top_tdf1_accum_3 tdf1_accum_3_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf1_accum_3_U0_ap_start),
    .ap_done(tdf1_accum_3_U0_ap_done),
    .ap_continue(tdf1_accum_3_U0_ap_continue),
    .ap_idle(tdf1_accum_3_U0_ap_idle),
    .ap_ready(tdf1_accum_3_U0_ap_ready),
    .accum_in_18(tdf1_accum_3_U0_accum_in_18),
    .accum_in_18_ap_vld(tdf1_accum_3_U0_accum_in_18_ap_vld),
    .accum_in_address0(tdf1_accum_3_U0_accum_in_address0),
    .accum_in_ce0(tdf1_accum_3_U0_accum_in_ce0),
    .accum_in_q0(accum2_out_0_t_q0)
);

td_fused_top_Block_entry_proc_proc Block_entry_proc_proc_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(Block_entry_proc_proc_U0_ap_start),
    .ap_done(Block_entry_proc_proc_U0_ap_done),
    .ap_continue(Block_entry_proc_proc_U0_ap_continue),
    .ap_idle(Block_entry_proc_proc_U0_ap_idle),
    .ap_ready(Block_entry_proc_proc_U0_ap_ready),
    .tmp(tmp_channel_dout),
    .ap_return(Block_entry_proc_proc_U0_ap_return)
);

td_fused_top_tdf1_adjust tdf1_adjust_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf1_adjust_U0_ap_start),
    .ap_done(tdf1_adjust_U0_ap_done),
    .ap_continue(tdf1_adjust_U0_ap_continue),
    .ap_idle(tdf1_adjust_U0_ap_idle),
    .ap_ready(tdf1_adjust_U0_ap_ready),
    .sums_read(sums_0_dout),
    .adjustments_address0(tdf1_adjust_U0_adjustments_address0),
    .adjustments_ce0(tdf1_adjust_U0_adjustments_ce0),
    .adjustments_q0(adjustments_q0),
    .input_indices_23_dout(input_indices_23_c1_dout),
    .input_indices_23_empty_n(input_indices_23_c1_empty_n),
    .input_indices_23_read(tdf1_adjust_U0_input_indices_23_read),
    .ap_return(tdf1_adjust_U0_ap_return)
);

td_fused_top_tdf1_poolOutputs tdf1_poolOutputs_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf1_poolOutputs_U0_ap_start),
    .ap_done(tdf1_poolOutputs_U0_ap_done),
    .ap_continue(tdf1_poolOutputs_U0_ap_continue),
    .ap_idle(tdf1_poolOutputs_U0_ap_idle),
    .ap_ready(tdf1_poolOutputs_U0_ap_ready),
    .output_indices_04_dout(output_indices_04_c_dout),
    .output_indices_04_empty_n(output_indices_04_c_empty_n),
    .output_indices_04_read(tdf1_poolOutputs_U0_output_indices_04_read),
    .output_indices_15_dout(output_indices_15_c_dout),
    .output_indices_15_empty_n(output_indices_15_c_empty_n),
    .output_indices_15_read(tdf1_poolOutputs_U0_output_indices_15_read),
    .resetMaximum6_dout(resetMaximum6_c_dout),
    .resetMaximum6_empty_n(resetMaximum6_c_empty_n),
    .resetMaximum6_read(tdf1_poolOutputs_U0_resetMaximum6_read),
    .storeOutput7_dout(storeOutput7_c_dout),
    .storeOutput7_empty_n(storeOutput7_c_empty_n),
    .storeOutput7_read(tdf1_poolOutputs_U0_storeOutput7_read),
    .p_read(outputs_0_dout),
    .out_data_address1(tdf1_poolOutputs_U0_out_data_address1),
    .out_data_ce1(tdf1_poolOutputs_U0_out_data_ce1),
    .out_data_we1(tdf1_poolOutputs_U0_out_data_we1),
    .out_data_d1(tdf1_poolOutputs_U0_out_data_d1)
);

td_fused_top_fifo_w4_d2_S input_indices_23_c_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(input_indices_23_c_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf1_readFilters18_U0_input_indices_23_read),
    .if_dout(input_indices_23_c_dout),
    .if_full_n(input_indices_23_c_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf1_get_next_ijk_U0_input_indices_2_out_write),
    .if_din(tdf1_get_next_ijk_U0_input_indices_2_out_din)
);

td_fused_top_fifo_w4_d8_S input_indices_23_c1_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(input_indices_23_c1_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf1_adjust_U0_input_indices_23_read),
    .if_dout(input_indices_23_c1_dout),
    .if_full_n(input_indices_23_c1_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf1_get_next_ijk_U0_input_indices_2_out1_write),
    .if_din(tdf1_get_next_ijk_U0_input_indices_2_out1_din)
);

td_fused_top_fifo_w7_d9_S output_indices_04_c_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(output_indices_04_c_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf1_poolOutputs_U0_output_indices_04_read),
    .if_dout(output_indices_04_c_dout),
    .if_full_n(output_indices_04_c_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf1_get_next_ijk_U0_output_indices_0_write),
    .if_din(tdf1_get_next_ijk_U0_output_indices_0_din)
);

td_fused_top_fifo_w14_d9_S output_indices_15_c_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(output_indices_15_c_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf1_poolOutputs_U0_output_indices_15_read),
    .if_dout(output_indices_15_c_dout),
    .if_full_n(output_indices_15_c_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf1_get_next_ijk_U0_output_indices_1_write),
    .if_din(tdf1_get_next_ijk_U0_output_indices_1_din)
);

td_fused_top_fifo_w1_d9_S resetMaximum6_c_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(resetMaximum6_c_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf1_poolOutputs_U0_resetMaximum6_read),
    .if_dout(resetMaximum6_c_dout),
    .if_full_n(resetMaximum6_c_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf1_get_next_ijk_U0_resetMaximum_write),
    .if_din(resetMaximum6_c_din)
);

td_fused_top_fifo_w1_d9_S storeOutput7_c_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(storeOutput7_c_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf1_poolOutputs_U0_storeOutput7_read),
    .if_dout(storeOutput7_c_dout),
    .if_full_n(storeOutput7_c_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf1_get_next_ijk_U0_storeOutput_write),
    .if_din(storeOutput7_c_din)
);

td_fused_top_fifo_w16_d2_S input_indices_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(input_indices_0_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf1_readInputs19_U0_ap_ready),
    .if_dout(input_indices_0_dout),
    .if_full_n(input_indices_0_full_n),
    .if_write_ce(1'b1),
    .if_write(ap_channel_done_input_indices_0),
    .if_din(tdf1_get_next_ijk_U0_ap_return_0)
);

td_fused_top_fifo_w16_d2_S input_indices_1_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(input_indices_1_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf1_readInputs19_U0_ap_ready),
    .if_dout(input_indices_1_dout),
    .if_full_n(input_indices_1_full_n),
    .if_write_ce(1'b1),
    .if_write(ap_channel_done_input_indices_1),
    .if_din(tdf1_get_next_ijk_U0_ap_return_1)
);

td_fused_top_fifo_w16_d2_S tmp_channel_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(tmp_channel_empty_n),
    .if_read_ce(1'b1),
    .if_read(Block_entry_proc_proc_U0_ap_ready),
    .if_dout(tmp_channel_dout),
    .if_full_n(tmp_channel_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf1_accum_3_U0_ap_done),
    .if_din(tdf1_accum_3_U0_accum_in_18)
);

td_fused_top_fifo_w16_d2_S sums_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(sums_0_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf1_adjust_U0_ap_ready),
    .if_dout(sums_0_dout),
    .if_full_n(sums_0_full_n),
    .if_write_ce(1'b1),
    .if_write(Block_entry_proc_proc_U0_ap_done),
    .if_din(Block_entry_proc_proc_U0_ap_return)
);

td_fused_top_fifo_w16_d2_S outputs_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(outputs_0_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf1_poolOutputs_U0_ap_ready),
    .if_dout(outputs_0_dout),
    .if_full_n(outputs_0_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf1_adjust_U0_ap_done),
    .if_din(tdf1_adjust_U0_ap_return)
);

td_fused_top_start_for_tdf1_readFilters18_U0 start_for_tdf1_readFilters18_U0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(start_for_tdf1_readFilters18_U0_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf1_readFilters18_U0_ap_ready),
    .if_dout(start_for_tdf1_readFilters18_U0_dout),
    .if_full_n(start_for_tdf1_readFilters18_U0_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf1_get_next_ijk_U0_start_write),
    .if_din(start_for_tdf1_readFilters18_U0_din)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_sync_reg_channel_write_input_indices_0 <= 1'b0;
    end else begin
        if (((tdf1_get_next_ijk_U0_ap_done & tdf1_get_next_ijk_U0_ap_continue) == 1'b1)) begin
            ap_sync_reg_channel_write_input_indices_0 <= 1'b0;
        end else begin
            ap_sync_reg_channel_write_input_indices_0 <= ap_sync_channel_write_input_indices_0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_sync_reg_channel_write_input_indices_1 <= 1'b0;
    end else begin
        if (((tdf1_get_next_ijk_U0_ap_done & tdf1_get_next_ijk_U0_ap_continue) == 1'b1)) begin
            ap_sync_reg_channel_write_input_indices_1 <= 1'b0;
        end else begin
            ap_sync_reg_channel_write_input_indices_1 <= ap_sync_channel_write_input_indices_1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_sync_reg_tdf1_get_next_ijk_U0_ap_ready <= 1'b0;
    end else begin
        if (((ap_sync_ready & ap_start) == 1'b1)) begin
            ap_sync_reg_tdf1_get_next_ijk_U0_ap_ready <= 1'b0;
        end else begin
            ap_sync_reg_tdf1_get_next_ijk_U0_ap_ready <= ap_sync_tdf1_get_next_ijk_U0_ap_ready;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_sync_reg_tdf1_readInputs19_U0_ap_ready <= 1'b0;
    end else begin
        if (((ap_sync_ready & ap_start) == 1'b1)) begin
            ap_sync_reg_tdf1_readInputs19_U0_ap_ready <= 1'b0;
        end else begin
            ap_sync_reg_tdf1_readInputs19_U0_ap_ready <= ap_sync_tdf1_readInputs19_U0_ap_ready;
        end
    end
end

assign Block_entry_proc_proc_U0_ap_continue = sums_0_full_n;

assign Block_entry_proc_proc_U0_ap_start = tmp_channel_empty_n;

assign Block_entry_proc_proc_U0_start_full_n = 1'b1;

assign Block_entry_proc_proc_U0_start_write = 1'b0;

assign accum1_out_0_t_d1 = 16'd0;

assign accum1_out_0_t_we1 = 1'b0;

assign adjustments_address0 = tdf1_adjust_U0_adjustments_address0;

assign adjustments_address1 = 4'd0;

assign adjustments_ce0 = tdf1_adjust_U0_adjustments_ce0;

assign adjustments_ce1 = 1'b0;

assign adjustments_d0 = 48'd0;

assign adjustments_d1 = 48'd0;

assign adjustments_we0 = 1'b0;

assign adjustments_we1 = 1'b0;

assign ap_channel_done_accum1_out_0 = tdf1_accum_1_U0_ap_done;

assign ap_channel_done_accum2_out_0 = tdf1_accum_2_U0_ap_done;

assign ap_channel_done_ifmap_vec = tdf1_readInputs19_U0_ap_done;

assign ap_channel_done_input_indices_0 = (tdf1_get_next_ijk_U0_ap_done & (ap_sync_reg_channel_write_input_indices_0 ^ 1'b1));

assign ap_channel_done_input_indices_1 = (tdf1_get_next_ijk_U0_ap_done & (ap_sync_reg_channel_write_input_indices_1 ^ 1'b1));

assign ap_channel_done_outputs_0 = tdf1_adjust_U0_ap_done;

assign ap_channel_done_products_0 = tdf1_dot_product_U0_ap_done;

assign ap_channel_done_sums_0 = Block_entry_proc_proc_U0_ap_done;

assign ap_channel_done_tmp_channel = tdf1_accum_3_U0_ap_done;

assign ap_channel_done_weight_vecs_0 = tdf1_readFilters18_U0_ap_done;

assign ap_done = tdf1_poolOutputs_U0_ap_done;

assign ap_idle = (tdf1_readInputs19_U0_ap_idle & tdf1_readFilters18_U0_ap_idle & tdf1_poolOutputs_U0_ap_idle & tdf1_get_next_ijk_U0_ap_idle & tdf1_dot_product_U0_ap_idle & tdf1_adjust_U0_ap_idle & tdf1_accum_3_U0_ap_idle & tdf1_accum_2_U0_ap_idle & tdf1_accum_1_U0_ap_idle & (outputs_0_empty_n ^ 1'b1) & (sums_0_empty_n ^ 1'b1) & (tmp_channel_empty_n ^ 1'b1) & (input_indices_1_empty_n ^ 1'b1) & (input_indices_0_empty_n ^ 1'b1) & (products_0_t_empty_n ^ 1'b1) & (weight_vecs_0_t_empty_n ^ 1'b1) & (ifmap_vec_t_empty_n ^ 1'b1) & (1'b1 ^ accum2_out_0_t_empty_n) & (1'b1 ^ accum1_out_0_t_empty_n) & Block_entry_proc_proc_U0_ap_idle);

assign ap_ready = ap_sync_ready;

assign ap_sync_channel_write_input_indices_0 = ((input_indices_0_full_n & ap_channel_done_input_indices_0) | ap_sync_reg_channel_write_input_indices_0);

assign ap_sync_channel_write_input_indices_1 = ((input_indices_1_full_n & ap_channel_done_input_indices_1) | ap_sync_reg_channel_write_input_indices_1);

assign ap_sync_continue = ap_continue;

assign ap_sync_done = tdf1_poolOutputs_U0_ap_done;

assign ap_sync_ready = (ap_sync_tdf1_readInputs19_U0_ap_ready & ap_sync_tdf1_get_next_ijk_U0_ap_ready);

assign ap_sync_tdf1_get_next_ijk_U0_ap_ready = (tdf1_get_next_ijk_U0_ap_ready | ap_sync_reg_tdf1_get_next_ijk_U0_ap_ready);

assign ap_sync_tdf1_readInputs19_U0_ap_ready = (tdf1_readInputs19_U0_ap_ready | ap_sync_reg_tdf1_readInputs19_U0_ap_ready);

assign filter_data_address0 = tdf1_readFilters18_U0_filter_data_address0;

assign filter_data_address1 = 9'd0;

assign filter_data_ce0 = tdf1_readFilters18_U0_filter_data_ce0;

assign filter_data_ce1 = 1'b0;

assign filter_data_d0 = 16'd0;

assign filter_data_d1 = 16'd0;

assign filter_data_we0 = 1'b0;

assign filter_data_we1 = 1'b0;

assign in_data_address0 = tdf1_readInputs19_U0_in_data_address0;

assign in_data_address1 = 16'd0;

assign in_data_ce0 = tdf1_readInputs19_U0_in_data_ce0;

assign in_data_ce1 = 1'b0;

assign in_data_d0 = 64'd0;

assign in_data_d1 = 64'd0;

assign in_data_read = tdf1_readInputs19_U0_in_data_write;

assign in_data_we0 = 1'b0;

assign in_data_we1 = 1'b0;

assign out_data_address0 = 16'd0;

assign out_data_address1 = tdf1_poolOutputs_U0_out_data_address1;

assign out_data_ce0 = 1'b0;

assign out_data_ce1 = tdf1_poolOutputs_U0_out_data_ce1;

assign out_data_d0 = 64'd0;

assign out_data_d1 = tdf1_poolOutputs_U0_out_data_d1;

assign out_data_we0 = 1'b0;

assign out_data_we1 = tdf1_poolOutputs_U0_out_data_we1;

assign out_data_write = tdf1_poolOutputs_U0_out_data_write;

assign products_0_t_d1 = 16'd0;

assign products_0_t_we1 = 1'b0;

assign resetMaximum6_c_din = tdf1_get_next_ijk_U0_resetMaximum_din;

assign start_for_tdf1_readFilters18_U0_din = 1'b1;

assign storeOutput7_c_din = tdf1_get_next_ijk_U0_storeOutput_din;

assign tdf1_accum_1_U0_accum_out_full_n = accum1_out_0_i_full_n;

assign tdf1_accum_1_U0_ap_continue = accum1_out_0_i_full_n;

assign tdf1_accum_1_U0_ap_start = products_0_t_empty_n;

assign tdf1_accum_1_U0_start_full_n = 1'b1;

assign tdf1_accum_1_U0_start_write = 1'b0;

assign tdf1_accum_2_U0_accum_out_full_n = accum2_out_0_i_full_n;

assign tdf1_accum_2_U0_ap_continue = accum2_out_0_i_full_n;

assign tdf1_accum_2_U0_ap_start = accum1_out_0_t_empty_n;

assign tdf1_accum_2_U0_start_full_n = 1'b1;

assign tdf1_accum_2_U0_start_write = 1'b0;

assign tdf1_accum_3_U0_ap_continue = tmp_channel_full_n;

assign tdf1_accum_3_U0_ap_start = accum2_out_0_t_empty_n;

assign tdf1_accum_3_U0_start_full_n = 1'b1;

assign tdf1_accum_3_U0_start_write = 1'b0;

assign tdf1_adjust_U0_ap_continue = outputs_0_full_n;

assign tdf1_adjust_U0_ap_start = sums_0_empty_n;

assign tdf1_adjust_U0_start_full_n = 1'b1;

assign tdf1_adjust_U0_start_write = 1'b0;

assign tdf1_dot_product_U0_ap_continue = products_0_i_full_n;

assign tdf1_dot_product_U0_ap_start = (weight_vecs_0_t_empty_n & ifmap_vec_t_empty_n);

assign tdf1_dot_product_U0_products_0_full_n = products_0_i_full_n;

assign tdf1_dot_product_U0_start_full_n = 1'b1;

assign tdf1_dot_product_U0_start_write = 1'b0;

assign tdf1_get_next_ijk_U0_ap_continue = (ap_sync_channel_write_input_indices_1 & ap_sync_channel_write_input_indices_0);

assign tdf1_get_next_ijk_U0_ap_start = ((ap_sync_reg_tdf1_get_next_ijk_U0_ap_ready ^ 1'b1) & ap_start);

assign tdf1_poolOutputs_U0_ap_continue = ap_continue;

assign tdf1_poolOutputs_U0_ap_start = outputs_0_empty_n;

assign tdf1_poolOutputs_U0_out_data_full_n = out_data_full_n;

assign tdf1_poolOutputs_U0_out_data_write = 1'b0;

assign tdf1_poolOutputs_U0_start_full_n = 1'b1;

assign tdf1_poolOutputs_U0_start_write = 1'b0;

assign tdf1_readFilters18_U0_ap_continue = weight_vecs_0_i_full_n;

assign tdf1_readFilters18_U0_ap_start = start_for_tdf1_readFilters18_U0_empty_n;

assign tdf1_readFilters18_U0_start_full_n = 1'b1;

assign tdf1_readFilters18_U0_start_write = 1'b0;

assign tdf1_readFilters18_U0_weight_vecs_0_full_n = weight_vecs_0_i_full_n;

assign tdf1_readInputs19_U0_ap_continue = ifmap_vec_i_full_n;

assign tdf1_readInputs19_U0_ap_start = (input_indices_1_empty_n & input_indices_0_empty_n & (ap_sync_reg_tdf1_readInputs19_U0_ap_ready ^ 1'b1) & ap_start);

assign tdf1_readInputs19_U0_ifmap_vec_full_n = ifmap_vec_i_full_n;

assign tdf1_readInputs19_U0_in_data_full_n = in_data_empty_n;

assign tdf1_readInputs19_U0_in_data_write = 1'b0;

assign tdf1_readInputs19_U0_start_full_n = 1'b1;

assign tdf1_readInputs19_U0_start_write = 1'b0;

endmodule //td_fused_top_dataflow_in_loop_TOP_LOOP38116
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP38270_accum1_out_0_memcore_ram (addr0, ce0, d0, we0, q0, addr1, ce1, d1, we1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 3;
parameter MEM_SIZE = 8;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
input clk;

reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];




always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1) 
            ram[addr1] <= d1; 
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP38270_accum1_out_0_memcore(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    q0,
    address1,
    ce1,
    we1,
    d1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd8;
parameter AddressWidth = 32'd3;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;



td_fused_top_dataflow_in_loop_TOP_LOOP38270_accum1_out_0_memcore_ram td_fused_top_dataflow_in_loop_TOP_LOOP38270_accum1_out_0_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_dataflow_in_loop_TOP_LOOP38270_accum1_out_0
#(parameter
    DataWidth    = 16,
    AddressRange = 32,
    AddressWidth = 3,
    BufferCount  = 2,
    MemLatency   = 1,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire                    i_we0,
    input  wire [AddressWidth-1:0] i_address0,
    input  wire [DataWidth-1:0]    i_d0,
    output wire [DataWidth-1:0]    i_q0,
    input  wire                    i_ce1,
    input  wire                    i_we1,
    input  wire [AddressWidth-1:0] i_address1,
    input  wire [DataWidth-1:0]    i_d1,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire                    t_we0,
    input  wire [AddressWidth-1:0] t_address0,
    input  wire [DataWidth-1:0]    t_d0,
    output wire [DataWidth-1:0]    t_q0,
    input  wire                    t_ce1,
    input  wire                    t_we1,
    input  wire [AddressWidth-1:0] t_address1,
    input  wire [DataWidth-1:0]    t_d1
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth-1:0]   prev_iptr    = 1'b0; // previous initiator index
reg  [IndexWidth-1:0]   prev_tptr    = 1'b0; // previous target index
reg  [DataWidth-1:0]    reg_q0      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid0    = 1'b0; // buffer has valid data
reg  [DataWidth-1:0]    reg_q1      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid1    = 1'b0; // buffer has valid data
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
// buffer signals
wire [BufferCount-1:0] buf_ce0;
wire [BufferCount-1:0] buf_we0;
wire [AddressWidth-1:0] buf_a0_0, buf_a0_1;
wire [DataWidth-1:0] buf_d0_0, buf_d0_1;
wire [DataWidth-1:0] buf_q0_0, buf_q0_1;
wire [BufferCount-1:0] buf_ce1;
wire [BufferCount-1:0] buf_we1;
wire [AddressWidth-1:0] buf_a1_0, buf_a1_1;
wire [DataWidth-1:0] buf_d1_0, buf_d1_1;
//------------------------Instantiation------------------
//genvar i;
        td_fused_top_dataflow_in_loop_TOP_LOOP38270_accum1_out_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP38270_accum1_out_0_memcore_U_0 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_0 ),
            .ce0      ( buf_ce0[ 0 ] ),
            .we0      ( buf_we0[ 0 ] ),
            .d0       ( buf_d0_0 ),
            .q0       ( buf_q0_0 ),
            .address1 ( buf_a1_0 ),
            .ce1      ( buf_ce1[ 0 ] ),
            .we1      ( buf_we1[ 0 ] ),
            .d1       ( buf_d1_0 )
        );
        td_fused_top_dataflow_in_loop_TOP_LOOP38270_accum1_out_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP38270_accum1_out_0_memcore_U_1 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_1 ),
            .ce0      ( buf_ce0[ 1 ] ),
            .we0      ( buf_we0[ 1 ] ),
            .d0       ( buf_d0_1 ),
            .q0       ( buf_q0_1 ),
            .address1 ( buf_a1_1 ),
            .ce1      ( buf_ce1[ 1 ] ),
            .we1      ( buf_we1[ 1 ] ),
            .d1       ( buf_d1_1 )
        );

//++++++++++++++++++++++++buffer signals+++++++++++++++++
        assign buf_ce0[ 0 ] = (tptr ==  0  && empty_n) ? t_ce0
                             : (iptr ==  0 ) ? i_ce0 : 1'b0;
        assign buf_a0_0  = (tptr ==  0  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 0 ] = (tptr ==  0  && empty_n)  ? t_we0
                             : (iptr ==  0 ) ? i_we0 : 1'b0;
        assign buf_d0_0  = (tptr ==  0  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 0 ] = (tptr ==  0  && empty_n) ? t_ce1
                             : (iptr ==  0 ) ? i_ce1 : 1'b0;
        assign buf_a1_0  = (tptr ==  0  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 0 ] = (tptr ==  0  && empty_n)  ? t_we1
                             : (iptr ==  0 ) ? i_we1 : 1'b0;
        assign buf_d1_0  = (tptr ==  0  && empty_n) ? t_d1       : i_d1;
        assign buf_ce0[ 1 ] = (tptr ==  1  && empty_n) ? t_ce0
                             : (iptr ==  1 ) ? i_ce0 : 1'b0;
        assign buf_a0_1  = (tptr ==  1  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 1 ] = (tptr ==  1  && empty_n)  ? t_we0
                             : (iptr ==  1 ) ? i_we0 : 1'b0;
        assign buf_d0_1  = (tptr ==  1  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 1 ] = (tptr ==  1  && empty_n) ? t_ce1
                             : (iptr ==  1 ) ? i_ce1 : 1'b0;
        assign buf_a1_1  = (tptr ==  1  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 1 ] = (tptr ==  1  && empty_n)  ? t_we1
                             : (iptr ==  1 ) ? i_we1 : 1'b0;
        assign buf_d1_1  = (tptr ==  1  && empty_n) ? t_d1       : i_d1;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//------------------------Body---------------------------
assign i_q0      = (prev_iptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign t_q0      = reg_valid0 ? reg_q0 : (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// prev_iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_iptr <= 1'b0;
    else begin
        prev_iptr <= iptr;
    end
end

// prev_tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_tptr <= 1'b0;
    else begin
        prev_tptr <= tptr;
    end
end

// reg_q0 and reg_valid0
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q0     <= 1'b0;
        reg_valid0 <= 1'b0;
    end else if (!t_ce0 && !reg_valid0) begin
        reg_q0     <= (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
        reg_valid0 <= 1'b1;
    end else if (t_ce0) begin
        reg_valid0 <= 1'b0;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP38270_ifmap_vec_memcore_ram (addr0, ce0, d0, we0, q0, addr1, ce1, d1, we1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 10;
parameter MEM_SIZE = 576;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
input clk;

reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];




always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1) 
            ram[addr1] <= d1; 
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP38270_ifmap_vec_memcore(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    q0,
    address1,
    ce1,
    we1,
    d1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd576;
parameter AddressWidth = 32'd10;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;



td_fused_top_dataflow_in_loop_TOP_LOOP38270_ifmap_vec_memcore_ram td_fused_top_dataflow_in_loop_TOP_LOOP38270_ifmap_vec_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_dataflow_in_loop_TOP_LOOP38270_ifmap_vec
#(parameter
    DataWidth    = 16,
    AddressRange = 32,
    AddressWidth = 10,
    BufferCount  = 2,
    MemLatency   = 1,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire                    i_we0,
    input  wire [AddressWidth-1:0] i_address0,
    input  wire [DataWidth-1:0]    i_d0,
    output wire [DataWidth-1:0]    i_q0,
    input  wire                    i_ce1,
    input  wire                    i_we1,
    input  wire [AddressWidth-1:0] i_address1,
    input  wire [DataWidth-1:0]    i_d1,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire                    t_we0,
    input  wire [AddressWidth-1:0] t_address0,
    input  wire [DataWidth-1:0]    t_d0,
    output wire [DataWidth-1:0]    t_q0,
    input  wire                    t_ce1,
    input  wire                    t_we1,
    input  wire [AddressWidth-1:0] t_address1,
    input  wire [DataWidth-1:0]    t_d1
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth-1:0]   prev_iptr    = 1'b0; // previous initiator index
reg  [IndexWidth-1:0]   prev_tptr    = 1'b0; // previous target index
reg  [DataWidth-1:0]    reg_q0      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid0    = 1'b0; // buffer has valid data
reg  [DataWidth-1:0]    reg_q1      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid1    = 1'b0; // buffer has valid data
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
// buffer signals
wire [BufferCount-1:0] buf_ce0;
wire [BufferCount-1:0] buf_we0;
wire [AddressWidth-1:0] buf_a0_0, buf_a0_1;
wire [DataWidth-1:0] buf_d0_0, buf_d0_1;
wire [DataWidth-1:0] buf_q0_0, buf_q0_1;
wire [BufferCount-1:0] buf_ce1;
wire [BufferCount-1:0] buf_we1;
wire [AddressWidth-1:0] buf_a1_0, buf_a1_1;
wire [DataWidth-1:0] buf_d1_0, buf_d1_1;
//------------------------Instantiation------------------
//genvar i;
        td_fused_top_dataflow_in_loop_TOP_LOOP38270_ifmap_vec_memcore td_fused_top_dataflow_in_loop_TOP_LOOP38270_ifmap_vec_memcore_U_0 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_0 ),
            .ce0      ( buf_ce0[ 0 ] ),
            .we0      ( buf_we0[ 0 ] ),
            .d0       ( buf_d0_0 ),
            .q0       ( buf_q0_0 ),
            .address1 ( buf_a1_0 ),
            .ce1      ( buf_ce1[ 0 ] ),
            .we1      ( buf_we1[ 0 ] ),
            .d1       ( buf_d1_0 )
        );
        td_fused_top_dataflow_in_loop_TOP_LOOP38270_ifmap_vec_memcore td_fused_top_dataflow_in_loop_TOP_LOOP38270_ifmap_vec_memcore_U_1 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_1 ),
            .ce0      ( buf_ce0[ 1 ] ),
            .we0      ( buf_we0[ 1 ] ),
            .d0       ( buf_d0_1 ),
            .q0       ( buf_q0_1 ),
            .address1 ( buf_a1_1 ),
            .ce1      ( buf_ce1[ 1 ] ),
            .we1      ( buf_we1[ 1 ] ),
            .d1       ( buf_d1_1 )
        );

//++++++++++++++++++++++++buffer signals+++++++++++++++++
        assign buf_ce0[ 0 ] = (tptr ==  0  && empty_n) ? t_ce0
                             : (iptr ==  0 ) ? i_ce0 : 1'b0;
        assign buf_a0_0  = (tptr ==  0  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 0 ] = (tptr ==  0  && empty_n)  ? t_we0
                             : (iptr ==  0 ) ? i_we0 : 1'b0;
        assign buf_d0_0  = (tptr ==  0  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 0 ] = (tptr ==  0  && empty_n) ? t_ce1
                             : (iptr ==  0 ) ? i_ce1 : 1'b0;
        assign buf_a1_0  = (tptr ==  0  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 0 ] = (tptr ==  0  && empty_n)  ? t_we1
                             : (iptr ==  0 ) ? i_we1 : 1'b0;
        assign buf_d1_0  = (tptr ==  0  && empty_n) ? t_d1       : i_d1;
        assign buf_ce0[ 1 ] = (tptr ==  1  && empty_n) ? t_ce0
                             : (iptr ==  1 ) ? i_ce0 : 1'b0;
        assign buf_a0_1  = (tptr ==  1  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 1 ] = (tptr ==  1  && empty_n)  ? t_we0
                             : (iptr ==  1 ) ? i_we0 : 1'b0;
        assign buf_d0_1  = (tptr ==  1  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 1 ] = (tptr ==  1  && empty_n) ? t_ce1
                             : (iptr ==  1 ) ? i_ce1 : 1'b0;
        assign buf_a1_1  = (tptr ==  1  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 1 ] = (tptr ==  1  && empty_n)  ? t_we1
                             : (iptr ==  1 ) ? i_we1 : 1'b0;
        assign buf_d1_1  = (tptr ==  1  && empty_n) ? t_d1       : i_d1;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//------------------------Body---------------------------
assign i_q0      = (prev_iptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign t_q0      = reg_valid0 ? reg_q0 : (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// prev_iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_iptr <= 1'b0;
    else begin
        prev_iptr <= iptr;
    end
end

// prev_tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_tptr <= 1'b0;
    else begin
        prev_tptr <= tptr;
    end
end

// reg_q0 and reg_valid0
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q0     <= 1'b0;
        reg_valid0 <= 1'b0;
    end else if (!t_ce0 && !reg_valid0) begin
        reg_q0     <= (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
        reg_valid0 <= 1'b1;
    end else if (t_ce0) begin
        reg_valid0 <= 1'b0;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP38270_l2_products_memcore_ram (addr0, ce0, d0, we0, q0, addr1, ce1, d1, we1, q1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 8;
parameter MEM_SIZE = 256;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
output reg[DWIDTH-1:0] q1;
input clk;

 reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];




always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1) 
            ram[addr1] <= d1; 
        q1 <= ram[addr1];
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP38270_l2_products_memcore(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    q0,
    address1,
    ce1,
    we1,
    d1,
    q1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd256;
parameter AddressWidth = 32'd8;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;
output[DataWidth - 1:0] q1;



td_fused_top_dataflow_in_loop_TOP_LOOP38270_l2_products_memcore_ram td_fused_top_dataflow_in_loop_TOP_LOOP38270_l2_products_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 ),
    .q1( q1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_dataflow_in_loop_TOP_LOOP38270_l2_products
#(parameter
    DataWidth    = 16,
    AddressRange = 32,
    AddressWidth = 7,
    BufferCount  = 2,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire                    i_we0,
    input  wire [AddressWidth-1:0] i_address0,
    input  wire [DataWidth-1:0]    i_d0,
    output wire [DataWidth-1:0]    i_q0,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire                    t_we0,
    input  wire [AddressWidth-1:0] t_address0,
    input  wire [DataWidth-1:0]    t_d0,
    output wire [DataWidth-1:0]    t_q0
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
wire [AddressWidth+IndexWidth-1:0]   memcore_iaddr;
wire [AddressWidth+IndexWidth-1:0]   memcore_taddr;

//------------------------Instantiation------------------
assign memcore_iaddr = {i_address0, iptr};
assign memcore_taddr = {t_address0, tptr};
td_fused_top_dataflow_in_loop_TOP_LOOP38270_l2_products_memcore td_fused_top_dataflow_in_loop_TOP_LOOP38270_l2_products_memcore_U (
    .reset    ( reset ),
    .clk      ( clk ),
    .address0 ( memcore_iaddr ),
    .ce0      ( i_ce0 ),
    .we0      ( i_we0),
    .d0       ( i_d0 ),
    .q0       ( i_q0 ),
    .address1 ( memcore_taddr ),
    .ce1      ( t_ce0 ),
    .we1      ( t_we0),
    .d1       ( t_d0 ),
    .q1       ( t_q0 )

);

//------------------------Body---------------------------

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP38270_products_0_memcore_ram (addr0, ce0, d0, we0, q0, addr1, ce1, q1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 10;
parameter MEM_SIZE = 576;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
output reg[DWIDTH-1:0] q1;
input clk;

reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];




always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        q1 <= ram[addr1];
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP38270_products_0_memcore(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    q0,
    address1,
    ce1,
    q1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd576;
parameter AddressWidth = 32'd10;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
output[DataWidth - 1:0] q1;



td_fused_top_dataflow_in_loop_TOP_LOOP38270_products_0_memcore_ram td_fused_top_dataflow_in_loop_TOP_LOOP38270_products_0_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .q1( q1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_dataflow_in_loop_TOP_LOOP38270_products_0
#(parameter
    DataWidth    = 16,
    AddressRange = 32,
    AddressWidth = 10,
    BufferCount  = 2,
    MemLatency   = 1,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire                    i_we0,
    input  wire [AddressWidth-1:0] i_address0,
    input  wire [DataWidth-1:0]    i_d0,
    output wire [DataWidth-1:0]    i_q0,
    input  wire                    i_ce1,
    input  wire [AddressWidth-1:0] i_address1,
    output wire [DataWidth-1:0]    i_q1,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire                    t_we0,
    input  wire [AddressWidth-1:0] t_address0,
    input  wire [DataWidth-1:0]    t_d0,
    output wire [DataWidth-1:0]    t_q0,
    input  wire                    t_ce1,
    input  wire [AddressWidth-1:0] t_address1,
    output wire [DataWidth-1:0]    t_q1
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth-1:0]   prev_iptr    = 1'b0; // previous initiator index
reg  [IndexWidth-1:0]   prev_tptr    = 1'b0; // previous target index
reg  [DataWidth-1:0]    reg_q0      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid0    = 1'b0; // buffer has valid data
reg  [DataWidth-1:0]    reg_q1      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid1    = 1'b0; // buffer has valid data
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
// buffer signals
wire [BufferCount-1:0] buf_ce0;
wire [BufferCount-1:0] buf_we0;
wire [AddressWidth-1:0] buf_a0_0, buf_a0_1;
wire [DataWidth-1:0] buf_d0_0, buf_d0_1;
wire [DataWidth-1:0] buf_q0_0, buf_q0_1;
wire [BufferCount-1:0] buf_ce1;
wire [AddressWidth-1:0] buf_a1_0, buf_a1_1;
wire [DataWidth-1:0] buf_q1_0, buf_q1_1;
//------------------------Instantiation------------------
//genvar i;
        td_fused_top_dataflow_in_loop_TOP_LOOP38270_products_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP38270_products_0_memcore_U_0 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_0 ),
            .ce0      ( buf_ce0[ 0 ] ),
            .we0      ( buf_we0[ 0 ] ),
            .d0       ( buf_d0_0 ),
            .q0       ( buf_q0_0 ),
            .address1 ( buf_a1_0 ),
            .ce1      ( buf_ce1[ 0 ] ),
            .q1       ( buf_q1_0 )
        );
        td_fused_top_dataflow_in_loop_TOP_LOOP38270_products_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP38270_products_0_memcore_U_1 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_1 ),
            .ce0      ( buf_ce0[ 1 ] ),
            .we0      ( buf_we0[ 1 ] ),
            .d0       ( buf_d0_1 ),
            .q0       ( buf_q0_1 ),
            .address1 ( buf_a1_1 ),
            .ce1      ( buf_ce1[ 1 ] ),
            .q1       ( buf_q1_1 )
        );

//++++++++++++++++++++++++buffer signals+++++++++++++++++
        assign buf_ce0[ 0 ] = (tptr ==  0  && empty_n) ? t_ce0
                             : (iptr ==  0 ) ? i_ce0 : 1'b0;
        assign buf_a0_0  = (tptr ==  0  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 0 ] = (tptr ==  0  && empty_n)  ? t_we0
                             : (iptr ==  0 ) ? i_we0 : 1'b0;
        assign buf_d0_0  = (tptr ==  0  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 0 ] = (tptr ==  0  && empty_n) ? t_ce1
                             : (iptr ==  0 ) ? i_ce1 : 1'b0;
        assign buf_a1_0  = (tptr ==  0  && empty_n) ?  t_address1 : i_address1;
        assign buf_ce0[ 1 ] = (tptr ==  1  && empty_n) ? t_ce0
                             : (iptr ==  1 ) ? i_ce0 : 1'b0;
        assign buf_a0_1  = (tptr ==  1  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 1 ] = (tptr ==  1  && empty_n)  ? t_we0
                             : (iptr ==  1 ) ? i_we0 : 1'b0;
        assign buf_d0_1  = (tptr ==  1  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 1 ] = (tptr ==  1  && empty_n) ? t_ce1
                             : (iptr ==  1 ) ? i_ce1 : 1'b0;
        assign buf_a1_1  = (tptr ==  1  && empty_n) ?  t_address1 : i_address1;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//------------------------Body---------------------------
assign i_q0      = (prev_iptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign t_q0      = reg_valid0 ? reg_q0 : (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign i_q1      = (prev_iptr == 1'b1 ? buf_q1_1 : buf_q1_0);
assign t_q1      = reg_valid1 ? reg_q1 : (prev_tptr == 1'b1 ? buf_q1_1 : buf_q1_0);

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// prev_iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_iptr <= 1'b0;
    else begin
        prev_iptr <= iptr;
    end
end

// prev_tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_tptr <= 1'b0;
    else begin
        prev_tptr <= tptr;
    end
end

// reg_q0 and reg_valid0
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q0     <= 1'b0;
        reg_valid0 <= 1'b0;
    end else if (!t_ce0 && !reg_valid0) begin
        reg_q0     <= (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
        reg_valid0 <= 1'b1;
    end else if (t_ce0) begin
        reg_valid0 <= 1'b0;
    end
end

// reg_q1 and reg_valid1
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q1     <= 1'b0;
        reg_valid1 <= 1'b0;
    end else if (!t_ce1 && !reg_valid1) begin
        reg_q1     <= (prev_tptr == 1'b1 ? buf_q1_1 : buf_q1_0);
        reg_valid1 <= 1'b1;
    end else if (t_ce1) begin
        reg_valid1 <= 1'b0;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_dataflow_in_loop_TOP_LOOP38270 (
        ap_clk,
        ap_rst,
        in_data_address0,
        in_data_ce0,
        in_data_d0,
        in_data_q0,
        in_data_we0,
        in_data_address1,
        in_data_ce1,
        in_data_d1,
        in_data_q1,
        in_data_we1,
        l1_filter_data_address0,
        l1_filter_data_ce0,
        l1_filter_data_d0,
        l1_filter_data_q0,
        l1_filter_data_we0,
        l1_filter_data_address1,
        l1_filter_data_ce1,
        l1_filter_data_d1,
        l1_filter_data_q1,
        l1_filter_data_we1,
        l1_adjustments_address0,
        l1_adjustments_ce0,
        l1_adjustments_d0,
        l1_adjustments_q0,
        l1_adjustments_we0,
        l1_adjustments_address1,
        l1_adjustments_ce1,
        l1_adjustments_d1,
        l1_adjustments_q1,
        l1_adjustments_we1,
        l2_filter_data_address0,
        l2_filter_data_ce0,
        l2_filter_data_d0,
        l2_filter_data_q0,
        l2_filter_data_we0,
        l2_filter_data_address1,
        l2_filter_data_ce1,
        l2_filter_data_d1,
        l2_filter_data_q1,
        l2_filter_data_we1,
        out_data_address0,
        out_data_ce0,
        out_data_d0,
        out_data_q0,
        out_data_we0,
        out_data_address1,
        out_data_ce1,
        out_data_d1,
        out_data_q1,
        out_data_we1,
        l2_adjustments_address0,
        l2_adjustments_ce0,
        l2_adjustments_d0,
        l2_adjustments_q0,
        l2_adjustments_we0,
        l2_adjustments_address1,
        l2_adjustments_ce1,
        l2_adjustments_d1,
        l2_adjustments_q1,
        l2_adjustments_we1,
        ap_start,
        in_data_empty_n,
        in_data_read,
        out_data_full_n,
        out_data_write,
        ap_done,
        ap_ready,
        ap_idle,
        ap_continue
);


input   ap_clk;
input   ap_rst;
output  [11:0] in_data_address0;
output   in_data_ce0;
output  [63:0] in_data_d0;
input  [63:0] in_data_q0;
output   in_data_we0;
output  [11:0] in_data_address1;
output   in_data_ce1;
output  [63:0] in_data_d1;
input  [63:0] in_data_q1;
output   in_data_we1;
output  [16:0] l1_filter_data_address0;
output   l1_filter_data_ce0;
output  [63:0] l1_filter_data_d0;
input  [63:0] l1_filter_data_q0;
output   l1_filter_data_we0;
output  [16:0] l1_filter_data_address1;
output   l1_filter_data_ce1;
output  [63:0] l1_filter_data_d1;
input  [63:0] l1_filter_data_q1;
output   l1_filter_data_we1;
output  [8:0] l1_adjustments_address0;
output   l1_adjustments_ce0;
output  [47:0] l1_adjustments_d0;
input  [47:0] l1_adjustments_q0;
output   l1_adjustments_we0;
output  [8:0] l1_adjustments_address1;
output   l1_adjustments_ce1;
output  [47:0] l1_adjustments_d1;
input  [47:0] l1_adjustments_q1;
output   l1_adjustments_we1;
output  [15:0] l2_filter_data_address0;
output   l2_filter_data_ce0;
output  [15:0] l2_filter_data_d0;
input  [15:0] l2_filter_data_q0;
output   l2_filter_data_we0;
output  [15:0] l2_filter_data_address1;
output   l2_filter_data_ce1;
output  [15:0] l2_filter_data_d1;
input  [15:0] l2_filter_data_q1;
output   l2_filter_data_we1;
output  [12:0] out_data_address0;
output   out_data_ce0;
output  [63:0] out_data_d0;
input  [63:0] out_data_q0;
output   out_data_we0;
output  [12:0] out_data_address1;
output   out_data_ce1;
output  [63:0] out_data_d1;
input  [63:0] out_data_q1;
output   out_data_we1;
output  [6:0] l2_adjustments_address0;
output   l2_adjustments_ce0;
output  [47:0] l2_adjustments_d0;
input  [47:0] l2_adjustments_q0;
output   l2_adjustments_we0;
output  [6:0] l2_adjustments_address1;
output   l2_adjustments_ce1;
output  [47:0] l2_adjustments_d1;
input  [47:0] l2_adjustments_q1;
output   l2_adjustments_we1;
input   ap_start;
input   in_data_empty_n;
output   in_data_read;
input   out_data_full_n;
output   out_data_write;
output   ap_done;
output   ap_ready;
output   ap_idle;
input   ap_continue;

wire   [15:0] ifmap_vec_i_q0;
wire   [15:0] ifmap_vec_t_q0;
wire   [15:0] weight_vecs_0_i_q0;
wire   [15:0] weight_vecs_0_t_q0;
wire   [15:0] products_0_i_q0;
wire   [15:0] products_0_i_q1;
wire   [15:0] products_0_t_q0;
wire   [15:0] products_0_t_q1;
wire   [15:0] accum1_out_0_i_q0;
wire   [15:0] accum1_out_0_t_q0;
wire   [15:0] l2_products_i_q0;
wire   [15:0] l2_products_t_q0;
wire    tdf11_get_next_ijk_U0_ap_start;
wire    tdf11_get_next_ijk_U0_ap_done;
wire    tdf11_get_next_ijk_U0_ap_continue;
wire    tdf11_get_next_ijk_U0_ap_idle;
wire    tdf11_get_next_ijk_U0_ap_ready;
wire    tdf11_get_next_ijk_U0_start_out;
wire    tdf11_get_next_ijk_U0_start_write;
wire   [15:0] tdf11_get_next_ijk_U0_indices_0_din;
wire    tdf11_get_next_ijk_U0_indices_0_write;
wire   [15:0] tdf11_get_next_ijk_U0_indices_1_din;
wire    tdf11_get_next_ijk_U0_indices_1_write;
wire   [8:0] tdf11_get_next_ijk_U0_indices_2_out_din;
wire    tdf11_get_next_ijk_U0_indices_2_out_write;
wire   [8:0] tdf11_get_next_ijk_U0_indices_2_out1_din;
wire    tdf11_get_next_ijk_U0_indices_2_out1_write;
wire    tdf11_get_next_ijk_U0_write_r_din;
wire    tdf11_get_next_ijk_U0_write_r_write;
wire    tdf11_readInputs75_U0_ap_start;
wire    tdf11_readInputs75_U0_ap_done;
wire    tdf11_readInputs75_U0_ap_continue;
wire    tdf11_readInputs75_U0_ap_idle;
wire    tdf11_readInputs75_U0_ap_ready;
wire   [11:0] tdf11_readInputs75_U0_in_data_address0;
wire    tdf11_readInputs75_U0_in_data_ce0;
wire    tdf11_readInputs75_U0_indices_01_read;
wire    tdf11_readInputs75_U0_indices_12_read;
wire   [9:0] tdf11_readInputs75_U0_ifmap_vec_address0;
wire    tdf11_readInputs75_U0_ifmap_vec_ce0;
wire    tdf11_readInputs75_U0_ifmap_vec_we0;
wire   [15:0] tdf11_readInputs75_U0_ifmap_vec_d0;
wire   [9:0] tdf11_readInputs75_U0_ifmap_vec_address1;
wire    tdf11_readInputs75_U0_ifmap_vec_ce1;
wire    tdf11_readInputs75_U0_ifmap_vec_we1;
wire   [15:0] tdf11_readInputs75_U0_ifmap_vec_d1;
wire   [3:0] tdf11_readInputs75_U0_indices_01_out_din;
wire    tdf11_readInputs75_U0_indices_01_out_write;
wire   [7:0] tdf11_readInputs75_U0_indices_12_out_din;
wire    tdf11_readInputs75_U0_indices_12_out_write;
wire    tdf11_readInputs75_U0_in_data_full_n;
wire    tdf11_readInputs75_U0_in_data_write;
wire    ap_channel_done_ifmap_vec;
wire    tdf11_readInputs75_U0_ifmap_vec_full_n;
wire    tdf11_readFilters74_U0_ap_start;
wire    tdf11_readFilters74_U0_ap_done;
wire    tdf11_readFilters74_U0_ap_continue;
wire    tdf11_readFilters74_U0_ap_idle;
wire    tdf11_readFilters74_U0_ap_ready;
wire   [16:0] tdf11_readFilters74_U0_filter_data_address0;
wire    tdf11_readFilters74_U0_filter_data_ce0;
wire    tdf11_readFilters74_U0_indices_23_read;
wire   [9:0] tdf11_readFilters74_U0_weight_vecs_0_address0;
wire    tdf11_readFilters74_U0_weight_vecs_0_ce0;
wire    tdf11_readFilters74_U0_weight_vecs_0_we0;
wire   [15:0] tdf11_readFilters74_U0_weight_vecs_0_d0;
wire   [9:0] tdf11_readFilters74_U0_weight_vecs_0_address1;
wire    tdf11_readFilters74_U0_weight_vecs_0_ce1;
wire    tdf11_readFilters74_U0_weight_vecs_0_we1;
wire   [15:0] tdf11_readFilters74_U0_weight_vecs_0_d1;
wire    ap_channel_done_weight_vecs_0;
wire    tdf11_readFilters74_U0_weight_vecs_0_full_n;
wire    tdf11_dot_product_U0_ap_start;
wire    tdf11_dot_product_U0_ap_done;
wire    tdf11_dot_product_U0_ap_continue;
wire    tdf11_dot_product_U0_ap_idle;
wire    tdf11_dot_product_U0_ap_ready;
wire   [9:0] tdf11_dot_product_U0_ifmap_vec_address0;
wire    tdf11_dot_product_U0_ifmap_vec_ce0;
wire   [9:0] tdf11_dot_product_U0_weight_vecs_0_address0;
wire    tdf11_dot_product_U0_weight_vecs_0_ce0;
wire   [9:0] tdf11_dot_product_U0_products_0_address0;
wire    tdf11_dot_product_U0_products_0_ce0;
wire    tdf11_dot_product_U0_products_0_we0;
wire   [15:0] tdf11_dot_product_U0_products_0_d0;
wire    ap_channel_done_products_0;
wire    tdf11_dot_product_U0_products_0_full_n;
wire    tdf11_accum_1_U0_ap_start;
wire    tdf11_accum_1_U0_ap_done;
wire    tdf11_accum_1_U0_ap_continue;
wire    tdf11_accum_1_U0_ap_idle;
wire    tdf11_accum_1_U0_ap_ready;
wire   [9:0] tdf11_accum_1_U0_accum_in_0_address0;
wire    tdf11_accum_1_U0_accum_in_0_ce0;
wire   [9:0] tdf11_accum_1_U0_accum_in_0_address1;
wire    tdf11_accum_1_U0_accum_in_0_ce1;
wire   [2:0] tdf11_accum_1_U0_accum_out_address0;
wire    tdf11_accum_1_U0_accum_out_ce0;
wire    tdf11_accum_1_U0_accum_out_we0;
wire   [15:0] tdf11_accum_1_U0_accum_out_d0;
wire   [2:0] tdf11_accum_1_U0_accum_out_address1;
wire    tdf11_accum_1_U0_accum_out_ce1;
wire    tdf11_accum_1_U0_accum_out_we1;
wire   [15:0] tdf11_accum_1_U0_accum_out_d1;
wire    ap_channel_done_accum1_out_0;
wire    tdf11_accum_1_U0_accum_out_full_n;
wire    tdf11_accum_2_U0_ap_start;
wire    tdf11_accum_2_U0_ap_done;
wire    tdf11_accum_2_U0_ap_continue;
wire    tdf11_accum_2_U0_ap_idle;
wire    tdf11_accum_2_U0_ap_ready;
wire   [15:0] tdf11_accum_2_U0_accum_in_22;
wire    tdf11_accum_2_U0_accum_in_22_ap_vld;
wire   [2:0] tdf11_accum_2_U0_accum_in_address0;
wire    tdf11_accum_2_U0_accum_in_ce0;
wire    ap_channel_done_tmp_channel;
wire    tmp_channel_full_n;
wire    Block_entry_proc_proc441_U0_ap_start;
wire    Block_entry_proc_proc441_U0_ap_done;
wire    Block_entry_proc_proc441_U0_ap_continue;
wire    Block_entry_proc_proc441_U0_ap_idle;
wire    Block_entry_proc_proc441_U0_ap_ready;
wire   [15:0] Block_entry_proc_proc441_U0_ap_return;
wire    ap_channel_done_sums_0;
wire    sums_0_full_n;
wire    tdf11_adjust_U0_ap_start;
wire    tdf11_adjust_U0_ap_done;
wire    tdf11_adjust_U0_ap_continue;
wire    tdf11_adjust_U0_ap_idle;
wire    tdf11_adjust_U0_ap_ready;
wire   [8:0] tdf11_adjust_U0_adjustments_address0;
wire    tdf11_adjust_U0_adjustments_ce0;
wire    tdf11_adjust_U0_indices_23_read;
wire   [8:0] tdf11_adjust_U0_indices_23_out_din;
wire    tdf11_adjust_U0_indices_23_out_write;
wire   [15:0] tdf11_adjust_U0_ap_return;
wire    ap_channel_done_intermediate_fmaps_0;
wire    intermediate_fmaps_0_full_n;
wire    tdf11_l2_multiply72_U0_ap_start;
wire    tdf11_l2_multiply72_U0_ap_done;
wire    tdf11_l2_multiply72_U0_ap_continue;
wire    tdf11_l2_multiply72_U0_ap_idle;
wire    tdf11_l2_multiply72_U0_ap_ready;
wire   [15:0] tdf11_l2_multiply72_U0_l2_filter_data_address0;
wire    tdf11_l2_multiply72_U0_l2_filter_data_ce0;
wire   [6:0] tdf11_l2_multiply72_U0_l2_products_address0;
wire    tdf11_l2_multiply72_U0_l2_products_ce0;
wire    tdf11_l2_multiply72_U0_l2_products_we0;
wire   [15:0] tdf11_l2_multiply72_U0_l2_products_d0;
wire    tdf11_l2_multiply72_U0_indices_23_read;
wire    ap_channel_done_l2_products;
wire    tdf11_l2_multiply72_U0_l2_products_full_n;
wire    tdf11_l2_writeOutputs_171_U0_ap_start;
wire    tdf11_l2_writeOutputs_171_U0_ap_done;
wire    tdf11_l2_writeOutputs_171_U0_ap_continue;
wire    tdf11_l2_writeOutputs_171_U0_ap_idle;
wire    tdf11_l2_writeOutputs_171_U0_ap_ready;
wire    tdf11_l2_writeOutputs_171_U0_indices_01_read;
wire    tdf11_l2_writeOutputs_171_U0_indices_12_read;
wire    tdf11_l2_writeOutputs_171_U0_write4_read;
wire   [6:0] tdf11_l2_writeOutputs_171_U0_l2_partial_sums_address0;
wire    tdf11_l2_writeOutputs_171_U0_l2_partial_sums_ce0;
wire   [12:0] tdf11_l2_writeOutputs_171_U0_out_data_address1;
wire    tdf11_l2_writeOutputs_171_U0_out_data_ce1;
wire    tdf11_l2_writeOutputs_171_U0_out_data_we1;
wire   [63:0] tdf11_l2_writeOutputs_171_U0_out_data_d1;
wire   [6:0] tdf11_l2_writeOutputs_171_U0_l2_adjustments_address0;
wire    tdf11_l2_writeOutputs_171_U0_l2_adjustments_ce0;
wire    tdf11_l2_writeOutputs_171_U0_out_data_full_n;
wire    tdf11_l2_writeOutputs_171_U0_out_data_write;
wire    ap_sync_continue;
wire    ifmap_vec_i_full_n;
wire    ifmap_vec_t_empty_n;
wire    weight_vecs_0_i_full_n;
wire    weight_vecs_0_t_empty_n;
wire    products_0_i_full_n;
wire    products_0_t_empty_n;
wire   [15:0] products_0_t_d1;
wire    products_0_t_we1;
wire    accum1_out_0_i_full_n;
wire    accum1_out_0_t_empty_n;
wire    l2_products_i_full_n;
wire    l2_products_t_empty_n;
wire    indices_01_c_full_n;
wire   [15:0] indices_01_c_dout;
wire    indices_01_c_empty_n;
wire    indices_12_c_full_n;
wire   [15:0] indices_12_c_dout;
wire    indices_12_c_empty_n;
wire    indices_23_c_full_n;
wire   [8:0] indices_23_c_dout;
wire    indices_23_c_empty_n;
wire    indices_23_c1_full_n;
wire   [8:0] indices_23_c1_dout;
wire    indices_23_c1_empty_n;
wire   [0:0] write4_c_din;
wire    write4_c_full_n;
wire   [0:0] write4_c_dout;
wire    write4_c_empty_n;
wire    indices_01_c2_full_n;
wire   [3:0] indices_01_c2_dout;
wire    indices_01_c2_empty_n;
wire    indices_12_c3_full_n;
wire   [7:0] indices_12_c3_dout;
wire    indices_12_c3_empty_n;
wire   [15:0] tmp_channel_dout;
wire    tmp_channel_empty_n;
wire   [15:0] sums_0_dout;
wire    sums_0_empty_n;
wire    indices_23_c4_full_n;
wire   [8:0] indices_23_c4_dout;
wire    indices_23_c4_empty_n;
wire   [15:0] intermediate_fmaps_0_dout;
wire    intermediate_fmaps_0_empty_n;
wire    ap_sync_done;
wire    ap_sync_ready;
reg    ap_sync_reg_tdf11_get_next_ijk_U0_ap_ready;
wire    ap_sync_tdf11_get_next_ijk_U0_ap_ready;
reg    ap_sync_reg_tdf11_readInputs75_U0_ap_ready;
wire    ap_sync_tdf11_readInputs75_U0_ap_ready;
wire   [0:0] start_for_tdf11_readFilters74_U0_din;
wire    start_for_tdf11_readFilters74_U0_full_n;
wire   [0:0] start_for_tdf11_readFilters74_U0_dout;
wire    start_for_tdf11_readFilters74_U0_empty_n;
wire    tdf11_readInputs75_U0_start_full_n;
wire    tdf11_readInputs75_U0_start_write;
wire    tdf11_readFilters74_U0_start_full_n;
wire    tdf11_readFilters74_U0_start_write;
wire    tdf11_dot_product_U0_start_full_n;
wire    tdf11_dot_product_U0_start_write;
wire    tdf11_accum_1_U0_start_full_n;
wire    tdf11_accum_1_U0_start_write;
wire    tdf11_accum_2_U0_start_full_n;
wire    tdf11_accum_2_U0_start_write;
wire    Block_entry_proc_proc441_U0_start_full_n;
wire    Block_entry_proc_proc441_U0_start_write;
wire    tdf11_adjust_U0_start_full_n;
wire    tdf11_adjust_U0_start_write;
wire    tdf11_l2_multiply72_U0_start_full_n;
wire    tdf11_l2_multiply72_U0_start_write;
wire    tdf11_l2_writeOutputs_171_U0_start_full_n;
wire    tdf11_l2_writeOutputs_171_U0_start_write;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_sync_reg_tdf11_get_next_ijk_U0_ap_ready = 1'b0;
#0 ap_sync_reg_tdf11_readInputs75_U0_ap_ready = 1'b0;
end

td_fused_top_dataflow_in_loop_TOP_LOOP38270_ifmap_vec #(
    .DataWidth( 16 ),
    .AddressRange( 576 ),
    .AddressWidth( 10 ))
ifmap_vec_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf11_readInputs75_U0_ap_done),
    .i_full_n(ifmap_vec_i_full_n),
    .i_ce0(tdf11_readInputs75_U0_ifmap_vec_ce0),
    .i_we0(tdf11_readInputs75_U0_ifmap_vec_we0),
    .i_address0(tdf11_readInputs75_U0_ifmap_vec_address0),
    .i_d0(tdf11_readInputs75_U0_ifmap_vec_d0),
    .i_q0(ifmap_vec_i_q0),
    .i_ce1(tdf11_readInputs75_U0_ifmap_vec_ce1),
    .i_we1(tdf11_readInputs75_U0_ifmap_vec_we1),
    .i_address1(tdf11_readInputs75_U0_ifmap_vec_address1),
    .i_d1(tdf11_readInputs75_U0_ifmap_vec_d1),
    .t_ce(1'b1),
    .t_read(tdf11_dot_product_U0_ap_ready),
    .t_empty_n(ifmap_vec_t_empty_n),
    .t_ce0(tdf11_dot_product_U0_ifmap_vec_ce0),
    .t_we0(1'b0),
    .t_address0(tdf11_dot_product_U0_ifmap_vec_address0),
    .t_d0(16'd0),
    .t_q0(ifmap_vec_t_q0),
    .t_ce1(1'b0),
    .t_we1(1'b0),
    .t_address1(10'd0),
    .t_d1(16'd0)
);

td_fused_top_dataflow_in_loop_TOP_LOOP38270_ifmap_vec #(
    .DataWidth( 16 ),
    .AddressRange( 576 ),
    .AddressWidth( 10 ))
weight_vecs_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf11_readFilters74_U0_ap_done),
    .i_full_n(weight_vecs_0_i_full_n),
    .i_ce0(tdf11_readFilters74_U0_weight_vecs_0_ce0),
    .i_we0(tdf11_readFilters74_U0_weight_vecs_0_we0),
    .i_address0(tdf11_readFilters74_U0_weight_vecs_0_address0),
    .i_d0(tdf11_readFilters74_U0_weight_vecs_0_d0),
    .i_q0(weight_vecs_0_i_q0),
    .i_ce1(tdf11_readFilters74_U0_weight_vecs_0_ce1),
    .i_we1(tdf11_readFilters74_U0_weight_vecs_0_we1),
    .i_address1(tdf11_readFilters74_U0_weight_vecs_0_address1),
    .i_d1(tdf11_readFilters74_U0_weight_vecs_0_d1),
    .t_ce(1'b1),
    .t_read(tdf11_dot_product_U0_ap_ready),
    .t_empty_n(weight_vecs_0_t_empty_n),
    .t_ce0(tdf11_dot_product_U0_weight_vecs_0_ce0),
    .t_we0(1'b0),
    .t_address0(tdf11_dot_product_U0_weight_vecs_0_address0),
    .t_d0(16'd0),
    .t_q0(weight_vecs_0_t_q0),
    .t_ce1(1'b0),
    .t_we1(1'b0),
    .t_address1(10'd0),
    .t_d1(16'd0)
);

td_fused_top_dataflow_in_loop_TOP_LOOP38270_products_0 #(
    .DataWidth( 16 ),
    .AddressRange( 576 ),
    .AddressWidth( 10 ))
products_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf11_dot_product_U0_ap_done),
    .i_full_n(products_0_i_full_n),
    .i_ce0(tdf11_dot_product_U0_products_0_ce0),
    .i_we0(tdf11_dot_product_U0_products_0_we0),
    .i_address0(tdf11_dot_product_U0_products_0_address0),
    .i_d0(tdf11_dot_product_U0_products_0_d0),
    .i_q0(products_0_i_q0),
    .i_ce1(1'b0),
    .i_address1(10'd0),
    .i_q1(products_0_i_q1),
    .t_ce(1'b1),
    .t_read(tdf11_accum_1_U0_ap_ready),
    .t_empty_n(products_0_t_empty_n),
    .t_ce0(tdf11_accum_1_U0_accum_in_0_ce0),
    .t_we0(1'b0),
    .t_address0(tdf11_accum_1_U0_accum_in_0_address0),
    .t_d0(16'd0),
    .t_q0(products_0_t_q0),
    .t_ce1(tdf11_accum_1_U0_accum_in_0_ce1),
    .t_address1(tdf11_accum_1_U0_accum_in_0_address1),
    .t_q1(products_0_t_q1)
);

td_fused_top_dataflow_in_loop_TOP_LOOP38270_accum1_out_0 #(
    .DataWidth( 16 ),
    .AddressRange( 8 ),
    .AddressWidth( 3 ))
accum1_out_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf11_accum_1_U0_ap_done),
    .i_full_n(accum1_out_0_i_full_n),
    .i_ce0(tdf11_accum_1_U0_accum_out_ce0),
    .i_we0(tdf11_accum_1_U0_accum_out_we0),
    .i_address0(tdf11_accum_1_U0_accum_out_address0),
    .i_d0(tdf11_accum_1_U0_accum_out_d0),
    .i_q0(accum1_out_0_i_q0),
    .i_ce1(tdf11_accum_1_U0_accum_out_ce1),
    .i_we1(tdf11_accum_1_U0_accum_out_we1),
    .i_address1(tdf11_accum_1_U0_accum_out_address1),
    .i_d1(tdf11_accum_1_U0_accum_out_d1),
    .t_ce(1'b1),
    .t_read(tdf11_accum_2_U0_ap_ready),
    .t_empty_n(accum1_out_0_t_empty_n),
    .t_ce0(tdf11_accum_2_U0_accum_in_ce0),
    .t_we0(1'b0),
    .t_address0(tdf11_accum_2_U0_accum_in_address0),
    .t_d0(16'd0),
    .t_q0(accum1_out_0_t_q0),
    .t_ce1(1'b0),
    .t_we1(1'b0),
    .t_address1(3'd0),
    .t_d1(16'd0)
);

td_fused_top_dataflow_in_loop_TOP_LOOP38270_l2_products #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
l2_products_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf11_l2_multiply72_U0_ap_done),
    .i_full_n(l2_products_i_full_n),
    .i_ce0(tdf11_l2_multiply72_U0_l2_products_ce0),
    .i_we0(tdf11_l2_multiply72_U0_l2_products_we0),
    .i_address0(tdf11_l2_multiply72_U0_l2_products_address0),
    .i_d0(tdf11_l2_multiply72_U0_l2_products_d0),
    .i_q0(l2_products_i_q0),
    .t_ce(1'b1),
    .t_read(tdf11_l2_writeOutputs_171_U0_ap_ready),
    .t_empty_n(l2_products_t_empty_n),
    .t_ce0(tdf11_l2_writeOutputs_171_U0_l2_partial_sums_ce0),
    .t_we0(1'b0),
    .t_address0(tdf11_l2_writeOutputs_171_U0_l2_partial_sums_address0),
    .t_d0(16'd0),
    .t_q0(l2_products_t_q0)
);

td_fused_top_tdf11_get_next_ijk tdf11_get_next_ijk_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf11_get_next_ijk_U0_ap_start),
    .start_full_n(start_for_tdf11_readFilters74_U0_full_n),
    .ap_done(tdf11_get_next_ijk_U0_ap_done),
    .ap_continue(tdf11_get_next_ijk_U0_ap_continue),
    .ap_idle(tdf11_get_next_ijk_U0_ap_idle),
    .ap_ready(tdf11_get_next_ijk_U0_ap_ready),
    .start_out(tdf11_get_next_ijk_U0_start_out),
    .start_write(tdf11_get_next_ijk_U0_start_write),
    .indices_0_din(tdf11_get_next_ijk_U0_indices_0_din),
    .indices_0_full_n(indices_01_c_full_n),
    .indices_0_write(tdf11_get_next_ijk_U0_indices_0_write),
    .indices_1_din(tdf11_get_next_ijk_U0_indices_1_din),
    .indices_1_full_n(indices_12_c_full_n),
    .indices_1_write(tdf11_get_next_ijk_U0_indices_1_write),
    .indices_2_out_din(tdf11_get_next_ijk_U0_indices_2_out_din),
    .indices_2_out_full_n(indices_23_c_full_n),
    .indices_2_out_write(tdf11_get_next_ijk_U0_indices_2_out_write),
    .indices_2_out1_din(tdf11_get_next_ijk_U0_indices_2_out1_din),
    .indices_2_out1_full_n(indices_23_c1_full_n),
    .indices_2_out1_write(tdf11_get_next_ijk_U0_indices_2_out1_write),
    .write_r_din(tdf11_get_next_ijk_U0_write_r_din),
    .write_r_full_n(write4_c_full_n),
    .write_r_write(tdf11_get_next_ijk_U0_write_r_write)
);

td_fused_top_tdf11_readInputs75 tdf11_readInputs75_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf11_readInputs75_U0_ap_start),
    .ap_done(tdf11_readInputs75_U0_ap_done),
    .ap_continue(tdf11_readInputs75_U0_ap_continue),
    .ap_idle(tdf11_readInputs75_U0_ap_idle),
    .ap_ready(tdf11_readInputs75_U0_ap_ready),
    .in_data_address0(tdf11_readInputs75_U0_in_data_address0),
    .in_data_ce0(tdf11_readInputs75_U0_in_data_ce0),
    .in_data_q0(in_data_q0),
    .indices_01_dout(indices_01_c_dout),
    .indices_01_empty_n(indices_01_c_empty_n),
    .indices_01_read(tdf11_readInputs75_U0_indices_01_read),
    .indices_12_dout(indices_12_c_dout),
    .indices_12_empty_n(indices_12_c_empty_n),
    .indices_12_read(tdf11_readInputs75_U0_indices_12_read),
    .ifmap_vec_address0(tdf11_readInputs75_U0_ifmap_vec_address0),
    .ifmap_vec_ce0(tdf11_readInputs75_U0_ifmap_vec_ce0),
    .ifmap_vec_we0(tdf11_readInputs75_U0_ifmap_vec_we0),
    .ifmap_vec_d0(tdf11_readInputs75_U0_ifmap_vec_d0),
    .ifmap_vec_address1(tdf11_readInputs75_U0_ifmap_vec_address1),
    .ifmap_vec_ce1(tdf11_readInputs75_U0_ifmap_vec_ce1),
    .ifmap_vec_we1(tdf11_readInputs75_U0_ifmap_vec_we1),
    .ifmap_vec_d1(tdf11_readInputs75_U0_ifmap_vec_d1),
    .indices_01_out_din(tdf11_readInputs75_U0_indices_01_out_din),
    .indices_01_out_full_n(indices_01_c2_full_n),
    .indices_01_out_write(tdf11_readInputs75_U0_indices_01_out_write),
    .indices_12_out_din(tdf11_readInputs75_U0_indices_12_out_din),
    .indices_12_out_full_n(indices_12_c3_full_n),
    .indices_12_out_write(tdf11_readInputs75_U0_indices_12_out_write)
);

td_fused_top_tdf11_readFilters74 tdf11_readFilters74_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf11_readFilters74_U0_ap_start),
    .ap_done(tdf11_readFilters74_U0_ap_done),
    .ap_continue(tdf11_readFilters74_U0_ap_continue),
    .ap_idle(tdf11_readFilters74_U0_ap_idle),
    .ap_ready(tdf11_readFilters74_U0_ap_ready),
    .filter_data_address0(tdf11_readFilters74_U0_filter_data_address0),
    .filter_data_ce0(tdf11_readFilters74_U0_filter_data_ce0),
    .filter_data_q0(l1_filter_data_q0),
    .indices_23_dout(indices_23_c_dout),
    .indices_23_empty_n(indices_23_c_empty_n),
    .indices_23_read(tdf11_readFilters74_U0_indices_23_read),
    .weight_vecs_0_address0(tdf11_readFilters74_U0_weight_vecs_0_address0),
    .weight_vecs_0_ce0(tdf11_readFilters74_U0_weight_vecs_0_ce0),
    .weight_vecs_0_we0(tdf11_readFilters74_U0_weight_vecs_0_we0),
    .weight_vecs_0_d0(tdf11_readFilters74_U0_weight_vecs_0_d0),
    .weight_vecs_0_address1(tdf11_readFilters74_U0_weight_vecs_0_address1),
    .weight_vecs_0_ce1(tdf11_readFilters74_U0_weight_vecs_0_ce1),
    .weight_vecs_0_we1(tdf11_readFilters74_U0_weight_vecs_0_we1),
    .weight_vecs_0_d1(tdf11_readFilters74_U0_weight_vecs_0_d1)
);

td_fused_top_tdf11_dot_product tdf11_dot_product_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf11_dot_product_U0_ap_start),
    .ap_done(tdf11_dot_product_U0_ap_done),
    .ap_continue(tdf11_dot_product_U0_ap_continue),
    .ap_idle(tdf11_dot_product_U0_ap_idle),
    .ap_ready(tdf11_dot_product_U0_ap_ready),
    .ifmap_vec_address0(tdf11_dot_product_U0_ifmap_vec_address0),
    .ifmap_vec_ce0(tdf11_dot_product_U0_ifmap_vec_ce0),
    .ifmap_vec_q0(ifmap_vec_t_q0),
    .weight_vecs_0_address0(tdf11_dot_product_U0_weight_vecs_0_address0),
    .weight_vecs_0_ce0(tdf11_dot_product_U0_weight_vecs_0_ce0),
    .weight_vecs_0_q0(weight_vecs_0_t_q0),
    .products_0_address0(tdf11_dot_product_U0_products_0_address0),
    .products_0_ce0(tdf11_dot_product_U0_products_0_ce0),
    .products_0_we0(tdf11_dot_product_U0_products_0_we0),
    .products_0_d0(tdf11_dot_product_U0_products_0_d0)
);

td_fused_top_tdf11_accum_1 tdf11_accum_1_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf11_accum_1_U0_ap_start),
    .ap_done(tdf11_accum_1_U0_ap_done),
    .ap_continue(tdf11_accum_1_U0_ap_continue),
    .ap_idle(tdf11_accum_1_U0_ap_idle),
    .ap_ready(tdf11_accum_1_U0_ap_ready),
    .accum_in_0_address0(tdf11_accum_1_U0_accum_in_0_address0),
    .accum_in_0_ce0(tdf11_accum_1_U0_accum_in_0_ce0),
    .accum_in_0_q0(products_0_t_q0),
    .accum_in_0_address1(tdf11_accum_1_U0_accum_in_0_address1),
    .accum_in_0_ce1(tdf11_accum_1_U0_accum_in_0_ce1),
    .accum_in_0_q1(products_0_t_q1),
    .accum_out_address0(tdf11_accum_1_U0_accum_out_address0),
    .accum_out_ce0(tdf11_accum_1_U0_accum_out_ce0),
    .accum_out_we0(tdf11_accum_1_U0_accum_out_we0),
    .accum_out_d0(tdf11_accum_1_U0_accum_out_d0),
    .accum_out_address1(tdf11_accum_1_U0_accum_out_address1),
    .accum_out_ce1(tdf11_accum_1_U0_accum_out_ce1),
    .accum_out_we1(tdf11_accum_1_U0_accum_out_we1),
    .accum_out_d1(tdf11_accum_1_U0_accum_out_d1)
);

td_fused_top_tdf11_accum_2 tdf11_accum_2_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf11_accum_2_U0_ap_start),
    .ap_done(tdf11_accum_2_U0_ap_done),
    .ap_continue(tdf11_accum_2_U0_ap_continue),
    .ap_idle(tdf11_accum_2_U0_ap_idle),
    .ap_ready(tdf11_accum_2_U0_ap_ready),
    .accum_in_22(tdf11_accum_2_U0_accum_in_22),
    .accum_in_22_ap_vld(tdf11_accum_2_U0_accum_in_22_ap_vld),
    .accum_in_address0(tdf11_accum_2_U0_accum_in_address0),
    .accum_in_ce0(tdf11_accum_2_U0_accum_in_ce0),
    .accum_in_q0(accum1_out_0_t_q0)
);

td_fused_top_Block_entry_proc_proc441 Block_entry_proc_proc441_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(Block_entry_proc_proc441_U0_ap_start),
    .ap_done(Block_entry_proc_proc441_U0_ap_done),
    .ap_continue(Block_entry_proc_proc441_U0_ap_continue),
    .ap_idle(Block_entry_proc_proc441_U0_ap_idle),
    .ap_ready(Block_entry_proc_proc441_U0_ap_ready),
    .tmp(tmp_channel_dout),
    .ap_return(Block_entry_proc_proc441_U0_ap_return)
);

td_fused_top_tdf11_adjust tdf11_adjust_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf11_adjust_U0_ap_start),
    .ap_done(tdf11_adjust_U0_ap_done),
    .ap_continue(tdf11_adjust_U0_ap_continue),
    .ap_idle(tdf11_adjust_U0_ap_idle),
    .ap_ready(tdf11_adjust_U0_ap_ready),
    .sums_read(sums_0_dout),
    .adjustments_address0(tdf11_adjust_U0_adjustments_address0),
    .adjustments_ce0(tdf11_adjust_U0_adjustments_ce0),
    .adjustments_q0(l1_adjustments_q0),
    .indices_23_dout(indices_23_c1_dout),
    .indices_23_empty_n(indices_23_c1_empty_n),
    .indices_23_read(tdf11_adjust_U0_indices_23_read),
    .indices_23_out_din(tdf11_adjust_U0_indices_23_out_din),
    .indices_23_out_full_n(indices_23_c4_full_n),
    .indices_23_out_write(tdf11_adjust_U0_indices_23_out_write),
    .ap_return(tdf11_adjust_U0_ap_return)
);

td_fused_top_tdf11_l2_multiply72 tdf11_l2_multiply72_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf11_l2_multiply72_U0_ap_start),
    .ap_done(tdf11_l2_multiply72_U0_ap_done),
    .ap_continue(tdf11_l2_multiply72_U0_ap_continue),
    .ap_idle(tdf11_l2_multiply72_U0_ap_idle),
    .ap_ready(tdf11_l2_multiply72_U0_ap_ready),
    .intermediate_fmaps_read(intermediate_fmaps_0_dout),
    .l2_filter_data_address0(tdf11_l2_multiply72_U0_l2_filter_data_address0),
    .l2_filter_data_ce0(tdf11_l2_multiply72_U0_l2_filter_data_ce0),
    .l2_filter_data_q0(l2_filter_data_q0),
    .l2_products_address0(tdf11_l2_multiply72_U0_l2_products_address0),
    .l2_products_ce0(tdf11_l2_multiply72_U0_l2_products_ce0),
    .l2_products_we0(tdf11_l2_multiply72_U0_l2_products_we0),
    .l2_products_d0(tdf11_l2_multiply72_U0_l2_products_d0),
    .indices_23_dout(indices_23_c4_dout),
    .indices_23_empty_n(indices_23_c4_empty_n),
    .indices_23_read(tdf11_l2_multiply72_U0_indices_23_read)
);

td_fused_top_tdf11_l2_writeOutputs_171 tdf11_l2_writeOutputs_171_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf11_l2_writeOutputs_171_U0_ap_start),
    .ap_done(tdf11_l2_writeOutputs_171_U0_ap_done),
    .ap_continue(tdf11_l2_writeOutputs_171_U0_ap_continue),
    .ap_idle(tdf11_l2_writeOutputs_171_U0_ap_idle),
    .ap_ready(tdf11_l2_writeOutputs_171_U0_ap_ready),
    .indices_01_dout(indices_01_c2_dout),
    .indices_01_empty_n(indices_01_c2_empty_n),
    .indices_01_read(tdf11_l2_writeOutputs_171_U0_indices_01_read),
    .indices_12_dout(indices_12_c3_dout),
    .indices_12_empty_n(indices_12_c3_empty_n),
    .indices_12_read(tdf11_l2_writeOutputs_171_U0_indices_12_read),
    .write4_dout(write4_c_dout),
    .write4_empty_n(write4_c_empty_n),
    .write4_read(tdf11_l2_writeOutputs_171_U0_write4_read),
    .l2_partial_sums_address0(tdf11_l2_writeOutputs_171_U0_l2_partial_sums_address0),
    .l2_partial_sums_ce0(tdf11_l2_writeOutputs_171_U0_l2_partial_sums_ce0),
    .l2_partial_sums_q0(l2_products_t_q0),
    .out_data_address1(tdf11_l2_writeOutputs_171_U0_out_data_address1),
    .out_data_ce1(tdf11_l2_writeOutputs_171_U0_out_data_ce1),
    .out_data_we1(tdf11_l2_writeOutputs_171_U0_out_data_we1),
    .out_data_d1(tdf11_l2_writeOutputs_171_U0_out_data_d1),
    .l2_adjustments_address0(tdf11_l2_writeOutputs_171_U0_l2_adjustments_address0),
    .l2_adjustments_ce0(tdf11_l2_writeOutputs_171_U0_l2_adjustments_ce0),
    .l2_adjustments_q0(l2_adjustments_q0)
);

td_fused_top_fifo_w16_d2_S_x8 indices_01_c_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(indices_01_c_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf11_readInputs75_U0_indices_01_read),
    .if_dout(indices_01_c_dout),
    .if_full_n(indices_01_c_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf11_get_next_ijk_U0_indices_0_write),
    .if_din(tdf11_get_next_ijk_U0_indices_0_din)
);

td_fused_top_fifo_w16_d2_S_x8 indices_12_c_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(indices_12_c_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf11_readInputs75_U0_indices_12_read),
    .if_dout(indices_12_c_dout),
    .if_full_n(indices_12_c_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf11_get_next_ijk_U0_indices_1_write),
    .if_din(tdf11_get_next_ijk_U0_indices_1_din)
);

td_fused_top_fifo_w9_d2_S_x indices_23_c_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(indices_23_c_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf11_readFilters74_U0_indices_23_read),
    .if_dout(indices_23_c_dout),
    .if_full_n(indices_23_c_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf11_get_next_ijk_U0_indices_2_out_write),
    .if_din(tdf11_get_next_ijk_U0_indices_2_out_din)
);

td_fused_top_fifo_w9_d7_S indices_23_c1_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(indices_23_c1_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf11_adjust_U0_indices_23_read),
    .if_dout(indices_23_c1_dout),
    .if_full_n(indices_23_c1_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf11_get_next_ijk_U0_indices_2_out1_write),
    .if_din(tdf11_get_next_ijk_U0_indices_2_out1_din)
);

td_fused_top_fifo_w1_d9_S_x2 write4_c_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(write4_c_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf11_l2_writeOutputs_171_U0_write4_read),
    .if_dout(write4_c_dout),
    .if_full_n(write4_c_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf11_get_next_ijk_U0_write_r_write),
    .if_din(write4_c_din)
);

td_fused_top_fifo_w4_d8_S_x1 indices_01_c2_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(indices_01_c2_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf11_l2_writeOutputs_171_U0_indices_01_read),
    .if_dout(indices_01_c2_dout),
    .if_full_n(indices_01_c2_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf11_readInputs75_U0_indices_01_out_write),
    .if_din(tdf11_readInputs75_U0_indices_01_out_din)
);

td_fused_top_fifo_w8_d8_S_x0 indices_12_c3_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(indices_12_c3_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf11_l2_writeOutputs_171_U0_indices_12_read),
    .if_dout(indices_12_c3_dout),
    .if_full_n(indices_12_c3_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf11_readInputs75_U0_indices_12_out_write),
    .if_din(tdf11_readInputs75_U0_indices_12_out_din)
);

td_fused_top_fifo_w16_d2_S_x8 tmp_channel_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(tmp_channel_empty_n),
    .if_read_ce(1'b1),
    .if_read(Block_entry_proc_proc441_U0_ap_ready),
    .if_dout(tmp_channel_dout),
    .if_full_n(tmp_channel_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf11_accum_2_U0_ap_done),
    .if_din(tdf11_accum_2_U0_accum_in_22)
);

td_fused_top_fifo_w16_d2_S_x8 sums_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(sums_0_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf11_adjust_U0_ap_ready),
    .if_dout(sums_0_dout),
    .if_full_n(sums_0_full_n),
    .if_write_ce(1'b1),
    .if_write(Block_entry_proc_proc441_U0_ap_done),
    .if_din(Block_entry_proc_proc441_U0_ap_return)
);

td_fused_top_fifo_w9_d2_S_x indices_23_c4_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(indices_23_c4_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf11_l2_multiply72_U0_indices_23_read),
    .if_dout(indices_23_c4_dout),
    .if_full_n(indices_23_c4_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf11_adjust_U0_indices_23_out_write),
    .if_din(tdf11_adjust_U0_indices_23_out_din)
);

td_fused_top_fifo_w16_d2_S_x8 intermediate_fmaps_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(intermediate_fmaps_0_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf11_l2_multiply72_U0_ap_ready),
    .if_dout(intermediate_fmaps_0_dout),
    .if_full_n(intermediate_fmaps_0_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf11_adjust_U0_ap_done),
    .if_din(tdf11_adjust_U0_ap_return)
);

td_fused_top_start_for_tdf11_readFilters74_U0 start_for_tdf11_readFilters74_U0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(start_for_tdf11_readFilters74_U0_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf11_readFilters74_U0_ap_ready),
    .if_dout(start_for_tdf11_readFilters74_U0_dout),
    .if_full_n(start_for_tdf11_readFilters74_U0_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf11_get_next_ijk_U0_start_write),
    .if_din(start_for_tdf11_readFilters74_U0_din)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_sync_reg_tdf11_get_next_ijk_U0_ap_ready <= 1'b0;
    end else begin
        if (((ap_sync_ready & ap_start) == 1'b1)) begin
            ap_sync_reg_tdf11_get_next_ijk_U0_ap_ready <= 1'b0;
        end else begin
            ap_sync_reg_tdf11_get_next_ijk_U0_ap_ready <= ap_sync_tdf11_get_next_ijk_U0_ap_ready;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_sync_reg_tdf11_readInputs75_U0_ap_ready <= 1'b0;
    end else begin
        if (((ap_sync_ready & ap_start) == 1'b1)) begin
            ap_sync_reg_tdf11_readInputs75_U0_ap_ready <= 1'b0;
        end else begin
            ap_sync_reg_tdf11_readInputs75_U0_ap_ready <= ap_sync_tdf11_readInputs75_U0_ap_ready;
        end
    end
end

assign Block_entry_proc_proc441_U0_ap_continue = sums_0_full_n;

assign Block_entry_proc_proc441_U0_ap_start = tmp_channel_empty_n;

assign Block_entry_proc_proc441_U0_start_full_n = 1'b1;

assign Block_entry_proc_proc441_U0_start_write = 1'b0;

assign ap_channel_done_accum1_out_0 = tdf11_accum_1_U0_ap_done;

assign ap_channel_done_ifmap_vec = tdf11_readInputs75_U0_ap_done;

assign ap_channel_done_intermediate_fmaps_0 = tdf11_adjust_U0_ap_done;

assign ap_channel_done_l2_products = tdf11_l2_multiply72_U0_ap_done;

assign ap_channel_done_products_0 = tdf11_dot_product_U0_ap_done;

assign ap_channel_done_sums_0 = Block_entry_proc_proc441_U0_ap_done;

assign ap_channel_done_tmp_channel = tdf11_accum_2_U0_ap_done;

assign ap_channel_done_weight_vecs_0 = tdf11_readFilters74_U0_ap_done;

assign ap_done = tdf11_l2_writeOutputs_171_U0_ap_done;

assign ap_idle = (tdf11_readInputs75_U0_ap_idle & tdf11_readFilters74_U0_ap_idle & tdf11_l2_writeOutputs_171_U0_ap_idle & tdf11_l2_multiply72_U0_ap_idle & tdf11_get_next_ijk_U0_ap_idle & tdf11_dot_product_U0_ap_idle & tdf11_adjust_U0_ap_idle & tdf11_accum_2_U0_ap_idle & tdf11_accum_1_U0_ap_idle & (intermediate_fmaps_0_empty_n ^ 1'b1) & (sums_0_empty_n ^ 1'b1) & (tmp_channel_empty_n ^ 1'b1) & (l2_products_t_empty_n ^ 1'b1) & (products_0_t_empty_n ^ 1'b1) & (weight_vecs_0_t_empty_n ^ 1'b1) & (ifmap_vec_t_empty_n ^ 1'b1) & (1'b1 ^ accum1_out_0_t_empty_n) & Block_entry_proc_proc441_U0_ap_idle);

assign ap_ready = ap_sync_ready;

assign ap_sync_continue = ap_continue;

assign ap_sync_done = tdf11_l2_writeOutputs_171_U0_ap_done;

assign ap_sync_ready = (ap_sync_tdf11_readInputs75_U0_ap_ready & ap_sync_tdf11_get_next_ijk_U0_ap_ready);

assign ap_sync_tdf11_get_next_ijk_U0_ap_ready = (tdf11_get_next_ijk_U0_ap_ready | ap_sync_reg_tdf11_get_next_ijk_U0_ap_ready);

assign ap_sync_tdf11_readInputs75_U0_ap_ready = (tdf11_readInputs75_U0_ap_ready | ap_sync_reg_tdf11_readInputs75_U0_ap_ready);

assign in_data_address0 = tdf11_readInputs75_U0_in_data_address0;

assign in_data_address1 = 12'd0;

assign in_data_ce0 = tdf11_readInputs75_U0_in_data_ce0;

assign in_data_ce1 = 1'b0;

assign in_data_d0 = 64'd0;

assign in_data_d1 = 64'd0;

assign in_data_read = tdf11_readInputs75_U0_in_data_write;

assign in_data_we0 = 1'b0;

assign in_data_we1 = 1'b0;

assign l1_adjustments_address0 = tdf11_adjust_U0_adjustments_address0;

assign l1_adjustments_address1 = 9'd0;

assign l1_adjustments_ce0 = tdf11_adjust_U0_adjustments_ce0;

assign l1_adjustments_ce1 = 1'b0;

assign l1_adjustments_d0 = 48'd0;

assign l1_adjustments_d1 = 48'd0;

assign l1_adjustments_we0 = 1'b0;

assign l1_adjustments_we1 = 1'b0;

assign l1_filter_data_address0 = tdf11_readFilters74_U0_filter_data_address0;

assign l1_filter_data_address1 = 17'd0;

assign l1_filter_data_ce0 = tdf11_readFilters74_U0_filter_data_ce0;

assign l1_filter_data_ce1 = 1'b0;

assign l1_filter_data_d0 = 64'd0;

assign l1_filter_data_d1 = 64'd0;

assign l1_filter_data_we0 = 1'b0;

assign l1_filter_data_we1 = 1'b0;

assign l2_adjustments_address0 = tdf11_l2_writeOutputs_171_U0_l2_adjustments_address0;

assign l2_adjustments_address1 = 7'd0;

assign l2_adjustments_ce0 = tdf11_l2_writeOutputs_171_U0_l2_adjustments_ce0;

assign l2_adjustments_ce1 = 1'b0;

assign l2_adjustments_d0 = 48'd0;

assign l2_adjustments_d1 = 48'd0;

assign l2_adjustments_we0 = 1'b0;

assign l2_adjustments_we1 = 1'b0;

assign l2_filter_data_address0 = tdf11_l2_multiply72_U0_l2_filter_data_address0;

assign l2_filter_data_address1 = 16'd0;

assign l2_filter_data_ce0 = tdf11_l2_multiply72_U0_l2_filter_data_ce0;

assign l2_filter_data_ce1 = 1'b0;

assign l2_filter_data_d0 = 16'd0;

assign l2_filter_data_d1 = 16'd0;

assign l2_filter_data_we0 = 1'b0;

assign l2_filter_data_we1 = 1'b0;

assign out_data_address0 = 13'd0;

assign out_data_address1 = tdf11_l2_writeOutputs_171_U0_out_data_address1;

assign out_data_ce0 = 1'b0;

assign out_data_ce1 = tdf11_l2_writeOutputs_171_U0_out_data_ce1;

assign out_data_d0 = 64'd0;

assign out_data_d1 = tdf11_l2_writeOutputs_171_U0_out_data_d1;

assign out_data_we0 = 1'b0;

assign out_data_we1 = tdf11_l2_writeOutputs_171_U0_out_data_we1;

assign out_data_write = tdf11_l2_writeOutputs_171_U0_out_data_write;

assign products_0_t_d1 = 16'd0;

assign products_0_t_we1 = 1'b0;

assign start_for_tdf11_readFilters74_U0_din = 1'b1;

assign tdf11_accum_1_U0_accum_out_full_n = accum1_out_0_i_full_n;

assign tdf11_accum_1_U0_ap_continue = accum1_out_0_i_full_n;

assign tdf11_accum_1_U0_ap_start = products_0_t_empty_n;

assign tdf11_accum_1_U0_start_full_n = 1'b1;

assign tdf11_accum_1_U0_start_write = 1'b0;

assign tdf11_accum_2_U0_ap_continue = tmp_channel_full_n;

assign tdf11_accum_2_U0_ap_start = accum1_out_0_t_empty_n;

assign tdf11_accum_2_U0_start_full_n = 1'b1;

assign tdf11_accum_2_U0_start_write = 1'b0;

assign tdf11_adjust_U0_ap_continue = intermediate_fmaps_0_full_n;

assign tdf11_adjust_U0_ap_start = sums_0_empty_n;

assign tdf11_adjust_U0_start_full_n = 1'b1;

assign tdf11_adjust_U0_start_write = 1'b0;

assign tdf11_dot_product_U0_ap_continue = products_0_i_full_n;

assign tdf11_dot_product_U0_ap_start = (weight_vecs_0_t_empty_n & ifmap_vec_t_empty_n);

assign tdf11_dot_product_U0_products_0_full_n = products_0_i_full_n;

assign tdf11_dot_product_U0_start_full_n = 1'b1;

assign tdf11_dot_product_U0_start_write = 1'b0;

assign tdf11_get_next_ijk_U0_ap_continue = 1'b1;

assign tdf11_get_next_ijk_U0_ap_start = ((ap_sync_reg_tdf11_get_next_ijk_U0_ap_ready ^ 1'b1) & ap_start);

assign tdf11_l2_multiply72_U0_ap_continue = l2_products_i_full_n;

assign tdf11_l2_multiply72_U0_ap_start = intermediate_fmaps_0_empty_n;

assign tdf11_l2_multiply72_U0_l2_products_full_n = l2_products_i_full_n;

assign tdf11_l2_multiply72_U0_start_full_n = 1'b1;

assign tdf11_l2_multiply72_U0_start_write = 1'b0;

assign tdf11_l2_writeOutputs_171_U0_ap_continue = ap_continue;

assign tdf11_l2_writeOutputs_171_U0_ap_start = l2_products_t_empty_n;

assign tdf11_l2_writeOutputs_171_U0_out_data_full_n = out_data_full_n;

assign tdf11_l2_writeOutputs_171_U0_out_data_write = 1'b0;

assign tdf11_l2_writeOutputs_171_U0_start_full_n = 1'b1;

assign tdf11_l2_writeOutputs_171_U0_start_write = 1'b0;

assign tdf11_readFilters74_U0_ap_continue = weight_vecs_0_i_full_n;

assign tdf11_readFilters74_U0_ap_start = start_for_tdf11_readFilters74_U0_empty_n;

assign tdf11_readFilters74_U0_start_full_n = 1'b1;

assign tdf11_readFilters74_U0_start_write = 1'b0;

assign tdf11_readFilters74_U0_weight_vecs_0_full_n = weight_vecs_0_i_full_n;

assign tdf11_readInputs75_U0_ap_continue = ifmap_vec_i_full_n;

assign tdf11_readInputs75_U0_ap_start = ((ap_sync_reg_tdf11_readInputs75_U0_ap_ready ^ 1'b1) & ap_start);

assign tdf11_readInputs75_U0_ifmap_vec_full_n = ifmap_vec_i_full_n;

assign tdf11_readInputs75_U0_in_data_full_n = in_data_empty_n;

assign tdf11_readInputs75_U0_in_data_write = 1'b0;

assign tdf11_readInputs75_U0_start_full_n = 1'b1;

assign tdf11_readInputs75_U0_start_write = 1'b0;

assign write4_c_din = tdf11_get_next_ijk_U0_write_r_din;

endmodule //td_fused_top_dataflow_in_loop_TOP_LOOP38270
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP38364_accum1_out_0_memcore_ram (addr0, ce0, d0, we0, q0, addr1, ce1, d1, we1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 3;
parameter MEM_SIZE = 8;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
input clk;

reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];




always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1) 
            ram[addr1] <= d1; 
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP38364_accum1_out_0_memcore(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    q0,
    address1,
    ce1,
    we1,
    d1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd8;
parameter AddressWidth = 32'd3;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;



td_fused_top_dataflow_in_loop_TOP_LOOP38364_accum1_out_0_memcore_ram td_fused_top_dataflow_in_loop_TOP_LOOP38364_accum1_out_0_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_dataflow_in_loop_TOP_LOOP38364_accum1_out_0
#(parameter
    DataWidth    = 16,
    AddressRange = 32,
    AddressWidth = 3,
    BufferCount  = 2,
    MemLatency   = 1,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire                    i_we0,
    input  wire [AddressWidth-1:0] i_address0,
    input  wire [DataWidth-1:0]    i_d0,
    output wire [DataWidth-1:0]    i_q0,
    input  wire                    i_ce1,
    input  wire                    i_we1,
    input  wire [AddressWidth-1:0] i_address1,
    input  wire [DataWidth-1:0]    i_d1,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire                    t_we0,
    input  wire [AddressWidth-1:0] t_address0,
    input  wire [DataWidth-1:0]    t_d0,
    output wire [DataWidth-1:0]    t_q0,
    input  wire                    t_ce1,
    input  wire                    t_we1,
    input  wire [AddressWidth-1:0] t_address1,
    input  wire [DataWidth-1:0]    t_d1
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth-1:0]   prev_iptr    = 1'b0; // previous initiator index
reg  [IndexWidth-1:0]   prev_tptr    = 1'b0; // previous target index
reg  [DataWidth-1:0]    reg_q0      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid0    = 1'b0; // buffer has valid data
reg  [DataWidth-1:0]    reg_q1      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid1    = 1'b0; // buffer has valid data
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
// buffer signals
wire [BufferCount-1:0] buf_ce0;
wire [BufferCount-1:0] buf_we0;
wire [AddressWidth-1:0] buf_a0_0, buf_a0_1;
wire [DataWidth-1:0] buf_d0_0, buf_d0_1;
wire [DataWidth-1:0] buf_q0_0, buf_q0_1;
wire [BufferCount-1:0] buf_ce1;
wire [BufferCount-1:0] buf_we1;
wire [AddressWidth-1:0] buf_a1_0, buf_a1_1;
wire [DataWidth-1:0] buf_d1_0, buf_d1_1;
//------------------------Instantiation------------------
//genvar i;
        td_fused_top_dataflow_in_loop_TOP_LOOP38364_accum1_out_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP38364_accum1_out_0_memcore_U_0 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_0 ),
            .ce0      ( buf_ce0[ 0 ] ),
            .we0      ( buf_we0[ 0 ] ),
            .d0       ( buf_d0_0 ),
            .q0       ( buf_q0_0 ),
            .address1 ( buf_a1_0 ),
            .ce1      ( buf_ce1[ 0 ] ),
            .we1      ( buf_we1[ 0 ] ),
            .d1       ( buf_d1_0 )
        );
        td_fused_top_dataflow_in_loop_TOP_LOOP38364_accum1_out_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP38364_accum1_out_0_memcore_U_1 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_1 ),
            .ce0      ( buf_ce0[ 1 ] ),
            .we0      ( buf_we0[ 1 ] ),
            .d0       ( buf_d0_1 ),
            .q0       ( buf_q0_1 ),
            .address1 ( buf_a1_1 ),
            .ce1      ( buf_ce1[ 1 ] ),
            .we1      ( buf_we1[ 1 ] ),
            .d1       ( buf_d1_1 )
        );

//++++++++++++++++++++++++buffer signals+++++++++++++++++
        assign buf_ce0[ 0 ] = (tptr ==  0  && empty_n) ? t_ce0
                             : (iptr ==  0 ) ? i_ce0 : 1'b0;
        assign buf_a0_0  = (tptr ==  0  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 0 ] = (tptr ==  0  && empty_n)  ? t_we0
                             : (iptr ==  0 ) ? i_we0 : 1'b0;
        assign buf_d0_0  = (tptr ==  0  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 0 ] = (tptr ==  0  && empty_n) ? t_ce1
                             : (iptr ==  0 ) ? i_ce1 : 1'b0;
        assign buf_a1_0  = (tptr ==  0  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 0 ] = (tptr ==  0  && empty_n)  ? t_we1
                             : (iptr ==  0 ) ? i_we1 : 1'b0;
        assign buf_d1_0  = (tptr ==  0  && empty_n) ? t_d1       : i_d1;
        assign buf_ce0[ 1 ] = (tptr ==  1  && empty_n) ? t_ce0
                             : (iptr ==  1 ) ? i_ce0 : 1'b0;
        assign buf_a0_1  = (tptr ==  1  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 1 ] = (tptr ==  1  && empty_n)  ? t_we0
                             : (iptr ==  1 ) ? i_we0 : 1'b0;
        assign buf_d0_1  = (tptr ==  1  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 1 ] = (tptr ==  1  && empty_n) ? t_ce1
                             : (iptr ==  1 ) ? i_ce1 : 1'b0;
        assign buf_a1_1  = (tptr ==  1  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 1 ] = (tptr ==  1  && empty_n)  ? t_we1
                             : (iptr ==  1 ) ? i_we1 : 1'b0;
        assign buf_d1_1  = (tptr ==  1  && empty_n) ? t_d1       : i_d1;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//------------------------Body---------------------------
assign i_q0      = (prev_iptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign t_q0      = reg_valid0 ? reg_q0 : (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// prev_iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_iptr <= 1'b0;
    else begin
        prev_iptr <= iptr;
    end
end

// prev_tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_tptr <= 1'b0;
    else begin
        prev_tptr <= tptr;
    end
end

// reg_q0 and reg_valid0
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q0     <= 1'b0;
        reg_valid0 <= 1'b0;
    end else if (!t_ce0 && !reg_valid0) begin
        reg_q0     <= (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
        reg_valid0 <= 1'b1;
    end else if (t_ce0) begin
        reg_valid0 <= 1'b0;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP38364_ifmap_vec_memcore_ram (addr0, ce0, d0, we0, q0, addr1, ce1, d1, we1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 10;
parameter MEM_SIZE = 576;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
input clk;

reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];




always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1) 
            ram[addr1] <= d1; 
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP38364_ifmap_vec_memcore(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    q0,
    address1,
    ce1,
    we1,
    d1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd576;
parameter AddressWidth = 32'd10;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;



td_fused_top_dataflow_in_loop_TOP_LOOP38364_ifmap_vec_memcore_ram td_fused_top_dataflow_in_loop_TOP_LOOP38364_ifmap_vec_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_dataflow_in_loop_TOP_LOOP38364_ifmap_vec
#(parameter
    DataWidth    = 16,
    AddressRange = 32,
    AddressWidth = 10,
    BufferCount  = 2,
    MemLatency   = 1,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire                    i_we0,
    input  wire [AddressWidth-1:0] i_address0,
    input  wire [DataWidth-1:0]    i_d0,
    output wire [DataWidth-1:0]    i_q0,
    input  wire                    i_ce1,
    input  wire                    i_we1,
    input  wire [AddressWidth-1:0] i_address1,
    input  wire [DataWidth-1:0]    i_d1,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire                    t_we0,
    input  wire [AddressWidth-1:0] t_address0,
    input  wire [DataWidth-1:0]    t_d0,
    output wire [DataWidth-1:0]    t_q0,
    input  wire                    t_ce1,
    input  wire                    t_we1,
    input  wire [AddressWidth-1:0] t_address1,
    input  wire [DataWidth-1:0]    t_d1
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth-1:0]   prev_iptr    = 1'b0; // previous initiator index
reg  [IndexWidth-1:0]   prev_tptr    = 1'b0; // previous target index
reg  [DataWidth-1:0]    reg_q0      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid0    = 1'b0; // buffer has valid data
reg  [DataWidth-1:0]    reg_q1      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid1    = 1'b0; // buffer has valid data
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
// buffer signals
wire [BufferCount-1:0] buf_ce0;
wire [BufferCount-1:0] buf_we0;
wire [AddressWidth-1:0] buf_a0_0, buf_a0_1;
wire [DataWidth-1:0] buf_d0_0, buf_d0_1;
wire [DataWidth-1:0] buf_q0_0, buf_q0_1;
wire [BufferCount-1:0] buf_ce1;
wire [BufferCount-1:0] buf_we1;
wire [AddressWidth-1:0] buf_a1_0, buf_a1_1;
wire [DataWidth-1:0] buf_d1_0, buf_d1_1;
//------------------------Instantiation------------------
//genvar i;
        td_fused_top_dataflow_in_loop_TOP_LOOP38364_ifmap_vec_memcore td_fused_top_dataflow_in_loop_TOP_LOOP38364_ifmap_vec_memcore_U_0 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_0 ),
            .ce0      ( buf_ce0[ 0 ] ),
            .we0      ( buf_we0[ 0 ] ),
            .d0       ( buf_d0_0 ),
            .q0       ( buf_q0_0 ),
            .address1 ( buf_a1_0 ),
            .ce1      ( buf_ce1[ 0 ] ),
            .we1      ( buf_we1[ 0 ] ),
            .d1       ( buf_d1_0 )
        );
        td_fused_top_dataflow_in_loop_TOP_LOOP38364_ifmap_vec_memcore td_fused_top_dataflow_in_loop_TOP_LOOP38364_ifmap_vec_memcore_U_1 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_1 ),
            .ce0      ( buf_ce0[ 1 ] ),
            .we0      ( buf_we0[ 1 ] ),
            .d0       ( buf_d0_1 ),
            .q0       ( buf_q0_1 ),
            .address1 ( buf_a1_1 ),
            .ce1      ( buf_ce1[ 1 ] ),
            .we1      ( buf_we1[ 1 ] ),
            .d1       ( buf_d1_1 )
        );

//++++++++++++++++++++++++buffer signals+++++++++++++++++
        assign buf_ce0[ 0 ] = (tptr ==  0  && empty_n) ? t_ce0
                             : (iptr ==  0 ) ? i_ce0 : 1'b0;
        assign buf_a0_0  = (tptr ==  0  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 0 ] = (tptr ==  0  && empty_n)  ? t_we0
                             : (iptr ==  0 ) ? i_we0 : 1'b0;
        assign buf_d0_0  = (tptr ==  0  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 0 ] = (tptr ==  0  && empty_n) ? t_ce1
                             : (iptr ==  0 ) ? i_ce1 : 1'b0;
        assign buf_a1_0  = (tptr ==  0  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 0 ] = (tptr ==  0  && empty_n)  ? t_we1
                             : (iptr ==  0 ) ? i_we1 : 1'b0;
        assign buf_d1_0  = (tptr ==  0  && empty_n) ? t_d1       : i_d1;
        assign buf_ce0[ 1 ] = (tptr ==  1  && empty_n) ? t_ce0
                             : (iptr ==  1 ) ? i_ce0 : 1'b0;
        assign buf_a0_1  = (tptr ==  1  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 1 ] = (tptr ==  1  && empty_n)  ? t_we0
                             : (iptr ==  1 ) ? i_we0 : 1'b0;
        assign buf_d0_1  = (tptr ==  1  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 1 ] = (tptr ==  1  && empty_n) ? t_ce1
                             : (iptr ==  1 ) ? i_ce1 : 1'b0;
        assign buf_a1_1  = (tptr ==  1  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 1 ] = (tptr ==  1  && empty_n)  ? t_we1
                             : (iptr ==  1 ) ? i_we1 : 1'b0;
        assign buf_d1_1  = (tptr ==  1  && empty_n) ? t_d1       : i_d1;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//------------------------Body---------------------------
assign i_q0      = (prev_iptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign t_q0      = reg_valid0 ? reg_q0 : (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// prev_iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_iptr <= 1'b0;
    else begin
        prev_iptr <= iptr;
    end
end

// prev_tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_tptr <= 1'b0;
    else begin
        prev_tptr <= tptr;
    end
end

// reg_q0 and reg_valid0
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q0     <= 1'b0;
        reg_valid0 <= 1'b0;
    end else if (!t_ce0 && !reg_valid0) begin
        reg_q0     <= (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
        reg_valid0 <= 1'b1;
    end else if (t_ce0) begin
        reg_valid0 <= 1'b0;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP38364_l2_products_memcore_ram (addr0, ce0, d0, we0, q0, addr1, ce1, d1, we1, q1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
output reg[DWIDTH-1:0] q1;
input clk;

 reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];




always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1) 
            ram[addr1] <= d1; 
        q1 <= ram[addr1];
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP38364_l2_products_memcore(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    q0,
    address1,
    ce1,
    we1,
    d1,
    q1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;
output[DataWidth - 1:0] q1;



td_fused_top_dataflow_in_loop_TOP_LOOP38364_l2_products_memcore_ram td_fused_top_dataflow_in_loop_TOP_LOOP38364_l2_products_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 ),
    .q1( q1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_dataflow_in_loop_TOP_LOOP38364_l2_products
#(parameter
    DataWidth    = 16,
    AddressRange = 32,
    AddressWidth = 6,
    BufferCount  = 2,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire                    i_we0,
    input  wire [AddressWidth-1:0] i_address0,
    input  wire [DataWidth-1:0]    i_d0,
    output wire [DataWidth-1:0]    i_q0,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire                    t_we0,
    input  wire [AddressWidth-1:0] t_address0,
    input  wire [DataWidth-1:0]    t_d0,
    output wire [DataWidth-1:0]    t_q0
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
wire [AddressWidth+IndexWidth-1:0]   memcore_iaddr;
wire [AddressWidth+IndexWidth-1:0]   memcore_taddr;

//------------------------Instantiation------------------
assign memcore_iaddr = {i_address0, iptr};
assign memcore_taddr = {t_address0, tptr};
td_fused_top_dataflow_in_loop_TOP_LOOP38364_l2_products_memcore td_fused_top_dataflow_in_loop_TOP_LOOP38364_l2_products_memcore_U (
    .reset    ( reset ),
    .clk      ( clk ),
    .address0 ( memcore_iaddr ),
    .ce0      ( i_ce0 ),
    .we0      ( i_we0),
    .d0       ( i_d0 ),
    .q0       ( i_q0 ),
    .address1 ( memcore_taddr ),
    .ce1      ( t_ce0 ),
    .we1      ( t_we0),
    .d1       ( t_d0 ),
    .q1       ( t_q0 )

);

//------------------------Body---------------------------

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP38364_products_0_memcore_ram (addr0, ce0, d0, we0, q0, addr1, ce1, q1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 10;
parameter MEM_SIZE = 576;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
output reg[DWIDTH-1:0] q1;
input clk;

reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];




always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        q1 <= ram[addr1];
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP38364_products_0_memcore(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    q0,
    address1,
    ce1,
    q1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd576;
parameter AddressWidth = 32'd10;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
output[DataWidth - 1:0] q1;



td_fused_top_dataflow_in_loop_TOP_LOOP38364_products_0_memcore_ram td_fused_top_dataflow_in_loop_TOP_LOOP38364_products_0_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .q1( q1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_dataflow_in_loop_TOP_LOOP38364_products_0
#(parameter
    DataWidth    = 16,
    AddressRange = 32,
    AddressWidth = 10,
    BufferCount  = 2,
    MemLatency   = 1,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire                    i_we0,
    input  wire [AddressWidth-1:0] i_address0,
    input  wire [DataWidth-1:0]    i_d0,
    output wire [DataWidth-1:0]    i_q0,
    input  wire                    i_ce1,
    input  wire [AddressWidth-1:0] i_address1,
    output wire [DataWidth-1:0]    i_q1,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire                    t_we0,
    input  wire [AddressWidth-1:0] t_address0,
    input  wire [DataWidth-1:0]    t_d0,
    output wire [DataWidth-1:0]    t_q0,
    input  wire                    t_ce1,
    input  wire [AddressWidth-1:0] t_address1,
    output wire [DataWidth-1:0]    t_q1
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth-1:0]   prev_iptr    = 1'b0; // previous initiator index
reg  [IndexWidth-1:0]   prev_tptr    = 1'b0; // previous target index
reg  [DataWidth-1:0]    reg_q0      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid0    = 1'b0; // buffer has valid data
reg  [DataWidth-1:0]    reg_q1      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid1    = 1'b0; // buffer has valid data
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
// buffer signals
wire [BufferCount-1:0] buf_ce0;
wire [BufferCount-1:0] buf_we0;
wire [AddressWidth-1:0] buf_a0_0, buf_a0_1;
wire [DataWidth-1:0] buf_d0_0, buf_d0_1;
wire [DataWidth-1:0] buf_q0_0, buf_q0_1;
wire [BufferCount-1:0] buf_ce1;
wire [AddressWidth-1:0] buf_a1_0, buf_a1_1;
wire [DataWidth-1:0] buf_q1_0, buf_q1_1;
//------------------------Instantiation------------------
//genvar i;
        td_fused_top_dataflow_in_loop_TOP_LOOP38364_products_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP38364_products_0_memcore_U_0 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_0 ),
            .ce0      ( buf_ce0[ 0 ] ),
            .we0      ( buf_we0[ 0 ] ),
            .d0       ( buf_d0_0 ),
            .q0       ( buf_q0_0 ),
            .address1 ( buf_a1_0 ),
            .ce1      ( buf_ce1[ 0 ] ),
            .q1       ( buf_q1_0 )
        );
        td_fused_top_dataflow_in_loop_TOP_LOOP38364_products_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP38364_products_0_memcore_U_1 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_1 ),
            .ce0      ( buf_ce0[ 1 ] ),
            .we0      ( buf_we0[ 1 ] ),
            .d0       ( buf_d0_1 ),
            .q0       ( buf_q0_1 ),
            .address1 ( buf_a1_1 ),
            .ce1      ( buf_ce1[ 1 ] ),
            .q1       ( buf_q1_1 )
        );

//++++++++++++++++++++++++buffer signals+++++++++++++++++
        assign buf_ce0[ 0 ] = (tptr ==  0  && empty_n) ? t_ce0
                             : (iptr ==  0 ) ? i_ce0 : 1'b0;
        assign buf_a0_0  = (tptr ==  0  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 0 ] = (tptr ==  0  && empty_n)  ? t_we0
                             : (iptr ==  0 ) ? i_we0 : 1'b0;
        assign buf_d0_0  = (tptr ==  0  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 0 ] = (tptr ==  0  && empty_n) ? t_ce1
                             : (iptr ==  0 ) ? i_ce1 : 1'b0;
        assign buf_a1_0  = (tptr ==  0  && empty_n) ?  t_address1 : i_address1;
        assign buf_ce0[ 1 ] = (tptr ==  1  && empty_n) ? t_ce0
                             : (iptr ==  1 ) ? i_ce0 : 1'b0;
        assign buf_a0_1  = (tptr ==  1  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 1 ] = (tptr ==  1  && empty_n)  ? t_we0
                             : (iptr ==  1 ) ? i_we0 : 1'b0;
        assign buf_d0_1  = (tptr ==  1  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 1 ] = (tptr ==  1  && empty_n) ? t_ce1
                             : (iptr ==  1 ) ? i_ce1 : 1'b0;
        assign buf_a1_1  = (tptr ==  1  && empty_n) ?  t_address1 : i_address1;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//------------------------Body---------------------------
assign i_q0      = (prev_iptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign t_q0      = reg_valid0 ? reg_q0 : (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign i_q1      = (prev_iptr == 1'b1 ? buf_q1_1 : buf_q1_0);
assign t_q1      = reg_valid1 ? reg_q1 : (prev_tptr == 1'b1 ? buf_q1_1 : buf_q1_0);

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// prev_iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_iptr <= 1'b0;
    else begin
        prev_iptr <= iptr;
    end
end

// prev_tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_tptr <= 1'b0;
    else begin
        prev_tptr <= tptr;
    end
end

// reg_q0 and reg_valid0
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q0     <= 1'b0;
        reg_valid0 <= 1'b0;
    end else if (!t_ce0 && !reg_valid0) begin
        reg_q0     <= (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
        reg_valid0 <= 1'b1;
    end else if (t_ce0) begin
        reg_valid0 <= 1'b0;
    end
end

// reg_q1 and reg_valid1
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q1     <= 1'b0;
        reg_valid1 <= 1'b0;
    end else if (!t_ce1 && !reg_valid1) begin
        reg_q1     <= (prev_tptr == 1'b1 ? buf_q1_1 : buf_q1_0);
        reg_valid1 <= 1'b1;
    end else if (t_ce1) begin
        reg_valid1 <= 1'b0;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_dataflow_in_loop_TOP_LOOP38364 (
        ap_clk,
        ap_rst,
        in_data_address0,
        in_data_ce0,
        in_data_d0,
        in_data_q0,
        in_data_we0,
        in_data_address1,
        in_data_ce1,
        in_data_d1,
        in_data_q1,
        in_data_we1,
        l1_filter_data_address0,
        l1_filter_data_ce0,
        l1_filter_data_d0,
        l1_filter_data_q0,
        l1_filter_data_we0,
        l1_filter_data_address1,
        l1_filter_data_ce1,
        l1_filter_data_d1,
        l1_filter_data_q1,
        l1_filter_data_we1,
        l1_adjustments_address0,
        l1_adjustments_ce0,
        l1_adjustments_d0,
        l1_adjustments_q0,
        l1_adjustments_we0,
        l1_adjustments_address1,
        l1_adjustments_ce1,
        l1_adjustments_d1,
        l1_adjustments_q1,
        l1_adjustments_we1,
        l2_filter_data_address0,
        l2_filter_data_ce0,
        l2_filter_data_d0,
        l2_filter_data_q0,
        l2_filter_data_we0,
        l2_filter_data_address1,
        l2_filter_data_ce1,
        l2_filter_data_d1,
        l2_filter_data_q1,
        l2_filter_data_we1,
        out_data_address0,
        out_data_ce0,
        out_data_d0,
        out_data_q0,
        out_data_we0,
        out_data_address1,
        out_data_ce1,
        out_data_d1,
        out_data_q1,
        out_data_we1,
        l2_adjustments_address0,
        l2_adjustments_ce0,
        l2_adjustments_d0,
        l2_adjustments_q0,
        l2_adjustments_we0,
        l2_adjustments_address1,
        l2_adjustments_ce1,
        l2_adjustments_d1,
        l2_adjustments_q1,
        l2_adjustments_we1,
        ap_start,
        in_data_empty_n,
        in_data_read,
        out_data_full_n,
        out_data_write,
        ap_done,
        ap_ready,
        ap_idle,
        ap_continue
);


input   ap_clk;
input   ap_rst;
output  [11:0] in_data_address0;
output   in_data_ce0;
output  [63:0] in_data_d0;
input  [63:0] in_data_q0;
output   in_data_we0;
output  [11:0] in_data_address1;
output   in_data_ce1;
output  [63:0] in_data_d1;
input  [63:0] in_data_q1;
output   in_data_we1;
output  [16:0] l1_filter_data_address0;
output   l1_filter_data_ce0;
output  [63:0] l1_filter_data_d0;
input  [63:0] l1_filter_data_q0;
output   l1_filter_data_we0;
output  [16:0] l1_filter_data_address1;
output   l1_filter_data_ce1;
output  [63:0] l1_filter_data_d1;
input  [63:0] l1_filter_data_q1;
output   l1_filter_data_we1;
output  [8:0] l1_adjustments_address0;
output   l1_adjustments_ce0;
output  [47:0] l1_adjustments_d0;
input  [47:0] l1_adjustments_q0;
output   l1_adjustments_we0;
output  [8:0] l1_adjustments_address1;
output   l1_adjustments_ce1;
output  [47:0] l1_adjustments_d1;
input  [47:0] l1_adjustments_q1;
output   l1_adjustments_we1;
output  [14:0] l2_filter_data_address0;
output   l2_filter_data_ce0;
output  [15:0] l2_filter_data_d0;
input  [15:0] l2_filter_data_q0;
output   l2_filter_data_we0;
output  [14:0] l2_filter_data_address1;
output   l2_filter_data_ce1;
output  [15:0] l2_filter_data_d1;
input  [15:0] l2_filter_data_q1;
output   l2_filter_data_we1;
output  [11:0] out_data_address0;
output   out_data_ce0;
output  [63:0] out_data_d0;
input  [63:0] out_data_q0;
output   out_data_we0;
output  [11:0] out_data_address1;
output   out_data_ce1;
output  [63:0] out_data_d1;
input  [63:0] out_data_q1;
output   out_data_we1;
output  [5:0] l2_adjustments_address0;
output   l2_adjustments_ce0;
output  [47:0] l2_adjustments_d0;
input  [47:0] l2_adjustments_q0;
output   l2_adjustments_we0;
output  [5:0] l2_adjustments_address1;
output   l2_adjustments_ce1;
output  [47:0] l2_adjustments_d1;
input  [47:0] l2_adjustments_q1;
output   l2_adjustments_we1;
input   ap_start;
input   in_data_empty_n;
output   in_data_read;
input   out_data_full_n;
output   out_data_write;
output   ap_done;
output   ap_ready;
output   ap_idle;
input   ap_continue;

wire   [15:0] ifmap_vec_i_q0;
wire   [15:0] ifmap_vec_t_q0;
wire   [15:0] weight_vecs_0_i_q0;
wire   [15:0] weight_vecs_0_t_q0;
wire   [15:0] products_0_i_q0;
wire   [15:0] products_0_i_q1;
wire   [15:0] products_0_t_q0;
wire   [15:0] products_0_t_q1;
wire   [15:0] accum1_out_0_i_q0;
wire   [15:0] accum1_out_0_t_q0;
wire   [15:0] l2_products_i_q0;
wire   [15:0] l2_products_t_q0;
wire    tdf10_get_next_ijk_U0_ap_start;
wire    tdf10_get_next_ijk_U0_ap_done;
wire    tdf10_get_next_ijk_U0_ap_continue;
wire    tdf10_get_next_ijk_U0_ap_idle;
wire    tdf10_get_next_ijk_U0_ap_ready;
wire    tdf10_get_next_ijk_U0_start_out;
wire    tdf10_get_next_ijk_U0_start_write;
wire   [15:0] tdf10_get_next_ijk_U0_indices_0_din;
wire    tdf10_get_next_ijk_U0_indices_0_write;
wire   [15:0] tdf10_get_next_ijk_U0_indices_1_din;
wire    tdf10_get_next_ijk_U0_indices_1_write;
wire   [8:0] tdf10_get_next_ijk_U0_indices_2_out_din;
wire    tdf10_get_next_ijk_U0_indices_2_out_write;
wire   [14:0] tdf10_get_next_ijk_U0_indices_2_out1_din;
wire    tdf10_get_next_ijk_U0_indices_2_out1_write;
wire    tdf10_get_next_ijk_U0_write_r_din;
wire    tdf10_get_next_ijk_U0_write_r_write;
wire    tdf10_readInputs69_U0_ap_start;
wire    tdf10_readInputs69_U0_ap_done;
wire    tdf10_readInputs69_U0_ap_continue;
wire    tdf10_readInputs69_U0_ap_idle;
wire    tdf10_readInputs69_U0_ap_ready;
wire   [11:0] tdf10_readInputs69_U0_in_data_address0;
wire    tdf10_readInputs69_U0_in_data_ce0;
wire    tdf10_readInputs69_U0_indices_01_read;
wire    tdf10_readInputs69_U0_indices_12_read;
wire   [9:0] tdf10_readInputs69_U0_ifmap_vec_address0;
wire    tdf10_readInputs69_U0_ifmap_vec_ce0;
wire    tdf10_readInputs69_U0_ifmap_vec_we0;
wire   [15:0] tdf10_readInputs69_U0_ifmap_vec_d0;
wire   [9:0] tdf10_readInputs69_U0_ifmap_vec_address1;
wire    tdf10_readInputs69_U0_ifmap_vec_ce1;
wire    tdf10_readInputs69_U0_ifmap_vec_we1;
wire   [15:0] tdf10_readInputs69_U0_ifmap_vec_d1;
wire   [3:0] tdf10_readInputs69_U0_indices_01_out_din;
wire    tdf10_readInputs69_U0_indices_01_out_write;
wire   [7:0] tdf10_readInputs69_U0_indices_12_out_din;
wire    tdf10_readInputs69_U0_indices_12_out_write;
wire    tdf10_readInputs69_U0_in_data_full_n;
wire    tdf10_readInputs69_U0_in_data_write;
wire    ap_channel_done_ifmap_vec;
wire    tdf10_readInputs69_U0_ifmap_vec_full_n;
wire    tdf10_readFilters68_U0_ap_start;
wire    tdf10_readFilters68_U0_ap_done;
wire    tdf10_readFilters68_U0_ap_continue;
wire    tdf10_readFilters68_U0_ap_idle;
wire    tdf10_readFilters68_U0_ap_ready;
wire   [16:0] tdf10_readFilters68_U0_filter_data_address0;
wire    tdf10_readFilters68_U0_filter_data_ce0;
wire    tdf10_readFilters68_U0_indices_23_read;
wire   [9:0] tdf10_readFilters68_U0_weight_vecs_0_address0;
wire    tdf10_readFilters68_U0_weight_vecs_0_ce0;
wire    tdf10_readFilters68_U0_weight_vecs_0_we0;
wire   [15:0] tdf10_readFilters68_U0_weight_vecs_0_d0;
wire   [9:0] tdf10_readFilters68_U0_weight_vecs_0_address1;
wire    tdf10_readFilters68_U0_weight_vecs_0_ce1;
wire    tdf10_readFilters68_U0_weight_vecs_0_we1;
wire   [15:0] tdf10_readFilters68_U0_weight_vecs_0_d1;
wire    ap_channel_done_weight_vecs_0;
wire    tdf10_readFilters68_U0_weight_vecs_0_full_n;
wire    tdf10_dot_product_U0_ap_start;
wire    tdf10_dot_product_U0_ap_done;
wire    tdf10_dot_product_U0_ap_continue;
wire    tdf10_dot_product_U0_ap_idle;
wire    tdf10_dot_product_U0_ap_ready;
wire   [9:0] tdf10_dot_product_U0_ifmap_vec_address0;
wire    tdf10_dot_product_U0_ifmap_vec_ce0;
wire   [9:0] tdf10_dot_product_U0_weight_vecs_0_address0;
wire    tdf10_dot_product_U0_weight_vecs_0_ce0;
wire   [9:0] tdf10_dot_product_U0_products_0_address0;
wire    tdf10_dot_product_U0_products_0_ce0;
wire    tdf10_dot_product_U0_products_0_we0;
wire   [15:0] tdf10_dot_product_U0_products_0_d0;
wire    ap_channel_done_products_0;
wire    tdf10_dot_product_U0_products_0_full_n;
wire    tdf10_accum_1_U0_ap_start;
wire    tdf10_accum_1_U0_ap_done;
wire    tdf10_accum_1_U0_ap_continue;
wire    tdf10_accum_1_U0_ap_idle;
wire    tdf10_accum_1_U0_ap_ready;
wire   [9:0] tdf10_accum_1_U0_accum_in_0_address0;
wire    tdf10_accum_1_U0_accum_in_0_ce0;
wire   [9:0] tdf10_accum_1_U0_accum_in_0_address1;
wire    tdf10_accum_1_U0_accum_in_0_ce1;
wire   [2:0] tdf10_accum_1_U0_accum_out_address0;
wire    tdf10_accum_1_U0_accum_out_ce0;
wire    tdf10_accum_1_U0_accum_out_we0;
wire   [15:0] tdf10_accum_1_U0_accum_out_d0;
wire   [2:0] tdf10_accum_1_U0_accum_out_address1;
wire    tdf10_accum_1_U0_accum_out_ce1;
wire    tdf10_accum_1_U0_accum_out_we1;
wire   [15:0] tdf10_accum_1_U0_accum_out_d1;
wire    ap_channel_done_accum1_out_0;
wire    tdf10_accum_1_U0_accum_out_full_n;
wire    tdf10_accum_2_U0_ap_start;
wire    tdf10_accum_2_U0_ap_done;
wire    tdf10_accum_2_U0_ap_continue;
wire    tdf10_accum_2_U0_ap_idle;
wire    tdf10_accum_2_U0_ap_ready;
wire   [15:0] tdf10_accum_2_U0_accum_in_24;
wire    tdf10_accum_2_U0_accum_in_24_ap_vld;
wire   [2:0] tdf10_accum_2_U0_accum_in_address0;
wire    tdf10_accum_2_U0_accum_in_ce0;
wire    ap_channel_done_tmp_channel;
wire    tmp_channel_full_n;
wire    Block_entry_proc_proc435_U0_ap_start;
wire    Block_entry_proc_proc435_U0_ap_done;
wire    Block_entry_proc_proc435_U0_ap_continue;
wire    Block_entry_proc_proc435_U0_ap_idle;
wire    Block_entry_proc_proc435_U0_ap_ready;
wire   [15:0] Block_entry_proc_proc435_U0_ap_return;
wire    ap_channel_done_sums_0;
wire    sums_0_full_n;
wire    tdf10_adjust_U0_ap_start;
wire    tdf10_adjust_U0_ap_done;
wire    tdf10_adjust_U0_ap_continue;
wire    tdf10_adjust_U0_ap_idle;
wire    tdf10_adjust_U0_ap_ready;
wire   [8:0] tdf10_adjust_U0_adjustments_address0;
wire    tdf10_adjust_U0_adjustments_ce0;
wire    tdf10_adjust_U0_indices_23_read;
wire   [14:0] tdf10_adjust_U0_indices_23_out_din;
wire    tdf10_adjust_U0_indices_23_out_write;
wire   [15:0] tdf10_adjust_U0_ap_return;
wire    ap_channel_done_intermediate_fmaps_0;
wire    intermediate_fmaps_0_full_n;
wire    tdf10_l2_multiply66_U0_ap_start;
wire    tdf10_l2_multiply66_U0_ap_done;
wire    tdf10_l2_multiply66_U0_ap_continue;
wire    tdf10_l2_multiply66_U0_ap_idle;
wire    tdf10_l2_multiply66_U0_ap_ready;
wire   [14:0] tdf10_l2_multiply66_U0_l2_filter_data_address0;
wire    tdf10_l2_multiply66_U0_l2_filter_data_ce0;
wire   [5:0] tdf10_l2_multiply66_U0_l2_products_address0;
wire    tdf10_l2_multiply66_U0_l2_products_ce0;
wire    tdf10_l2_multiply66_U0_l2_products_we0;
wire   [15:0] tdf10_l2_multiply66_U0_l2_products_d0;
wire    tdf10_l2_multiply66_U0_indices_23_read;
wire    ap_channel_done_l2_products;
wire    tdf10_l2_multiply66_U0_l2_products_full_n;
wire    tdf10_l2_writeOutputs_165_U0_ap_start;
wire    tdf10_l2_writeOutputs_165_U0_ap_done;
wire    tdf10_l2_writeOutputs_165_U0_ap_continue;
wire    tdf10_l2_writeOutputs_165_U0_ap_idle;
wire    tdf10_l2_writeOutputs_165_U0_ap_ready;
wire    tdf10_l2_writeOutputs_165_U0_indices_01_read;
wire    tdf10_l2_writeOutputs_165_U0_indices_12_read;
wire    tdf10_l2_writeOutputs_165_U0_write4_read;
wire   [5:0] tdf10_l2_writeOutputs_165_U0_l2_partial_sums_address0;
wire    tdf10_l2_writeOutputs_165_U0_l2_partial_sums_ce0;
wire   [11:0] tdf10_l2_writeOutputs_165_U0_out_data_address1;
wire    tdf10_l2_writeOutputs_165_U0_out_data_ce1;
wire    tdf10_l2_writeOutputs_165_U0_out_data_we1;
wire   [63:0] tdf10_l2_writeOutputs_165_U0_out_data_d1;
wire   [5:0] tdf10_l2_writeOutputs_165_U0_l2_adjustments_address0;
wire    tdf10_l2_writeOutputs_165_U0_l2_adjustments_ce0;
wire    tdf10_l2_writeOutputs_165_U0_out_data_full_n;
wire    tdf10_l2_writeOutputs_165_U0_out_data_write;
wire    ap_sync_continue;
wire    ifmap_vec_i_full_n;
wire    ifmap_vec_t_empty_n;
wire    weight_vecs_0_i_full_n;
wire    weight_vecs_0_t_empty_n;
wire    products_0_i_full_n;
wire    products_0_t_empty_n;
wire   [15:0] products_0_t_d1;
wire    products_0_t_we1;
wire    accum1_out_0_i_full_n;
wire    accum1_out_0_t_empty_n;
wire    l2_products_i_full_n;
wire    l2_products_t_empty_n;
wire    indices_01_c_full_n;
wire   [15:0] indices_01_c_dout;
wire    indices_01_c_empty_n;
wire    indices_12_c_full_n;
wire   [15:0] indices_12_c_dout;
wire    indices_12_c_empty_n;
wire    indices_23_c_full_n;
wire   [8:0] indices_23_c_dout;
wire    indices_23_c_empty_n;
wire    indices_23_c1_full_n;
wire   [14:0] indices_23_c1_dout;
wire    indices_23_c1_empty_n;
wire   [0:0] write4_c_din;
wire    write4_c_full_n;
wire   [0:0] write4_c_dout;
wire    write4_c_empty_n;
wire    indices_01_c2_full_n;
wire   [3:0] indices_01_c2_dout;
wire    indices_01_c2_empty_n;
wire    indices_12_c3_full_n;
wire   [7:0] indices_12_c3_dout;
wire    indices_12_c3_empty_n;
wire   [15:0] tmp_channel_dout;
wire    tmp_channel_empty_n;
wire   [15:0] sums_0_dout;
wire    sums_0_empty_n;
wire    indices_23_c4_full_n;
wire   [14:0] indices_23_c4_dout;
wire    indices_23_c4_empty_n;
wire   [15:0] intermediate_fmaps_0_dout;
wire    intermediate_fmaps_0_empty_n;
wire    ap_sync_done;
wire    ap_sync_ready;
reg    ap_sync_reg_tdf10_get_next_ijk_U0_ap_ready;
wire    ap_sync_tdf10_get_next_ijk_U0_ap_ready;
reg    ap_sync_reg_tdf10_readInputs69_U0_ap_ready;
wire    ap_sync_tdf10_readInputs69_U0_ap_ready;
wire   [0:0] start_for_tdf10_readFilters68_U0_din;
wire    start_for_tdf10_readFilters68_U0_full_n;
wire   [0:0] start_for_tdf10_readFilters68_U0_dout;
wire    start_for_tdf10_readFilters68_U0_empty_n;
wire    tdf10_readInputs69_U0_start_full_n;
wire    tdf10_readInputs69_U0_start_write;
wire    tdf10_readFilters68_U0_start_full_n;
wire    tdf10_readFilters68_U0_start_write;
wire    tdf10_dot_product_U0_start_full_n;
wire    tdf10_dot_product_U0_start_write;
wire    tdf10_accum_1_U0_start_full_n;
wire    tdf10_accum_1_U0_start_write;
wire    tdf10_accum_2_U0_start_full_n;
wire    tdf10_accum_2_U0_start_write;
wire    Block_entry_proc_proc435_U0_start_full_n;
wire    Block_entry_proc_proc435_U0_start_write;
wire    tdf10_adjust_U0_start_full_n;
wire    tdf10_adjust_U0_start_write;
wire    tdf10_l2_multiply66_U0_start_full_n;
wire    tdf10_l2_multiply66_U0_start_write;
wire    tdf10_l2_writeOutputs_165_U0_start_full_n;
wire    tdf10_l2_writeOutputs_165_U0_start_write;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_sync_reg_tdf10_get_next_ijk_U0_ap_ready = 1'b0;
#0 ap_sync_reg_tdf10_readInputs69_U0_ap_ready = 1'b0;
end

td_fused_top_dataflow_in_loop_TOP_LOOP38364_ifmap_vec #(
    .DataWidth( 16 ),
    .AddressRange( 576 ),
    .AddressWidth( 10 ))
ifmap_vec_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf10_readInputs69_U0_ap_done),
    .i_full_n(ifmap_vec_i_full_n),
    .i_ce0(tdf10_readInputs69_U0_ifmap_vec_ce0),
    .i_we0(tdf10_readInputs69_U0_ifmap_vec_we0),
    .i_address0(tdf10_readInputs69_U0_ifmap_vec_address0),
    .i_d0(tdf10_readInputs69_U0_ifmap_vec_d0),
    .i_q0(ifmap_vec_i_q0),
    .i_ce1(tdf10_readInputs69_U0_ifmap_vec_ce1),
    .i_we1(tdf10_readInputs69_U0_ifmap_vec_we1),
    .i_address1(tdf10_readInputs69_U0_ifmap_vec_address1),
    .i_d1(tdf10_readInputs69_U0_ifmap_vec_d1),
    .t_ce(1'b1),
    .t_read(tdf10_dot_product_U0_ap_ready),
    .t_empty_n(ifmap_vec_t_empty_n),
    .t_ce0(tdf10_dot_product_U0_ifmap_vec_ce0),
    .t_we0(1'b0),
    .t_address0(tdf10_dot_product_U0_ifmap_vec_address0),
    .t_d0(16'd0),
    .t_q0(ifmap_vec_t_q0),
    .t_ce1(1'b0),
    .t_we1(1'b0),
    .t_address1(10'd0),
    .t_d1(16'd0)
);

td_fused_top_dataflow_in_loop_TOP_LOOP38364_ifmap_vec #(
    .DataWidth( 16 ),
    .AddressRange( 576 ),
    .AddressWidth( 10 ))
weight_vecs_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf10_readFilters68_U0_ap_done),
    .i_full_n(weight_vecs_0_i_full_n),
    .i_ce0(tdf10_readFilters68_U0_weight_vecs_0_ce0),
    .i_we0(tdf10_readFilters68_U0_weight_vecs_0_we0),
    .i_address0(tdf10_readFilters68_U0_weight_vecs_0_address0),
    .i_d0(tdf10_readFilters68_U0_weight_vecs_0_d0),
    .i_q0(weight_vecs_0_i_q0),
    .i_ce1(tdf10_readFilters68_U0_weight_vecs_0_ce1),
    .i_we1(tdf10_readFilters68_U0_weight_vecs_0_we1),
    .i_address1(tdf10_readFilters68_U0_weight_vecs_0_address1),
    .i_d1(tdf10_readFilters68_U0_weight_vecs_0_d1),
    .t_ce(1'b1),
    .t_read(tdf10_dot_product_U0_ap_ready),
    .t_empty_n(weight_vecs_0_t_empty_n),
    .t_ce0(tdf10_dot_product_U0_weight_vecs_0_ce0),
    .t_we0(1'b0),
    .t_address0(tdf10_dot_product_U0_weight_vecs_0_address0),
    .t_d0(16'd0),
    .t_q0(weight_vecs_0_t_q0),
    .t_ce1(1'b0),
    .t_we1(1'b0),
    .t_address1(10'd0),
    .t_d1(16'd0)
);

td_fused_top_dataflow_in_loop_TOP_LOOP38364_products_0 #(
    .DataWidth( 16 ),
    .AddressRange( 576 ),
    .AddressWidth( 10 ))
products_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf10_dot_product_U0_ap_done),
    .i_full_n(products_0_i_full_n),
    .i_ce0(tdf10_dot_product_U0_products_0_ce0),
    .i_we0(tdf10_dot_product_U0_products_0_we0),
    .i_address0(tdf10_dot_product_U0_products_0_address0),
    .i_d0(tdf10_dot_product_U0_products_0_d0),
    .i_q0(products_0_i_q0),
    .i_ce1(1'b0),
    .i_address1(10'd0),
    .i_q1(products_0_i_q1),
    .t_ce(1'b1),
    .t_read(tdf10_accum_1_U0_ap_ready),
    .t_empty_n(products_0_t_empty_n),
    .t_ce0(tdf10_accum_1_U0_accum_in_0_ce0),
    .t_we0(1'b0),
    .t_address0(tdf10_accum_1_U0_accum_in_0_address0),
    .t_d0(16'd0),
    .t_q0(products_0_t_q0),
    .t_ce1(tdf10_accum_1_U0_accum_in_0_ce1),
    .t_address1(tdf10_accum_1_U0_accum_in_0_address1),
    .t_q1(products_0_t_q1)
);

td_fused_top_dataflow_in_loop_TOP_LOOP38364_accum1_out_0 #(
    .DataWidth( 16 ),
    .AddressRange( 8 ),
    .AddressWidth( 3 ))
accum1_out_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf10_accum_1_U0_ap_done),
    .i_full_n(accum1_out_0_i_full_n),
    .i_ce0(tdf10_accum_1_U0_accum_out_ce0),
    .i_we0(tdf10_accum_1_U0_accum_out_we0),
    .i_address0(tdf10_accum_1_U0_accum_out_address0),
    .i_d0(tdf10_accum_1_U0_accum_out_d0),
    .i_q0(accum1_out_0_i_q0),
    .i_ce1(tdf10_accum_1_U0_accum_out_ce1),
    .i_we1(tdf10_accum_1_U0_accum_out_we1),
    .i_address1(tdf10_accum_1_U0_accum_out_address1),
    .i_d1(tdf10_accum_1_U0_accum_out_d1),
    .t_ce(1'b1),
    .t_read(tdf10_accum_2_U0_ap_ready),
    .t_empty_n(accum1_out_0_t_empty_n),
    .t_ce0(tdf10_accum_2_U0_accum_in_ce0),
    .t_we0(1'b0),
    .t_address0(tdf10_accum_2_U0_accum_in_address0),
    .t_d0(16'd0),
    .t_q0(accum1_out_0_t_q0),
    .t_ce1(1'b0),
    .t_we1(1'b0),
    .t_address1(3'd0),
    .t_d1(16'd0)
);

td_fused_top_dataflow_in_loop_TOP_LOOP38364_l2_products #(
    .DataWidth( 16 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
l2_products_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf10_l2_multiply66_U0_ap_done),
    .i_full_n(l2_products_i_full_n),
    .i_ce0(tdf10_l2_multiply66_U0_l2_products_ce0),
    .i_we0(tdf10_l2_multiply66_U0_l2_products_we0),
    .i_address0(tdf10_l2_multiply66_U0_l2_products_address0),
    .i_d0(tdf10_l2_multiply66_U0_l2_products_d0),
    .i_q0(l2_products_i_q0),
    .t_ce(1'b1),
    .t_read(tdf10_l2_writeOutputs_165_U0_ap_ready),
    .t_empty_n(l2_products_t_empty_n),
    .t_ce0(tdf10_l2_writeOutputs_165_U0_l2_partial_sums_ce0),
    .t_we0(1'b0),
    .t_address0(tdf10_l2_writeOutputs_165_U0_l2_partial_sums_address0),
    .t_d0(16'd0),
    .t_q0(l2_products_t_q0)
);

td_fused_top_tdf10_get_next_ijk tdf10_get_next_ijk_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf10_get_next_ijk_U0_ap_start),
    .start_full_n(start_for_tdf10_readFilters68_U0_full_n),
    .ap_done(tdf10_get_next_ijk_U0_ap_done),
    .ap_continue(tdf10_get_next_ijk_U0_ap_continue),
    .ap_idle(tdf10_get_next_ijk_U0_ap_idle),
    .ap_ready(tdf10_get_next_ijk_U0_ap_ready),
    .start_out(tdf10_get_next_ijk_U0_start_out),
    .start_write(tdf10_get_next_ijk_U0_start_write),
    .indices_0_din(tdf10_get_next_ijk_U0_indices_0_din),
    .indices_0_full_n(indices_01_c_full_n),
    .indices_0_write(tdf10_get_next_ijk_U0_indices_0_write),
    .indices_1_din(tdf10_get_next_ijk_U0_indices_1_din),
    .indices_1_full_n(indices_12_c_full_n),
    .indices_1_write(tdf10_get_next_ijk_U0_indices_1_write),
    .indices_2_out_din(tdf10_get_next_ijk_U0_indices_2_out_din),
    .indices_2_out_full_n(indices_23_c_full_n),
    .indices_2_out_write(tdf10_get_next_ijk_U0_indices_2_out_write),
    .indices_2_out1_din(tdf10_get_next_ijk_U0_indices_2_out1_din),
    .indices_2_out1_full_n(indices_23_c1_full_n),
    .indices_2_out1_write(tdf10_get_next_ijk_U0_indices_2_out1_write),
    .write_r_din(tdf10_get_next_ijk_U0_write_r_din),
    .write_r_full_n(write4_c_full_n),
    .write_r_write(tdf10_get_next_ijk_U0_write_r_write)
);

td_fused_top_tdf10_readInputs69 tdf10_readInputs69_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf10_readInputs69_U0_ap_start),
    .ap_done(tdf10_readInputs69_U0_ap_done),
    .ap_continue(tdf10_readInputs69_U0_ap_continue),
    .ap_idle(tdf10_readInputs69_U0_ap_idle),
    .ap_ready(tdf10_readInputs69_U0_ap_ready),
    .in_data_address0(tdf10_readInputs69_U0_in_data_address0),
    .in_data_ce0(tdf10_readInputs69_U0_in_data_ce0),
    .in_data_q0(in_data_q0),
    .indices_01_dout(indices_01_c_dout),
    .indices_01_empty_n(indices_01_c_empty_n),
    .indices_01_read(tdf10_readInputs69_U0_indices_01_read),
    .indices_12_dout(indices_12_c_dout),
    .indices_12_empty_n(indices_12_c_empty_n),
    .indices_12_read(tdf10_readInputs69_U0_indices_12_read),
    .ifmap_vec_address0(tdf10_readInputs69_U0_ifmap_vec_address0),
    .ifmap_vec_ce0(tdf10_readInputs69_U0_ifmap_vec_ce0),
    .ifmap_vec_we0(tdf10_readInputs69_U0_ifmap_vec_we0),
    .ifmap_vec_d0(tdf10_readInputs69_U0_ifmap_vec_d0),
    .ifmap_vec_address1(tdf10_readInputs69_U0_ifmap_vec_address1),
    .ifmap_vec_ce1(tdf10_readInputs69_U0_ifmap_vec_ce1),
    .ifmap_vec_we1(tdf10_readInputs69_U0_ifmap_vec_we1),
    .ifmap_vec_d1(tdf10_readInputs69_U0_ifmap_vec_d1),
    .indices_01_out_din(tdf10_readInputs69_U0_indices_01_out_din),
    .indices_01_out_full_n(indices_01_c2_full_n),
    .indices_01_out_write(tdf10_readInputs69_U0_indices_01_out_write),
    .indices_12_out_din(tdf10_readInputs69_U0_indices_12_out_din),
    .indices_12_out_full_n(indices_12_c3_full_n),
    .indices_12_out_write(tdf10_readInputs69_U0_indices_12_out_write)
);

td_fused_top_tdf10_readFilters68 tdf10_readFilters68_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf10_readFilters68_U0_ap_start),
    .ap_done(tdf10_readFilters68_U0_ap_done),
    .ap_continue(tdf10_readFilters68_U0_ap_continue),
    .ap_idle(tdf10_readFilters68_U0_ap_idle),
    .ap_ready(tdf10_readFilters68_U0_ap_ready),
    .filter_data_address0(tdf10_readFilters68_U0_filter_data_address0),
    .filter_data_ce0(tdf10_readFilters68_U0_filter_data_ce0),
    .filter_data_q0(l1_filter_data_q0),
    .indices_23_dout(indices_23_c_dout),
    .indices_23_empty_n(indices_23_c_empty_n),
    .indices_23_read(tdf10_readFilters68_U0_indices_23_read),
    .weight_vecs_0_address0(tdf10_readFilters68_U0_weight_vecs_0_address0),
    .weight_vecs_0_ce0(tdf10_readFilters68_U0_weight_vecs_0_ce0),
    .weight_vecs_0_we0(tdf10_readFilters68_U0_weight_vecs_0_we0),
    .weight_vecs_0_d0(tdf10_readFilters68_U0_weight_vecs_0_d0),
    .weight_vecs_0_address1(tdf10_readFilters68_U0_weight_vecs_0_address1),
    .weight_vecs_0_ce1(tdf10_readFilters68_U0_weight_vecs_0_ce1),
    .weight_vecs_0_we1(tdf10_readFilters68_U0_weight_vecs_0_we1),
    .weight_vecs_0_d1(tdf10_readFilters68_U0_weight_vecs_0_d1)
);

td_fused_top_tdf10_dot_product tdf10_dot_product_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf10_dot_product_U0_ap_start),
    .ap_done(tdf10_dot_product_U0_ap_done),
    .ap_continue(tdf10_dot_product_U0_ap_continue),
    .ap_idle(tdf10_dot_product_U0_ap_idle),
    .ap_ready(tdf10_dot_product_U0_ap_ready),
    .ifmap_vec_address0(tdf10_dot_product_U0_ifmap_vec_address0),
    .ifmap_vec_ce0(tdf10_dot_product_U0_ifmap_vec_ce0),
    .ifmap_vec_q0(ifmap_vec_t_q0),
    .weight_vecs_0_address0(tdf10_dot_product_U0_weight_vecs_0_address0),
    .weight_vecs_0_ce0(tdf10_dot_product_U0_weight_vecs_0_ce0),
    .weight_vecs_0_q0(weight_vecs_0_t_q0),
    .products_0_address0(tdf10_dot_product_U0_products_0_address0),
    .products_0_ce0(tdf10_dot_product_U0_products_0_ce0),
    .products_0_we0(tdf10_dot_product_U0_products_0_we0),
    .products_0_d0(tdf10_dot_product_U0_products_0_d0)
);

td_fused_top_tdf10_accum_1 tdf10_accum_1_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf10_accum_1_U0_ap_start),
    .ap_done(tdf10_accum_1_U0_ap_done),
    .ap_continue(tdf10_accum_1_U0_ap_continue),
    .ap_idle(tdf10_accum_1_U0_ap_idle),
    .ap_ready(tdf10_accum_1_U0_ap_ready),
    .accum_in_0_address0(tdf10_accum_1_U0_accum_in_0_address0),
    .accum_in_0_ce0(tdf10_accum_1_U0_accum_in_0_ce0),
    .accum_in_0_q0(products_0_t_q0),
    .accum_in_0_address1(tdf10_accum_1_U0_accum_in_0_address1),
    .accum_in_0_ce1(tdf10_accum_1_U0_accum_in_0_ce1),
    .accum_in_0_q1(products_0_t_q1),
    .accum_out_address0(tdf10_accum_1_U0_accum_out_address0),
    .accum_out_ce0(tdf10_accum_1_U0_accum_out_ce0),
    .accum_out_we0(tdf10_accum_1_U0_accum_out_we0),
    .accum_out_d0(tdf10_accum_1_U0_accum_out_d0),
    .accum_out_address1(tdf10_accum_1_U0_accum_out_address1),
    .accum_out_ce1(tdf10_accum_1_U0_accum_out_ce1),
    .accum_out_we1(tdf10_accum_1_U0_accum_out_we1),
    .accum_out_d1(tdf10_accum_1_U0_accum_out_d1)
);

td_fused_top_tdf10_accum_2 tdf10_accum_2_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf10_accum_2_U0_ap_start),
    .ap_done(tdf10_accum_2_U0_ap_done),
    .ap_continue(tdf10_accum_2_U0_ap_continue),
    .ap_idle(tdf10_accum_2_U0_ap_idle),
    .ap_ready(tdf10_accum_2_U0_ap_ready),
    .accum_in_24(tdf10_accum_2_U0_accum_in_24),
    .accum_in_24_ap_vld(tdf10_accum_2_U0_accum_in_24_ap_vld),
    .accum_in_address0(tdf10_accum_2_U0_accum_in_address0),
    .accum_in_ce0(tdf10_accum_2_U0_accum_in_ce0),
    .accum_in_q0(accum1_out_0_t_q0)
);

td_fused_top_Block_entry_proc_proc435 Block_entry_proc_proc435_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(Block_entry_proc_proc435_U0_ap_start),
    .ap_done(Block_entry_proc_proc435_U0_ap_done),
    .ap_continue(Block_entry_proc_proc435_U0_ap_continue),
    .ap_idle(Block_entry_proc_proc435_U0_ap_idle),
    .ap_ready(Block_entry_proc_proc435_U0_ap_ready),
    .tmp(tmp_channel_dout),
    .ap_return(Block_entry_proc_proc435_U0_ap_return)
);

td_fused_top_tdf10_adjust tdf10_adjust_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf10_adjust_U0_ap_start),
    .ap_done(tdf10_adjust_U0_ap_done),
    .ap_continue(tdf10_adjust_U0_ap_continue),
    .ap_idle(tdf10_adjust_U0_ap_idle),
    .ap_ready(tdf10_adjust_U0_ap_ready),
    .sums_read(sums_0_dout),
    .adjustments_address0(tdf10_adjust_U0_adjustments_address0),
    .adjustments_ce0(tdf10_adjust_U0_adjustments_ce0),
    .adjustments_q0(l1_adjustments_q0),
    .indices_23_dout(indices_23_c1_dout),
    .indices_23_empty_n(indices_23_c1_empty_n),
    .indices_23_read(tdf10_adjust_U0_indices_23_read),
    .indices_23_out_din(tdf10_adjust_U0_indices_23_out_din),
    .indices_23_out_full_n(indices_23_c4_full_n),
    .indices_23_out_write(tdf10_adjust_U0_indices_23_out_write),
    .ap_return(tdf10_adjust_U0_ap_return)
);

td_fused_top_tdf10_l2_multiply66 tdf10_l2_multiply66_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf10_l2_multiply66_U0_ap_start),
    .ap_done(tdf10_l2_multiply66_U0_ap_done),
    .ap_continue(tdf10_l2_multiply66_U0_ap_continue),
    .ap_idle(tdf10_l2_multiply66_U0_ap_idle),
    .ap_ready(tdf10_l2_multiply66_U0_ap_ready),
    .intermediate_fmaps_read(intermediate_fmaps_0_dout),
    .l2_filter_data_address0(tdf10_l2_multiply66_U0_l2_filter_data_address0),
    .l2_filter_data_ce0(tdf10_l2_multiply66_U0_l2_filter_data_ce0),
    .l2_filter_data_q0(l2_filter_data_q0),
    .l2_products_address0(tdf10_l2_multiply66_U0_l2_products_address0),
    .l2_products_ce0(tdf10_l2_multiply66_U0_l2_products_ce0),
    .l2_products_we0(tdf10_l2_multiply66_U0_l2_products_we0),
    .l2_products_d0(tdf10_l2_multiply66_U0_l2_products_d0),
    .indices_23_dout(indices_23_c4_dout),
    .indices_23_empty_n(indices_23_c4_empty_n),
    .indices_23_read(tdf10_l2_multiply66_U0_indices_23_read)
);

td_fused_top_tdf10_l2_writeOutputs_165 tdf10_l2_writeOutputs_165_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf10_l2_writeOutputs_165_U0_ap_start),
    .ap_done(tdf10_l2_writeOutputs_165_U0_ap_done),
    .ap_continue(tdf10_l2_writeOutputs_165_U0_ap_continue),
    .ap_idle(tdf10_l2_writeOutputs_165_U0_ap_idle),
    .ap_ready(tdf10_l2_writeOutputs_165_U0_ap_ready),
    .indices_01_dout(indices_01_c2_dout),
    .indices_01_empty_n(indices_01_c2_empty_n),
    .indices_01_read(tdf10_l2_writeOutputs_165_U0_indices_01_read),
    .indices_12_dout(indices_12_c3_dout),
    .indices_12_empty_n(indices_12_c3_empty_n),
    .indices_12_read(tdf10_l2_writeOutputs_165_U0_indices_12_read),
    .write4_dout(write4_c_dout),
    .write4_empty_n(write4_c_empty_n),
    .write4_read(tdf10_l2_writeOutputs_165_U0_write4_read),
    .l2_partial_sums_address0(tdf10_l2_writeOutputs_165_U0_l2_partial_sums_address0),
    .l2_partial_sums_ce0(tdf10_l2_writeOutputs_165_U0_l2_partial_sums_ce0),
    .l2_partial_sums_q0(l2_products_t_q0),
    .out_data_address1(tdf10_l2_writeOutputs_165_U0_out_data_address1),
    .out_data_ce1(tdf10_l2_writeOutputs_165_U0_out_data_ce1),
    .out_data_we1(tdf10_l2_writeOutputs_165_U0_out_data_we1),
    .out_data_d1(tdf10_l2_writeOutputs_165_U0_out_data_d1),
    .l2_adjustments_address0(tdf10_l2_writeOutputs_165_U0_l2_adjustments_address0),
    .l2_adjustments_ce0(tdf10_l2_writeOutputs_165_U0_l2_adjustments_ce0),
    .l2_adjustments_q0(l2_adjustments_q0)
);

td_fused_top_fifo_w16_d2_S_x7 indices_01_c_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(indices_01_c_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf10_readInputs69_U0_indices_01_read),
    .if_dout(indices_01_c_dout),
    .if_full_n(indices_01_c_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf10_get_next_ijk_U0_indices_0_write),
    .if_din(tdf10_get_next_ijk_U0_indices_0_din)
);

td_fused_top_fifo_w16_d2_S_x7 indices_12_c_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(indices_12_c_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf10_readInputs69_U0_indices_12_read),
    .if_dout(indices_12_c_dout),
    .if_full_n(indices_12_c_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf10_get_next_ijk_U0_indices_1_write),
    .if_din(tdf10_get_next_ijk_U0_indices_1_din)
);

td_fused_top_fifo_w9_d2_S indices_23_c_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(indices_23_c_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf10_readFilters68_U0_indices_23_read),
    .if_dout(indices_23_c_dout),
    .if_full_n(indices_23_c_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf10_get_next_ijk_U0_indices_2_out_write),
    .if_din(tdf10_get_next_ijk_U0_indices_2_out_din)
);

td_fused_top_fifo_w15_d7_S indices_23_c1_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(indices_23_c1_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf10_adjust_U0_indices_23_read),
    .if_dout(indices_23_c1_dout),
    .if_full_n(indices_23_c1_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf10_get_next_ijk_U0_indices_2_out1_write),
    .if_din(tdf10_get_next_ijk_U0_indices_2_out1_din)
);

td_fused_top_fifo_w1_d9_S_x1 write4_c_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(write4_c_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf10_l2_writeOutputs_165_U0_write4_read),
    .if_dout(write4_c_dout),
    .if_full_n(write4_c_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf10_get_next_ijk_U0_write_r_write),
    .if_din(write4_c_din)
);

td_fused_top_fifo_w4_d8_S_x0 indices_01_c2_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(indices_01_c2_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf10_l2_writeOutputs_165_U0_indices_01_read),
    .if_dout(indices_01_c2_dout),
    .if_full_n(indices_01_c2_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf10_readInputs69_U0_indices_01_out_write),
    .if_din(tdf10_readInputs69_U0_indices_01_out_din)
);

td_fused_top_fifo_w8_d8_S_x indices_12_c3_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(indices_12_c3_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf10_l2_writeOutputs_165_U0_indices_12_read),
    .if_dout(indices_12_c3_dout),
    .if_full_n(indices_12_c3_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf10_readInputs69_U0_indices_12_out_write),
    .if_din(tdf10_readInputs69_U0_indices_12_out_din)
);

td_fused_top_fifo_w16_d2_S_x7 tmp_channel_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(tmp_channel_empty_n),
    .if_read_ce(1'b1),
    .if_read(Block_entry_proc_proc435_U0_ap_ready),
    .if_dout(tmp_channel_dout),
    .if_full_n(tmp_channel_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf10_accum_2_U0_ap_done),
    .if_din(tdf10_accum_2_U0_accum_in_24)
);

td_fused_top_fifo_w16_d2_S_x7 sums_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(sums_0_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf10_adjust_U0_ap_ready),
    .if_dout(sums_0_dout),
    .if_full_n(sums_0_full_n),
    .if_write_ce(1'b1),
    .if_write(Block_entry_proc_proc435_U0_ap_done),
    .if_din(Block_entry_proc_proc435_U0_ap_return)
);

td_fused_top_fifo_w15_d2_S indices_23_c4_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(indices_23_c4_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf10_l2_multiply66_U0_indices_23_read),
    .if_dout(indices_23_c4_dout),
    .if_full_n(indices_23_c4_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf10_adjust_U0_indices_23_out_write),
    .if_din(tdf10_adjust_U0_indices_23_out_din)
);

td_fused_top_fifo_w16_d2_S_x7 intermediate_fmaps_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(intermediate_fmaps_0_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf10_l2_multiply66_U0_ap_ready),
    .if_dout(intermediate_fmaps_0_dout),
    .if_full_n(intermediate_fmaps_0_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf10_adjust_U0_ap_done),
    .if_din(tdf10_adjust_U0_ap_return)
);

td_fused_top_start_for_tdf10_readFilters68_U0 start_for_tdf10_readFilters68_U0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(start_for_tdf10_readFilters68_U0_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf10_readFilters68_U0_ap_ready),
    .if_dout(start_for_tdf10_readFilters68_U0_dout),
    .if_full_n(start_for_tdf10_readFilters68_U0_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf10_get_next_ijk_U0_start_write),
    .if_din(start_for_tdf10_readFilters68_U0_din)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_sync_reg_tdf10_get_next_ijk_U0_ap_ready <= 1'b0;
    end else begin
        if (((ap_sync_ready & ap_start) == 1'b1)) begin
            ap_sync_reg_tdf10_get_next_ijk_U0_ap_ready <= 1'b0;
        end else begin
            ap_sync_reg_tdf10_get_next_ijk_U0_ap_ready <= ap_sync_tdf10_get_next_ijk_U0_ap_ready;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_sync_reg_tdf10_readInputs69_U0_ap_ready <= 1'b0;
    end else begin
        if (((ap_sync_ready & ap_start) == 1'b1)) begin
            ap_sync_reg_tdf10_readInputs69_U0_ap_ready <= 1'b0;
        end else begin
            ap_sync_reg_tdf10_readInputs69_U0_ap_ready <= ap_sync_tdf10_readInputs69_U0_ap_ready;
        end
    end
end

assign Block_entry_proc_proc435_U0_ap_continue = sums_0_full_n;

assign Block_entry_proc_proc435_U0_ap_start = tmp_channel_empty_n;

assign Block_entry_proc_proc435_U0_start_full_n = 1'b1;

assign Block_entry_proc_proc435_U0_start_write = 1'b0;

assign ap_channel_done_accum1_out_0 = tdf10_accum_1_U0_ap_done;

assign ap_channel_done_ifmap_vec = tdf10_readInputs69_U0_ap_done;

assign ap_channel_done_intermediate_fmaps_0 = tdf10_adjust_U0_ap_done;

assign ap_channel_done_l2_products = tdf10_l2_multiply66_U0_ap_done;

assign ap_channel_done_products_0 = tdf10_dot_product_U0_ap_done;

assign ap_channel_done_sums_0 = Block_entry_proc_proc435_U0_ap_done;

assign ap_channel_done_tmp_channel = tdf10_accum_2_U0_ap_done;

assign ap_channel_done_weight_vecs_0 = tdf10_readFilters68_U0_ap_done;

assign ap_done = tdf10_l2_writeOutputs_165_U0_ap_done;

assign ap_idle = (tdf10_readInputs69_U0_ap_idle & tdf10_readFilters68_U0_ap_idle & tdf10_l2_writeOutputs_165_U0_ap_idle & tdf10_l2_multiply66_U0_ap_idle & tdf10_get_next_ijk_U0_ap_idle & tdf10_dot_product_U0_ap_idle & tdf10_adjust_U0_ap_idle & tdf10_accum_2_U0_ap_idle & tdf10_accum_1_U0_ap_idle & (intermediate_fmaps_0_empty_n ^ 1'b1) & (sums_0_empty_n ^ 1'b1) & (tmp_channel_empty_n ^ 1'b1) & (l2_products_t_empty_n ^ 1'b1) & (products_0_t_empty_n ^ 1'b1) & (weight_vecs_0_t_empty_n ^ 1'b1) & (ifmap_vec_t_empty_n ^ 1'b1) & (1'b1 ^ accum1_out_0_t_empty_n) & Block_entry_proc_proc435_U0_ap_idle);

assign ap_ready = ap_sync_ready;

assign ap_sync_continue = ap_continue;

assign ap_sync_done = tdf10_l2_writeOutputs_165_U0_ap_done;

assign ap_sync_ready = (ap_sync_tdf10_readInputs69_U0_ap_ready & ap_sync_tdf10_get_next_ijk_U0_ap_ready);

assign ap_sync_tdf10_get_next_ijk_U0_ap_ready = (tdf10_get_next_ijk_U0_ap_ready | ap_sync_reg_tdf10_get_next_ijk_U0_ap_ready);

assign ap_sync_tdf10_readInputs69_U0_ap_ready = (tdf10_readInputs69_U0_ap_ready | ap_sync_reg_tdf10_readInputs69_U0_ap_ready);

assign in_data_address0 = tdf10_readInputs69_U0_in_data_address0;

assign in_data_address1 = 12'd0;

assign in_data_ce0 = tdf10_readInputs69_U0_in_data_ce0;

assign in_data_ce1 = 1'b0;

assign in_data_d0 = 64'd0;

assign in_data_d1 = 64'd0;

assign in_data_read = tdf10_readInputs69_U0_in_data_write;

assign in_data_we0 = 1'b0;

assign in_data_we1 = 1'b0;

assign l1_adjustments_address0 = tdf10_adjust_U0_adjustments_address0;

assign l1_adjustments_address1 = 9'd0;

assign l1_adjustments_ce0 = tdf10_adjust_U0_adjustments_ce0;

assign l1_adjustments_ce1 = 1'b0;

assign l1_adjustments_d0 = 48'd0;

assign l1_adjustments_d1 = 48'd0;

assign l1_adjustments_we0 = 1'b0;

assign l1_adjustments_we1 = 1'b0;

assign l1_filter_data_address0 = tdf10_readFilters68_U0_filter_data_address0;

assign l1_filter_data_address1 = 17'd0;

assign l1_filter_data_ce0 = tdf10_readFilters68_U0_filter_data_ce0;

assign l1_filter_data_ce1 = 1'b0;

assign l1_filter_data_d0 = 64'd0;

assign l1_filter_data_d1 = 64'd0;

assign l1_filter_data_we0 = 1'b0;

assign l1_filter_data_we1 = 1'b0;

assign l2_adjustments_address0 = tdf10_l2_writeOutputs_165_U0_l2_adjustments_address0;

assign l2_adjustments_address1 = 6'd0;

assign l2_adjustments_ce0 = tdf10_l2_writeOutputs_165_U0_l2_adjustments_ce0;

assign l2_adjustments_ce1 = 1'b0;

assign l2_adjustments_d0 = 48'd0;

assign l2_adjustments_d1 = 48'd0;

assign l2_adjustments_we0 = 1'b0;

assign l2_adjustments_we1 = 1'b0;

assign l2_filter_data_address0 = tdf10_l2_multiply66_U0_l2_filter_data_address0;

assign l2_filter_data_address1 = 15'd0;

assign l2_filter_data_ce0 = tdf10_l2_multiply66_U0_l2_filter_data_ce0;

assign l2_filter_data_ce1 = 1'b0;

assign l2_filter_data_d0 = 16'd0;

assign l2_filter_data_d1 = 16'd0;

assign l2_filter_data_we0 = 1'b0;

assign l2_filter_data_we1 = 1'b0;

assign out_data_address0 = 12'd0;

assign out_data_address1 = tdf10_l2_writeOutputs_165_U0_out_data_address1;

assign out_data_ce0 = 1'b0;

assign out_data_ce1 = tdf10_l2_writeOutputs_165_U0_out_data_ce1;

assign out_data_d0 = 64'd0;

assign out_data_d1 = tdf10_l2_writeOutputs_165_U0_out_data_d1;

assign out_data_we0 = 1'b0;

assign out_data_we1 = tdf10_l2_writeOutputs_165_U0_out_data_we1;

assign out_data_write = tdf10_l2_writeOutputs_165_U0_out_data_write;

assign products_0_t_d1 = 16'd0;

assign products_0_t_we1 = 1'b0;

assign start_for_tdf10_readFilters68_U0_din = 1'b1;

assign tdf10_accum_1_U0_accum_out_full_n = accum1_out_0_i_full_n;

assign tdf10_accum_1_U0_ap_continue = accum1_out_0_i_full_n;

assign tdf10_accum_1_U0_ap_start = products_0_t_empty_n;

assign tdf10_accum_1_U0_start_full_n = 1'b1;

assign tdf10_accum_1_U0_start_write = 1'b0;

assign tdf10_accum_2_U0_ap_continue = tmp_channel_full_n;

assign tdf10_accum_2_U0_ap_start = accum1_out_0_t_empty_n;

assign tdf10_accum_2_U0_start_full_n = 1'b1;

assign tdf10_accum_2_U0_start_write = 1'b0;

assign tdf10_adjust_U0_ap_continue = intermediate_fmaps_0_full_n;

assign tdf10_adjust_U0_ap_start = sums_0_empty_n;

assign tdf10_adjust_U0_start_full_n = 1'b1;

assign tdf10_adjust_U0_start_write = 1'b0;

assign tdf10_dot_product_U0_ap_continue = products_0_i_full_n;

assign tdf10_dot_product_U0_ap_start = (weight_vecs_0_t_empty_n & ifmap_vec_t_empty_n);

assign tdf10_dot_product_U0_products_0_full_n = products_0_i_full_n;

assign tdf10_dot_product_U0_start_full_n = 1'b1;

assign tdf10_dot_product_U0_start_write = 1'b0;

assign tdf10_get_next_ijk_U0_ap_continue = 1'b1;

assign tdf10_get_next_ijk_U0_ap_start = ((ap_sync_reg_tdf10_get_next_ijk_U0_ap_ready ^ 1'b1) & ap_start);

assign tdf10_l2_multiply66_U0_ap_continue = l2_products_i_full_n;

assign tdf10_l2_multiply66_U0_ap_start = intermediate_fmaps_0_empty_n;

assign tdf10_l2_multiply66_U0_l2_products_full_n = l2_products_i_full_n;

assign tdf10_l2_multiply66_U0_start_full_n = 1'b1;

assign tdf10_l2_multiply66_U0_start_write = 1'b0;

assign tdf10_l2_writeOutputs_165_U0_ap_continue = ap_continue;

assign tdf10_l2_writeOutputs_165_U0_ap_start = l2_products_t_empty_n;

assign tdf10_l2_writeOutputs_165_U0_out_data_full_n = out_data_full_n;

assign tdf10_l2_writeOutputs_165_U0_out_data_write = 1'b0;

assign tdf10_l2_writeOutputs_165_U0_start_full_n = 1'b1;

assign tdf10_l2_writeOutputs_165_U0_start_write = 1'b0;

assign tdf10_readFilters68_U0_ap_continue = weight_vecs_0_i_full_n;

assign tdf10_readFilters68_U0_ap_start = start_for_tdf10_readFilters68_U0_empty_n;

assign tdf10_readFilters68_U0_start_full_n = 1'b1;

assign tdf10_readFilters68_U0_start_write = 1'b0;

assign tdf10_readFilters68_U0_weight_vecs_0_full_n = weight_vecs_0_i_full_n;

assign tdf10_readInputs69_U0_ap_continue = ifmap_vec_i_full_n;

assign tdf10_readInputs69_U0_ap_start = ((ap_sync_reg_tdf10_readInputs69_U0_ap_ready ^ 1'b1) & ap_start);

assign tdf10_readInputs69_U0_ifmap_vec_full_n = ifmap_vec_i_full_n;

assign tdf10_readInputs69_U0_in_data_full_n = in_data_empty_n;

assign tdf10_readInputs69_U0_in_data_write = 1'b0;

assign tdf10_readInputs69_U0_start_full_n = 1'b1;

assign tdf10_readInputs69_U0_start_write = 1'b0;

assign write4_c_din = tdf10_get_next_ijk_U0_write_r_din;

endmodule //td_fused_top_dataflow_in_loop_TOP_LOOP38364
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP76_accum1_out_0_memcore_ram (addr0, ce0, d0, we0, q0, addr1, ce1, d1, we1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 3;
parameter MEM_SIZE = 8;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
input clk;

reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];




always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1) 
            ram[addr1] <= d1; 
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP76_accum1_out_0_memcore(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    q0,
    address1,
    ce1,
    we1,
    d1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd8;
parameter AddressWidth = 32'd3;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;



td_fused_top_dataflow_in_loop_TOP_LOOP76_accum1_out_0_memcore_ram td_fused_top_dataflow_in_loop_TOP_LOOP76_accum1_out_0_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_dataflow_in_loop_TOP_LOOP76_accum1_out_0
#(parameter
    DataWidth    = 16,
    AddressRange = 32,
    AddressWidth = 3,
    BufferCount  = 2,
    MemLatency   = 1,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire                    i_we0,
    input  wire [AddressWidth-1:0] i_address0,
    input  wire [DataWidth-1:0]    i_d0,
    output wire [DataWidth-1:0]    i_q0,
    input  wire                    i_ce1,
    input  wire                    i_we1,
    input  wire [AddressWidth-1:0] i_address1,
    input  wire [DataWidth-1:0]    i_d1,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire                    t_we0,
    input  wire [AddressWidth-1:0] t_address0,
    input  wire [DataWidth-1:0]    t_d0,
    output wire [DataWidth-1:0]    t_q0,
    input  wire                    t_ce1,
    input  wire                    t_we1,
    input  wire [AddressWidth-1:0] t_address1,
    input  wire [DataWidth-1:0]    t_d1
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth-1:0]   prev_iptr    = 1'b0; // previous initiator index
reg  [IndexWidth-1:0]   prev_tptr    = 1'b0; // previous target index
reg  [DataWidth-1:0]    reg_q0      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid0    = 1'b0; // buffer has valid data
reg  [DataWidth-1:0]    reg_q1      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid1    = 1'b0; // buffer has valid data
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
// buffer signals
wire [BufferCount-1:0] buf_ce0;
wire [BufferCount-1:0] buf_we0;
wire [AddressWidth-1:0] buf_a0_0, buf_a0_1;
wire [DataWidth-1:0] buf_d0_0, buf_d0_1;
wire [DataWidth-1:0] buf_q0_0, buf_q0_1;
wire [BufferCount-1:0] buf_ce1;
wire [BufferCount-1:0] buf_we1;
wire [AddressWidth-1:0] buf_a1_0, buf_a1_1;
wire [DataWidth-1:0] buf_d1_0, buf_d1_1;
//------------------------Instantiation------------------
//genvar i;
        td_fused_top_dataflow_in_loop_TOP_LOOP76_accum1_out_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP76_accum1_out_0_memcore_U_0 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_0 ),
            .ce0      ( buf_ce0[ 0 ] ),
            .we0      ( buf_we0[ 0 ] ),
            .d0       ( buf_d0_0 ),
            .q0       ( buf_q0_0 ),
            .address1 ( buf_a1_0 ),
            .ce1      ( buf_ce1[ 0 ] ),
            .we1      ( buf_we1[ 0 ] ),
            .d1       ( buf_d1_0 )
        );
        td_fused_top_dataflow_in_loop_TOP_LOOP76_accum1_out_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP76_accum1_out_0_memcore_U_1 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_1 ),
            .ce0      ( buf_ce0[ 1 ] ),
            .we0      ( buf_we0[ 1 ] ),
            .d0       ( buf_d0_1 ),
            .q0       ( buf_q0_1 ),
            .address1 ( buf_a1_1 ),
            .ce1      ( buf_ce1[ 1 ] ),
            .we1      ( buf_we1[ 1 ] ),
            .d1       ( buf_d1_1 )
        );

//++++++++++++++++++++++++buffer signals+++++++++++++++++
        assign buf_ce0[ 0 ] = (tptr ==  0  && empty_n) ? t_ce0
                             : (iptr ==  0 ) ? i_ce0 : 1'b0;
        assign buf_a0_0  = (tptr ==  0  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 0 ] = (tptr ==  0  && empty_n)  ? t_we0
                             : (iptr ==  0 ) ? i_we0 : 1'b0;
        assign buf_d0_0  = (tptr ==  0  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 0 ] = (tptr ==  0  && empty_n) ? t_ce1
                             : (iptr ==  0 ) ? i_ce1 : 1'b0;
        assign buf_a1_0  = (tptr ==  0  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 0 ] = (tptr ==  0  && empty_n)  ? t_we1
                             : (iptr ==  0 ) ? i_we1 : 1'b0;
        assign buf_d1_0  = (tptr ==  0  && empty_n) ? t_d1       : i_d1;
        assign buf_ce0[ 1 ] = (tptr ==  1  && empty_n) ? t_ce0
                             : (iptr ==  1 ) ? i_ce0 : 1'b0;
        assign buf_a0_1  = (tptr ==  1  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 1 ] = (tptr ==  1  && empty_n)  ? t_we0
                             : (iptr ==  1 ) ? i_we0 : 1'b0;
        assign buf_d0_1  = (tptr ==  1  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 1 ] = (tptr ==  1  && empty_n) ? t_ce1
                             : (iptr ==  1 ) ? i_ce1 : 1'b0;
        assign buf_a1_1  = (tptr ==  1  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 1 ] = (tptr ==  1  && empty_n)  ? t_we1
                             : (iptr ==  1 ) ? i_we1 : 1'b0;
        assign buf_d1_1  = (tptr ==  1  && empty_n) ? t_d1       : i_d1;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//------------------------Body---------------------------
assign i_q0      = (prev_iptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign t_q0      = reg_valid0 ? reg_q0 : (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// prev_iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_iptr <= 1'b0;
    else begin
        prev_iptr <= iptr;
    end
end

// prev_tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_tptr <= 1'b0;
    else begin
        prev_tptr <= tptr;
    end
end

// reg_q0 and reg_valid0
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q0     <= 1'b0;
        reg_valid0 <= 1'b0;
    end else if (!t_ce0 && !reg_valid0) begin
        reg_q0     <= (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
        reg_valid0 <= 1'b1;
    end else if (t_ce0) begin
        reg_valid0 <= 1'b0;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP76_ifmap_vec_0_0_memcore_ram (addr0, ce0, d0, we0, q0, addr1, ce1, d1, we1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
input clk;

reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];




always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1) 
            ram[addr1] <= d1; 
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP76_ifmap_vec_0_0_memcore(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    q0,
    address1,
    ce1,
    we1,
    d1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;



td_fused_top_dataflow_in_loop_TOP_LOOP76_ifmap_vec_0_0_memcore_ram td_fused_top_dataflow_in_loop_TOP_LOOP76_ifmap_vec_0_0_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_dataflow_in_loop_TOP_LOOP76_ifmap_vec_0_0
#(parameter
    DataWidth    = 16,
    AddressRange = 32,
    AddressWidth = 7,
    BufferCount  = 2,
    MemLatency   = 1,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire                    i_we0,
    input  wire [AddressWidth-1:0] i_address0,
    input  wire [DataWidth-1:0]    i_d0,
    output wire [DataWidth-1:0]    i_q0,
    input  wire                    i_ce1,
    input  wire                    i_we1,
    input  wire [AddressWidth-1:0] i_address1,
    input  wire [DataWidth-1:0]    i_d1,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire                    t_we0,
    input  wire [AddressWidth-1:0] t_address0,
    input  wire [DataWidth-1:0]    t_d0,
    output wire [DataWidth-1:0]    t_q0,
    input  wire                    t_ce1,
    input  wire                    t_we1,
    input  wire [AddressWidth-1:0] t_address1,
    input  wire [DataWidth-1:0]    t_d1
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth-1:0]   prev_iptr    = 1'b0; // previous initiator index
reg  [IndexWidth-1:0]   prev_tptr    = 1'b0; // previous target index
reg  [DataWidth-1:0]    reg_q0      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid0    = 1'b0; // buffer has valid data
reg  [DataWidth-1:0]    reg_q1      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid1    = 1'b0; // buffer has valid data
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
// buffer signals
wire [BufferCount-1:0] buf_ce0;
wire [BufferCount-1:0] buf_we0;
wire [AddressWidth-1:0] buf_a0_0, buf_a0_1;
wire [DataWidth-1:0] buf_d0_0, buf_d0_1;
wire [DataWidth-1:0] buf_q0_0, buf_q0_1;
wire [BufferCount-1:0] buf_ce1;
wire [BufferCount-1:0] buf_we1;
wire [AddressWidth-1:0] buf_a1_0, buf_a1_1;
wire [DataWidth-1:0] buf_d1_0, buf_d1_1;
//------------------------Instantiation------------------
//genvar i;
        td_fused_top_dataflow_in_loop_TOP_LOOP76_ifmap_vec_0_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP76_ifmap_vec_0_0_memcore_U_0 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_0 ),
            .ce0      ( buf_ce0[ 0 ] ),
            .we0      ( buf_we0[ 0 ] ),
            .d0       ( buf_d0_0 ),
            .q0       ( buf_q0_0 ),
            .address1 ( buf_a1_0 ),
            .ce1      ( buf_ce1[ 0 ] ),
            .we1      ( buf_we1[ 0 ] ),
            .d1       ( buf_d1_0 )
        );
        td_fused_top_dataflow_in_loop_TOP_LOOP76_ifmap_vec_0_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP76_ifmap_vec_0_0_memcore_U_1 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_1 ),
            .ce0      ( buf_ce0[ 1 ] ),
            .we0      ( buf_we0[ 1 ] ),
            .d0       ( buf_d0_1 ),
            .q0       ( buf_q0_1 ),
            .address1 ( buf_a1_1 ),
            .ce1      ( buf_ce1[ 1 ] ),
            .we1      ( buf_we1[ 1 ] ),
            .d1       ( buf_d1_1 )
        );

//++++++++++++++++++++++++buffer signals+++++++++++++++++
        assign buf_ce0[ 0 ] = (tptr ==  0  && empty_n) ? t_ce0
                             : (iptr ==  0 ) ? i_ce0 : 1'b0;
        assign buf_a0_0  = (tptr ==  0  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 0 ] = (tptr ==  0  && empty_n)  ? t_we0
                             : (iptr ==  0 ) ? i_we0 : 1'b0;
        assign buf_d0_0  = (tptr ==  0  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 0 ] = (tptr ==  0  && empty_n) ? t_ce1
                             : (iptr ==  0 ) ? i_ce1 : 1'b0;
        assign buf_a1_0  = (tptr ==  0  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 0 ] = (tptr ==  0  && empty_n)  ? t_we1
                             : (iptr ==  0 ) ? i_we1 : 1'b0;
        assign buf_d1_0  = (tptr ==  0  && empty_n) ? t_d1       : i_d1;
        assign buf_ce0[ 1 ] = (tptr ==  1  && empty_n) ? t_ce0
                             : (iptr ==  1 ) ? i_ce0 : 1'b0;
        assign buf_a0_1  = (tptr ==  1  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 1 ] = (tptr ==  1  && empty_n)  ? t_we0
                             : (iptr ==  1 ) ? i_we0 : 1'b0;
        assign buf_d0_1  = (tptr ==  1  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 1 ] = (tptr ==  1  && empty_n) ? t_ce1
                             : (iptr ==  1 ) ? i_ce1 : 1'b0;
        assign buf_a1_1  = (tptr ==  1  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 1 ] = (tptr ==  1  && empty_n)  ? t_we1
                             : (iptr ==  1 ) ? i_we1 : 1'b0;
        assign buf_d1_1  = (tptr ==  1  && empty_n) ? t_d1       : i_d1;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//------------------------Body---------------------------
assign i_q0      = (prev_iptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign t_q0      = reg_valid0 ? reg_q0 : (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// prev_iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_iptr <= 1'b0;
    else begin
        prev_iptr <= iptr;
    end
end

// prev_tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_tptr <= 1'b0;
    else begin
        prev_tptr <= tptr;
    end
end

// reg_q0 and reg_valid0
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q0     <= 1'b0;
        reg_valid0 <= 1'b0;
    end else if (!t_ce0 && !reg_valid0) begin
        reg_q0     <= (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
        reg_valid0 <= 1'b1;
    end else if (t_ce0) begin
        reg_valid0 <= 1'b0;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP76_products_0_memcore_ram (addr0, ce0, d0, we0, q0, addr1, ce1, q1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
output reg[DWIDTH-1:0] q1;
input clk;

reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];




always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        q1 <= ram[addr1];
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP76_products_0_memcore(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    q0,
    address1,
    ce1,
    q1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
output[DataWidth - 1:0] q1;



td_fused_top_dataflow_in_loop_TOP_LOOP76_products_0_memcore_ram td_fused_top_dataflow_in_loop_TOP_LOOP76_products_0_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .q1( q1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_dataflow_in_loop_TOP_LOOP76_products_0
#(parameter
    DataWidth    = 16,
    AddressRange = 32,
    AddressWidth = 7,
    BufferCount  = 2,
    MemLatency   = 1,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire                    i_we0,
    input  wire [AddressWidth-1:0] i_address0,
    input  wire [DataWidth-1:0]    i_d0,
    output wire [DataWidth-1:0]    i_q0,
    input  wire                    i_ce1,
    input  wire [AddressWidth-1:0] i_address1,
    output wire [DataWidth-1:0]    i_q1,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire                    t_we0,
    input  wire [AddressWidth-1:0] t_address0,
    input  wire [DataWidth-1:0]    t_d0,
    output wire [DataWidth-1:0]    t_q0,
    input  wire                    t_ce1,
    input  wire [AddressWidth-1:0] t_address1,
    output wire [DataWidth-1:0]    t_q1
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth-1:0]   prev_iptr    = 1'b0; // previous initiator index
reg  [IndexWidth-1:0]   prev_tptr    = 1'b0; // previous target index
reg  [DataWidth-1:0]    reg_q0      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid0    = 1'b0; // buffer has valid data
reg  [DataWidth-1:0]    reg_q1      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid1    = 1'b0; // buffer has valid data
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
// buffer signals
wire [BufferCount-1:0] buf_ce0;
wire [BufferCount-1:0] buf_we0;
wire [AddressWidth-1:0] buf_a0_0, buf_a0_1;
wire [DataWidth-1:0] buf_d0_0, buf_d0_1;
wire [DataWidth-1:0] buf_q0_0, buf_q0_1;
wire [BufferCount-1:0] buf_ce1;
wire [AddressWidth-1:0] buf_a1_0, buf_a1_1;
wire [DataWidth-1:0] buf_q1_0, buf_q1_1;
//------------------------Instantiation------------------
//genvar i;
        td_fused_top_dataflow_in_loop_TOP_LOOP76_products_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP76_products_0_memcore_U_0 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_0 ),
            .ce0      ( buf_ce0[ 0 ] ),
            .we0      ( buf_we0[ 0 ] ),
            .d0       ( buf_d0_0 ),
            .q0       ( buf_q0_0 ),
            .address1 ( buf_a1_0 ),
            .ce1      ( buf_ce1[ 0 ] ),
            .q1       ( buf_q1_0 )
        );
        td_fused_top_dataflow_in_loop_TOP_LOOP76_products_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP76_products_0_memcore_U_1 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_1 ),
            .ce0      ( buf_ce0[ 1 ] ),
            .we0      ( buf_we0[ 1 ] ),
            .d0       ( buf_d0_1 ),
            .q0       ( buf_q0_1 ),
            .address1 ( buf_a1_1 ),
            .ce1      ( buf_ce1[ 1 ] ),
            .q1       ( buf_q1_1 )
        );

//++++++++++++++++++++++++buffer signals+++++++++++++++++
        assign buf_ce0[ 0 ] = (tptr ==  0  && empty_n) ? t_ce0
                             : (iptr ==  0 ) ? i_ce0 : 1'b0;
        assign buf_a0_0  = (tptr ==  0  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 0 ] = (tptr ==  0  && empty_n)  ? t_we0
                             : (iptr ==  0 ) ? i_we0 : 1'b0;
        assign buf_d0_0  = (tptr ==  0  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 0 ] = (tptr ==  0  && empty_n) ? t_ce1
                             : (iptr ==  0 ) ? i_ce1 : 1'b0;
        assign buf_a1_0  = (tptr ==  0  && empty_n) ?  t_address1 : i_address1;
        assign buf_ce0[ 1 ] = (tptr ==  1  && empty_n) ? t_ce0
                             : (iptr ==  1 ) ? i_ce0 : 1'b0;
        assign buf_a0_1  = (tptr ==  1  && empty_n) ?  t_address0 : i_address0;
        assign buf_we0[ 1 ] = (tptr ==  1  && empty_n)  ? t_we0
                             : (iptr ==  1 ) ? i_we0 : 1'b0;
        assign buf_d0_1  = (tptr ==  1  && empty_n) ? t_d0       : i_d0;
        assign buf_ce1[ 1 ] = (tptr ==  1  && empty_n) ? t_ce1
                             : (iptr ==  1 ) ? i_ce1 : 1'b0;
        assign buf_a1_1  = (tptr ==  1  && empty_n) ?  t_address1 : i_address1;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//------------------------Body---------------------------
assign i_q0      = (prev_iptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign t_q0      = reg_valid0 ? reg_q0 : (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign i_q1      = (prev_iptr == 1'b1 ? buf_q1_1 : buf_q1_0);
assign t_q1      = reg_valid1 ? reg_q1 : (prev_tptr == 1'b1 ? buf_q1_1 : buf_q1_0);

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// prev_iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_iptr <= 1'b0;
    else begin
        prev_iptr <= iptr;
    end
end

// prev_tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_tptr <= 1'b0;
    else begin
        prev_tptr <= tptr;
    end
end

// reg_q0 and reg_valid0
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q0     <= 1'b0;
        reg_valid0 <= 1'b0;
    end else if (!t_ce0 && !reg_valid0) begin
        reg_q0     <= (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
        reg_valid0 <= 1'b1;
    end else if (t_ce0) begin
        reg_valid0 <= 1'b0;
    end
end

// reg_q1 and reg_valid1
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q1     <= 1'b0;
        reg_valid1 <= 1'b0;
    end else if (!t_ce1 && !reg_valid1) begin
        reg_q1     <= (prev_tptr == 1'b1 ? buf_q1_1 : buf_q1_0);
        reg_valid1 <= 1'b1;
    end else if (t_ce1) begin
        reg_valid1 <= 1'b0;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_dataflow_in_loop_TOP_LOOP76 (
        ap_clk,
        ap_rst,
        in_data_address0,
        in_data_ce0,
        in_data_d0,
        in_data_q0,
        in_data_we0,
        in_data_address1,
        in_data_ce1,
        in_data_d1,
        in_data_q1,
        in_data_we1,
        filter_data_address0,
        filter_data_ce0,
        filter_data_d0,
        filter_data_q0,
        filter_data_we0,
        filter_data_address1,
        filter_data_ce1,
        filter_data_d1,
        filter_data_q1,
        filter_data_we1,
        adjustments_address0,
        adjustments_ce0,
        adjustments_d0,
        adjustments_q0,
        adjustments_we0,
        adjustments_address1,
        adjustments_ce1,
        adjustments_d1,
        adjustments_q1,
        adjustments_we1,
        out_data_address0,
        out_data_ce0,
        out_data_d0,
        out_data_q0,
        out_data_we0,
        out_data_address1,
        out_data_ce1,
        out_data_d1,
        out_data_q1,
        out_data_we1,
        ap_start,
        in_data_empty_n,
        in_data_read,
        out_data_full_n,
        out_data_write,
        ap_done,
        ap_ready,
        ap_idle,
        ap_continue
);


input   ap_clk;
input   ap_rst;
output  [12:0] in_data_address0;
output   in_data_ce0;
output  [63:0] in_data_d0;
input  [63:0] in_data_q0;
output   in_data_we0;
output  [12:0] in_data_address1;
output   in_data_ce1;
output  [63:0] in_data_d1;
input  [63:0] in_data_q1;
output   in_data_we1;
output  [16:0] filter_data_address0;
output   filter_data_ce0;
output  [15:0] filter_data_d0;
input  [15:0] filter_data_q0;
output   filter_data_we0;
output  [16:0] filter_data_address1;
output   filter_data_ce1;
output  [15:0] filter_data_d1;
input  [15:0] filter_data_q1;
output   filter_data_we1;
output  [9:0] adjustments_address0;
output   adjustments_ce0;
output  [47:0] adjustments_d0;
input  [47:0] adjustments_q0;
output   adjustments_we0;
output  [9:0] adjustments_address1;
output   adjustments_ce1;
output  [47:0] adjustments_d1;
input  [47:0] adjustments_q1;
output   adjustments_we1;
output  [15:0] out_data_address0;
output   out_data_ce0;
output  [63:0] out_data_d0;
input  [63:0] out_data_q0;
output   out_data_we0;
output  [15:0] out_data_address1;
output   out_data_ce1;
output  [63:0] out_data_d1;
input  [63:0] out_data_q1;
output   out_data_we1;
input   ap_start;
input   in_data_empty_n;
output   in_data_read;
input   out_data_full_n;
output   out_data_write;
output   ap_done;
output   ap_ready;
output   ap_idle;
input   ap_continue;

wire   [15:0] ifmap_vec_0_0_i_q0;
wire   [15:0] ifmap_vec_0_0_t_q0;
wire   [15:0] weight_vecs_0_0_0_i_q0;
wire   [15:0] weight_vecs_0_0_0_t_q0;
wire   [15:0] products_0_i_q0;
wire   [15:0] products_0_i_q1;
wire   [15:0] products_0_t_q0;
wire   [15:0] products_0_t_q1;
wire   [15:0] accum1_out_0_i_q0;
wire   [15:0] accum1_out_0_t_q0;
wire    tdf12_get_next_ijk_U0_ap_start;
wire    tdf12_get_next_ijk_U0_ap_done;
wire    tdf12_get_next_ijk_U0_ap_continue;
wire    tdf12_get_next_ijk_U0_ap_idle;
wire    tdf12_get_next_ijk_U0_ap_ready;
wire    tdf12_get_next_ijk_U0_start_out;
wire    tdf12_get_next_ijk_U0_start_write;
wire   [15:0] tdf12_get_next_ijk_U0_indices_0_din;
wire    tdf12_get_next_ijk_U0_indices_0_write;
wire   [15:0] tdf12_get_next_ijk_U0_indices_1_din;
wire    tdf12_get_next_ijk_U0_indices_1_write;
wire   [9:0] tdf12_get_next_ijk_U0_indices_2_out_din;
wire    tdf12_get_next_ijk_U0_indices_2_out_write;
wire   [9:0] tdf12_get_next_ijk_U0_indices_2_out1_din;
wire    tdf12_get_next_ijk_U0_indices_2_out1_write;
wire    tdf12_readInputs_U0_ap_start;
wire    tdf12_readInputs_U0_ap_done;
wire    tdf12_readInputs_U0_ap_continue;
wire    tdf12_readInputs_U0_ap_idle;
wire    tdf12_readInputs_U0_ap_ready;
wire   [12:0] tdf12_readInputs_U0_in_data_address0;
wire    tdf12_readInputs_U0_in_data_ce0;
wire    tdf12_readInputs_U0_indices_01_read;
wire    tdf12_readInputs_U0_indices_12_read;
wire   [6:0] tdf12_readInputs_U0_ifmap_vec_0_0_address0;
wire    tdf12_readInputs_U0_ifmap_vec_0_0_ce0;
wire    tdf12_readInputs_U0_ifmap_vec_0_0_we0;
wire   [15:0] tdf12_readInputs_U0_ifmap_vec_0_0_d0;
wire   [6:0] tdf12_readInputs_U0_ifmap_vec_0_0_address1;
wire    tdf12_readInputs_U0_ifmap_vec_0_0_ce1;
wire    tdf12_readInputs_U0_ifmap_vec_0_0_we1;
wire   [15:0] tdf12_readInputs_U0_ifmap_vec_0_0_d1;
wire   [3:0] tdf12_readInputs_U0_indices_01_out_din;
wire    tdf12_readInputs_U0_indices_01_out_write;
wire   [7:0] tdf12_readInputs_U0_indices_12_out_din;
wire    tdf12_readInputs_U0_indices_12_out_write;
wire    tdf12_readInputs_U0_in_data_full_n;
wire    tdf12_readInputs_U0_in_data_write;
wire    ap_channel_done_ifmap_vec_0_0;
wire    tdf12_readInputs_U0_ifmap_vec_0_0_full_n;
wire    tdf12_readFilters78_U0_ap_start;
wire    tdf12_readFilters78_U0_ap_done;
wire    tdf12_readFilters78_U0_ap_continue;
wire    tdf12_readFilters78_U0_ap_idle;
wire    tdf12_readFilters78_U0_ap_ready;
wire   [16:0] tdf12_readFilters78_U0_filter_data_address0;
wire    tdf12_readFilters78_U0_filter_data_ce0;
wire    tdf12_readFilters78_U0_indices_23_read;
wire   [6:0] tdf12_readFilters78_U0_weight_vecs_0_0_0_address0;
wire    tdf12_readFilters78_U0_weight_vecs_0_0_0_ce0;
wire    tdf12_readFilters78_U0_weight_vecs_0_0_0_we0;
wire   [15:0] tdf12_readFilters78_U0_weight_vecs_0_0_0_d0;
wire    ap_channel_done_weight_vecs_0_0_0;
wire    tdf12_readFilters78_U0_weight_vecs_0_0_0_full_n;
wire    tdf12_dot_product_U0_ap_start;
wire    tdf12_dot_product_U0_ap_done;
wire    tdf12_dot_product_U0_ap_continue;
wire    tdf12_dot_product_U0_ap_idle;
wire    tdf12_dot_product_U0_ap_ready;
wire   [6:0] tdf12_dot_product_U0_ifmap_vec_0_0_address0;
wire    tdf12_dot_product_U0_ifmap_vec_0_0_ce0;
wire   [6:0] tdf12_dot_product_U0_weight_vecs_0_0_0_address0;
wire    tdf12_dot_product_U0_weight_vecs_0_0_0_ce0;
wire   [6:0] tdf12_dot_product_U0_products_0_address0;
wire    tdf12_dot_product_U0_products_0_ce0;
wire    tdf12_dot_product_U0_products_0_we0;
wire   [15:0] tdf12_dot_product_U0_products_0_d0;
wire    ap_channel_done_products_0;
wire    tdf12_dot_product_U0_products_0_full_n;
wire    tdf12_accum_1_U0_ap_start;
wire    tdf12_accum_1_U0_ap_done;
wire    tdf12_accum_1_U0_ap_continue;
wire    tdf12_accum_1_U0_ap_idle;
wire    tdf12_accum_1_U0_ap_ready;
wire   [6:0] tdf12_accum_1_U0_accum_in_0_address0;
wire    tdf12_accum_1_U0_accum_in_0_ce0;
wire   [6:0] tdf12_accum_1_U0_accum_in_0_address1;
wire    tdf12_accum_1_U0_accum_in_0_ce1;
wire   [2:0] tdf12_accum_1_U0_accum_out_address0;
wire    tdf12_accum_1_U0_accum_out_ce0;
wire    tdf12_accum_1_U0_accum_out_we0;
wire   [15:0] tdf12_accum_1_U0_accum_out_d0;
wire   [2:0] tdf12_accum_1_U0_accum_out_address1;
wire    tdf12_accum_1_U0_accum_out_ce1;
wire    tdf12_accum_1_U0_accum_out_we1;
wire   [15:0] tdf12_accum_1_U0_accum_out_d1;
wire    ap_channel_done_accum1_out_0;
wire    tdf12_accum_1_U0_accum_out_full_n;
wire    tdf12_accum_2_U0_ap_start;
wire    tdf12_accum_2_U0_ap_done;
wire    tdf12_accum_2_U0_ap_continue;
wire    tdf12_accum_2_U0_ap_idle;
wire    tdf12_accum_2_U0_ap_ready;
wire   [15:0] tdf12_accum_2_U0_accum_in_20;
wire    tdf12_accum_2_U0_accum_in_20_ap_vld;
wire   [2:0] tdf12_accum_2_U0_accum_in_address0;
wire    tdf12_accum_2_U0_accum_in_ce0;
wire    ap_channel_done_tmp_channel;
wire    tmp_channel_full_n;
wire    Block_entry_proc_proc446_U0_ap_start;
wire    Block_entry_proc_proc446_U0_ap_done;
wire    Block_entry_proc_proc446_U0_ap_continue;
wire    Block_entry_proc_proc446_U0_ap_idle;
wire    Block_entry_proc_proc446_U0_ap_ready;
wire   [15:0] Block_entry_proc_proc446_U0_ap_return;
wire    ap_channel_done_sums_0;
wire    sums_0_full_n;
wire    tdf12_adjust_U0_ap_start;
wire    tdf12_adjust_U0_ap_done;
wire    tdf12_adjust_U0_ap_continue;
wire    tdf12_adjust_U0_ap_idle;
wire    tdf12_adjust_U0_ap_ready;
wire   [9:0] tdf12_adjust_U0_adjustments_address0;
wire    tdf12_adjust_U0_adjustments_ce0;
wire    tdf12_adjust_U0_indices_23_read;
wire   [15:0] tdf12_adjust_U0_ap_return;
wire    ap_channel_done_outputs_0;
wire    outputs_0_full_n;
wire    tdf12_writeOutputs_unaligned_U0_ap_start;
wire    tdf12_writeOutputs_unaligned_U0_ap_done;
wire    tdf12_writeOutputs_unaligned_U0_ap_continue;
wire    tdf12_writeOutputs_unaligned_U0_ap_idle;
wire    tdf12_writeOutputs_unaligned_U0_ap_ready;
wire    tdf12_writeOutputs_unaligned_U0_indices_01_read;
wire    tdf12_writeOutputs_unaligned_U0_indices_12_read;
wire   [15:0] tdf12_writeOutputs_unaligned_U0_out_data_address1;
wire    tdf12_writeOutputs_unaligned_U0_out_data_ce1;
wire    tdf12_writeOutputs_unaligned_U0_out_data_we1;
wire   [63:0] tdf12_writeOutputs_unaligned_U0_out_data_d1;
wire    tdf12_writeOutputs_unaligned_U0_out_data_full_n;
wire    tdf12_writeOutputs_unaligned_U0_out_data_write;
wire    ap_sync_continue;
wire    ifmap_vec_0_0_i_full_n;
wire    ifmap_vec_0_0_t_empty_n;
wire    weight_vecs_0_0_0_i_full_n;
wire    weight_vecs_0_0_0_t_empty_n;
wire    products_0_i_full_n;
wire    products_0_t_empty_n;
wire   [15:0] products_0_t_d1;
wire    products_0_t_we1;
wire    accum1_out_0_i_full_n;
wire    accum1_out_0_t_empty_n;
wire    indices_01_c_full_n;
wire   [15:0] indices_01_c_dout;
wire    indices_01_c_empty_n;
wire    indices_12_c_full_n;
wire   [15:0] indices_12_c_dout;
wire    indices_12_c_empty_n;
wire    indices_23_c_full_n;
wire   [9:0] indices_23_c_dout;
wire    indices_23_c_empty_n;
wire    indices_23_c1_full_n;
wire   [9:0] indices_23_c1_dout;
wire    indices_23_c1_empty_n;
wire    indices_01_c2_full_n;
wire   [3:0] indices_01_c2_dout;
wire    indices_01_c2_empty_n;
wire    indices_12_c3_full_n;
wire   [7:0] indices_12_c3_dout;
wire    indices_12_c3_empty_n;
wire   [15:0] tmp_channel_dout;
wire    tmp_channel_empty_n;
wire   [15:0] sums_0_dout;
wire    sums_0_empty_n;
wire   [15:0] outputs_0_dout;
wire    outputs_0_empty_n;
wire    ap_sync_done;
wire    ap_sync_ready;
reg    ap_sync_reg_tdf12_get_next_ijk_U0_ap_ready;
wire    ap_sync_tdf12_get_next_ijk_U0_ap_ready;
reg    ap_sync_reg_tdf12_readInputs_U0_ap_ready;
wire    ap_sync_tdf12_readInputs_U0_ap_ready;
wire   [0:0] start_for_tdf12_readFilters78_U0_din;
wire    start_for_tdf12_readFilters78_U0_full_n;
wire   [0:0] start_for_tdf12_readFilters78_U0_dout;
wire    start_for_tdf12_readFilters78_U0_empty_n;
wire    tdf12_readInputs_U0_start_full_n;
wire    tdf12_readInputs_U0_start_write;
wire    tdf12_readFilters78_U0_start_full_n;
wire    tdf12_readFilters78_U0_start_write;
wire    tdf12_dot_product_U0_start_full_n;
wire    tdf12_dot_product_U0_start_write;
wire    tdf12_accum_1_U0_start_full_n;
wire    tdf12_accum_1_U0_start_write;
wire    tdf12_accum_2_U0_start_full_n;
wire    tdf12_accum_2_U0_start_write;
wire    Block_entry_proc_proc446_U0_start_full_n;
wire    Block_entry_proc_proc446_U0_start_write;
wire    tdf12_adjust_U0_start_full_n;
wire    tdf12_adjust_U0_start_write;
wire    tdf12_writeOutputs_unaligned_U0_start_full_n;
wire    tdf12_writeOutputs_unaligned_U0_start_write;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_sync_reg_tdf12_get_next_ijk_U0_ap_ready = 1'b0;
#0 ap_sync_reg_tdf12_readInputs_U0_ap_ready = 1'b0;
end

td_fused_top_dataflow_in_loop_TOP_LOOP76_ifmap_vec_0_0 #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
ifmap_vec_0_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf12_readInputs_U0_ap_done),
    .i_full_n(ifmap_vec_0_0_i_full_n),
    .i_ce0(tdf12_readInputs_U0_ifmap_vec_0_0_ce0),
    .i_we0(tdf12_readInputs_U0_ifmap_vec_0_0_we0),
    .i_address0(tdf12_readInputs_U0_ifmap_vec_0_0_address0),
    .i_d0(tdf12_readInputs_U0_ifmap_vec_0_0_d0),
    .i_q0(ifmap_vec_0_0_i_q0),
    .i_ce1(tdf12_readInputs_U0_ifmap_vec_0_0_ce1),
    .i_we1(tdf12_readInputs_U0_ifmap_vec_0_0_we1),
    .i_address1(tdf12_readInputs_U0_ifmap_vec_0_0_address1),
    .i_d1(tdf12_readInputs_U0_ifmap_vec_0_0_d1),
    .t_ce(1'b1),
    .t_read(tdf12_dot_product_U0_ap_ready),
    .t_empty_n(ifmap_vec_0_0_t_empty_n),
    .t_ce0(tdf12_dot_product_U0_ifmap_vec_0_0_ce0),
    .t_we0(1'b0),
    .t_address0(tdf12_dot_product_U0_ifmap_vec_0_0_address0),
    .t_d0(16'd0),
    .t_q0(ifmap_vec_0_0_t_q0),
    .t_ce1(1'b0),
    .t_we1(1'b0),
    .t_address1(7'd0),
    .t_d1(16'd0)
);

td_fused_top_dataflow_in_loop_TOP_LOOP76_weight_vecs_0_0_0 #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
weight_vecs_0_0_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf12_readFilters78_U0_ap_done),
    .i_full_n(weight_vecs_0_0_0_i_full_n),
    .i_ce0(tdf12_readFilters78_U0_weight_vecs_0_0_0_ce0),
    .i_we0(tdf12_readFilters78_U0_weight_vecs_0_0_0_we0),
    .i_address0(tdf12_readFilters78_U0_weight_vecs_0_0_0_address0),
    .i_d0(tdf12_readFilters78_U0_weight_vecs_0_0_0_d0),
    .i_q0(weight_vecs_0_0_0_i_q0),
    .t_ce(1'b1),
    .t_read(tdf12_dot_product_U0_ap_ready),
    .t_empty_n(weight_vecs_0_0_0_t_empty_n),
    .t_ce0(tdf12_dot_product_U0_weight_vecs_0_0_0_ce0),
    .t_we0(1'b0),
    .t_address0(tdf12_dot_product_U0_weight_vecs_0_0_0_address0),
    .t_d0(16'd0),
    .t_q0(weight_vecs_0_0_0_t_q0)
);

td_fused_top_dataflow_in_loop_TOP_LOOP76_products_0 #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
products_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf12_dot_product_U0_ap_done),
    .i_full_n(products_0_i_full_n),
    .i_ce0(tdf12_dot_product_U0_products_0_ce0),
    .i_we0(tdf12_dot_product_U0_products_0_we0),
    .i_address0(tdf12_dot_product_U0_products_0_address0),
    .i_d0(tdf12_dot_product_U0_products_0_d0),
    .i_q0(products_0_i_q0),
    .i_ce1(1'b0),
    .i_address1(7'd0),
    .i_q1(products_0_i_q1),
    .t_ce(1'b1),
    .t_read(tdf12_accum_1_U0_ap_ready),
    .t_empty_n(products_0_t_empty_n),
    .t_ce0(tdf12_accum_1_U0_accum_in_0_ce0),
    .t_we0(1'b0),
    .t_address0(tdf12_accum_1_U0_accum_in_0_address0),
    .t_d0(16'd0),
    .t_q0(products_0_t_q0),
    .t_ce1(tdf12_accum_1_U0_accum_in_0_ce1),
    .t_address1(tdf12_accum_1_U0_accum_in_0_address1),
    .t_q1(products_0_t_q1)
);

td_fused_top_dataflow_in_loop_TOP_LOOP76_accum1_out_0 #(
    .DataWidth( 16 ),
    .AddressRange( 8 ),
    .AddressWidth( 3 ))
accum1_out_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf12_accum_1_U0_ap_done),
    .i_full_n(accum1_out_0_i_full_n),
    .i_ce0(tdf12_accum_1_U0_accum_out_ce0),
    .i_we0(tdf12_accum_1_U0_accum_out_we0),
    .i_address0(tdf12_accum_1_U0_accum_out_address0),
    .i_d0(tdf12_accum_1_U0_accum_out_d0),
    .i_q0(accum1_out_0_i_q0),
    .i_ce1(tdf12_accum_1_U0_accum_out_ce1),
    .i_we1(tdf12_accum_1_U0_accum_out_we1),
    .i_address1(tdf12_accum_1_U0_accum_out_address1),
    .i_d1(tdf12_accum_1_U0_accum_out_d1),
    .t_ce(1'b1),
    .t_read(tdf12_accum_2_U0_ap_ready),
    .t_empty_n(accum1_out_0_t_empty_n),
    .t_ce0(tdf12_accum_2_U0_accum_in_ce0),
    .t_we0(1'b0),
    .t_address0(tdf12_accum_2_U0_accum_in_address0),
    .t_d0(16'd0),
    .t_q0(accum1_out_0_t_q0),
    .t_ce1(1'b0),
    .t_we1(1'b0),
    .t_address1(3'd0),
    .t_d1(16'd0)
);

td_fused_top_tdf12_get_next_ijk tdf12_get_next_ijk_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf12_get_next_ijk_U0_ap_start),
    .start_full_n(start_for_tdf12_readFilters78_U0_full_n),
    .ap_done(tdf12_get_next_ijk_U0_ap_done),
    .ap_continue(tdf12_get_next_ijk_U0_ap_continue),
    .ap_idle(tdf12_get_next_ijk_U0_ap_idle),
    .ap_ready(tdf12_get_next_ijk_U0_ap_ready),
    .start_out(tdf12_get_next_ijk_U0_start_out),
    .start_write(tdf12_get_next_ijk_U0_start_write),
    .indices_0_din(tdf12_get_next_ijk_U0_indices_0_din),
    .indices_0_full_n(indices_01_c_full_n),
    .indices_0_write(tdf12_get_next_ijk_U0_indices_0_write),
    .indices_1_din(tdf12_get_next_ijk_U0_indices_1_din),
    .indices_1_full_n(indices_12_c_full_n),
    .indices_1_write(tdf12_get_next_ijk_U0_indices_1_write),
    .indices_2_out_din(tdf12_get_next_ijk_U0_indices_2_out_din),
    .indices_2_out_full_n(indices_23_c_full_n),
    .indices_2_out_write(tdf12_get_next_ijk_U0_indices_2_out_write),
    .indices_2_out1_din(tdf12_get_next_ijk_U0_indices_2_out1_din),
    .indices_2_out1_full_n(indices_23_c1_full_n),
    .indices_2_out1_write(tdf12_get_next_ijk_U0_indices_2_out1_write)
);

td_fused_top_tdf12_readInputs tdf12_readInputs_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf12_readInputs_U0_ap_start),
    .ap_done(tdf12_readInputs_U0_ap_done),
    .ap_continue(tdf12_readInputs_U0_ap_continue),
    .ap_idle(tdf12_readInputs_U0_ap_idle),
    .ap_ready(tdf12_readInputs_U0_ap_ready),
    .in_data_address0(tdf12_readInputs_U0_in_data_address0),
    .in_data_ce0(tdf12_readInputs_U0_in_data_ce0),
    .in_data_q0(in_data_q0),
    .indices_01_dout(indices_01_c_dout),
    .indices_01_empty_n(indices_01_c_empty_n),
    .indices_01_read(tdf12_readInputs_U0_indices_01_read),
    .indices_12_dout(indices_12_c_dout),
    .indices_12_empty_n(indices_12_c_empty_n),
    .indices_12_read(tdf12_readInputs_U0_indices_12_read),
    .ifmap_vec_0_0_address0(tdf12_readInputs_U0_ifmap_vec_0_0_address0),
    .ifmap_vec_0_0_ce0(tdf12_readInputs_U0_ifmap_vec_0_0_ce0),
    .ifmap_vec_0_0_we0(tdf12_readInputs_U0_ifmap_vec_0_0_we0),
    .ifmap_vec_0_0_d0(tdf12_readInputs_U0_ifmap_vec_0_0_d0),
    .ifmap_vec_0_0_address1(tdf12_readInputs_U0_ifmap_vec_0_0_address1),
    .ifmap_vec_0_0_ce1(tdf12_readInputs_U0_ifmap_vec_0_0_ce1),
    .ifmap_vec_0_0_we1(tdf12_readInputs_U0_ifmap_vec_0_0_we1),
    .ifmap_vec_0_0_d1(tdf12_readInputs_U0_ifmap_vec_0_0_d1),
    .indices_01_out_din(tdf12_readInputs_U0_indices_01_out_din),
    .indices_01_out_full_n(indices_01_c2_full_n),
    .indices_01_out_write(tdf12_readInputs_U0_indices_01_out_write),
    .indices_12_out_din(tdf12_readInputs_U0_indices_12_out_din),
    .indices_12_out_full_n(indices_12_c3_full_n),
    .indices_12_out_write(tdf12_readInputs_U0_indices_12_out_write)
);

td_fused_top_tdf12_readFilters78 tdf12_readFilters78_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf12_readFilters78_U0_ap_start),
    .ap_done(tdf12_readFilters78_U0_ap_done),
    .ap_continue(tdf12_readFilters78_U0_ap_continue),
    .ap_idle(tdf12_readFilters78_U0_ap_idle),
    .ap_ready(tdf12_readFilters78_U0_ap_ready),
    .filter_data_address0(tdf12_readFilters78_U0_filter_data_address0),
    .filter_data_ce0(tdf12_readFilters78_U0_filter_data_ce0),
    .filter_data_q0(filter_data_q0),
    .indices_23_dout(indices_23_c_dout),
    .indices_23_empty_n(indices_23_c_empty_n),
    .indices_23_read(tdf12_readFilters78_U0_indices_23_read),
    .weight_vecs_0_0_0_address0(tdf12_readFilters78_U0_weight_vecs_0_0_0_address0),
    .weight_vecs_0_0_0_ce0(tdf12_readFilters78_U0_weight_vecs_0_0_0_ce0),
    .weight_vecs_0_0_0_we0(tdf12_readFilters78_U0_weight_vecs_0_0_0_we0),
    .weight_vecs_0_0_0_d0(tdf12_readFilters78_U0_weight_vecs_0_0_0_d0)
);

td_fused_top_tdf12_dot_product tdf12_dot_product_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf12_dot_product_U0_ap_start),
    .ap_done(tdf12_dot_product_U0_ap_done),
    .ap_continue(tdf12_dot_product_U0_ap_continue),
    .ap_idle(tdf12_dot_product_U0_ap_idle),
    .ap_ready(tdf12_dot_product_U0_ap_ready),
    .ifmap_vec_0_0_address0(tdf12_dot_product_U0_ifmap_vec_0_0_address0),
    .ifmap_vec_0_0_ce0(tdf12_dot_product_U0_ifmap_vec_0_0_ce0),
    .ifmap_vec_0_0_q0(ifmap_vec_0_0_t_q0),
    .weight_vecs_0_0_0_address0(tdf12_dot_product_U0_weight_vecs_0_0_0_address0),
    .weight_vecs_0_0_0_ce0(tdf12_dot_product_U0_weight_vecs_0_0_0_ce0),
    .weight_vecs_0_0_0_q0(weight_vecs_0_0_0_t_q0),
    .products_0_address0(tdf12_dot_product_U0_products_0_address0),
    .products_0_ce0(tdf12_dot_product_U0_products_0_ce0),
    .products_0_we0(tdf12_dot_product_U0_products_0_we0),
    .products_0_d0(tdf12_dot_product_U0_products_0_d0)
);

td_fused_top_tdf12_accum_1 tdf12_accum_1_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf12_accum_1_U0_ap_start),
    .ap_done(tdf12_accum_1_U0_ap_done),
    .ap_continue(tdf12_accum_1_U0_ap_continue),
    .ap_idle(tdf12_accum_1_U0_ap_idle),
    .ap_ready(tdf12_accum_1_U0_ap_ready),
    .accum_in_0_address0(tdf12_accum_1_U0_accum_in_0_address0),
    .accum_in_0_ce0(tdf12_accum_1_U0_accum_in_0_ce0),
    .accum_in_0_q0(products_0_t_q0),
    .accum_in_0_address1(tdf12_accum_1_U0_accum_in_0_address1),
    .accum_in_0_ce1(tdf12_accum_1_U0_accum_in_0_ce1),
    .accum_in_0_q1(products_0_t_q1),
    .accum_out_address0(tdf12_accum_1_U0_accum_out_address0),
    .accum_out_ce0(tdf12_accum_1_U0_accum_out_ce0),
    .accum_out_we0(tdf12_accum_1_U0_accum_out_we0),
    .accum_out_d0(tdf12_accum_1_U0_accum_out_d0),
    .accum_out_address1(tdf12_accum_1_U0_accum_out_address1),
    .accum_out_ce1(tdf12_accum_1_U0_accum_out_ce1),
    .accum_out_we1(tdf12_accum_1_U0_accum_out_we1),
    .accum_out_d1(tdf12_accum_1_U0_accum_out_d1)
);

td_fused_top_tdf12_accum_2 tdf12_accum_2_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf12_accum_2_U0_ap_start),
    .ap_done(tdf12_accum_2_U0_ap_done),
    .ap_continue(tdf12_accum_2_U0_ap_continue),
    .ap_idle(tdf12_accum_2_U0_ap_idle),
    .ap_ready(tdf12_accum_2_U0_ap_ready),
    .accum_in_20(tdf12_accum_2_U0_accum_in_20),
    .accum_in_20_ap_vld(tdf12_accum_2_U0_accum_in_20_ap_vld),
    .accum_in_address0(tdf12_accum_2_U0_accum_in_address0),
    .accum_in_ce0(tdf12_accum_2_U0_accum_in_ce0),
    .accum_in_q0(accum1_out_0_t_q0)
);

td_fused_top_Block_entry_proc_proc446 Block_entry_proc_proc446_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(Block_entry_proc_proc446_U0_ap_start),
    .ap_done(Block_entry_proc_proc446_U0_ap_done),
    .ap_continue(Block_entry_proc_proc446_U0_ap_continue),
    .ap_idle(Block_entry_proc_proc446_U0_ap_idle),
    .ap_ready(Block_entry_proc_proc446_U0_ap_ready),
    .tmp(tmp_channel_dout),
    .ap_return(Block_entry_proc_proc446_U0_ap_return)
);

td_fused_top_tdf12_adjust tdf12_adjust_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf12_adjust_U0_ap_start),
    .ap_done(tdf12_adjust_U0_ap_done),
    .ap_continue(tdf12_adjust_U0_ap_continue),
    .ap_idle(tdf12_adjust_U0_ap_idle),
    .ap_ready(tdf12_adjust_U0_ap_ready),
    .sums_read(sums_0_dout),
    .adjustments_address0(tdf12_adjust_U0_adjustments_address0),
    .adjustments_ce0(tdf12_adjust_U0_adjustments_ce0),
    .adjustments_q0(adjustments_q0),
    .indices_23_dout(indices_23_c1_dout),
    .indices_23_empty_n(indices_23_c1_empty_n),
    .indices_23_read(tdf12_adjust_U0_indices_23_read),
    .ap_return(tdf12_adjust_U0_ap_return)
);

td_fused_top_tdf12_writeOutputs_unaligned tdf12_writeOutputs_unaligned_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(tdf12_writeOutputs_unaligned_U0_ap_start),
    .ap_done(tdf12_writeOutputs_unaligned_U0_ap_done),
    .ap_continue(tdf12_writeOutputs_unaligned_U0_ap_continue),
    .ap_idle(tdf12_writeOutputs_unaligned_U0_ap_idle),
    .ap_ready(tdf12_writeOutputs_unaligned_U0_ap_ready),
    .indices_01_dout(indices_01_c2_dout),
    .indices_01_empty_n(indices_01_c2_empty_n),
    .indices_01_read(tdf12_writeOutputs_unaligned_U0_indices_01_read),
    .indices_12_dout(indices_12_c3_dout),
    .indices_12_empty_n(indices_12_c3_empty_n),
    .indices_12_read(tdf12_writeOutputs_unaligned_U0_indices_12_read),
    .p_read(outputs_0_dout),
    .out_data_address1(tdf12_writeOutputs_unaligned_U0_out_data_address1),
    .out_data_ce1(tdf12_writeOutputs_unaligned_U0_out_data_ce1),
    .out_data_we1(tdf12_writeOutputs_unaligned_U0_out_data_we1),
    .out_data_d1(tdf12_writeOutputs_unaligned_U0_out_data_d1)
);

td_fused_top_fifo_w16_d2_S_x9 indices_01_c_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(indices_01_c_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf12_readInputs_U0_indices_01_read),
    .if_dout(indices_01_c_dout),
    .if_full_n(indices_01_c_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf12_get_next_ijk_U0_indices_0_write),
    .if_din(tdf12_get_next_ijk_U0_indices_0_din)
);

td_fused_top_fifo_w16_d2_S_x9 indices_12_c_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(indices_12_c_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf12_readInputs_U0_indices_12_read),
    .if_dout(indices_12_c_dout),
    .if_full_n(indices_12_c_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf12_get_next_ijk_U0_indices_1_write),
    .if_din(tdf12_get_next_ijk_U0_indices_1_din)
);

td_fused_top_fifo_w10_d2_S indices_23_c_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(indices_23_c_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf12_readFilters78_U0_indices_23_read),
    .if_dout(indices_23_c_dout),
    .if_full_n(indices_23_c_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf12_get_next_ijk_U0_indices_2_out_write),
    .if_din(tdf12_get_next_ijk_U0_indices_2_out_din)
);

td_fused_top_fifo_w10_d7_S_x indices_23_c1_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(indices_23_c1_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf12_adjust_U0_indices_23_read),
    .if_dout(indices_23_c1_dout),
    .if_full_n(indices_23_c1_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf12_get_next_ijk_U0_indices_2_out1_write),
    .if_din(tdf12_get_next_ijk_U0_indices_2_out1_din)
);

td_fused_top_fifo_w4_d7_S_x0 indices_01_c2_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(indices_01_c2_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf12_writeOutputs_unaligned_U0_indices_01_read),
    .if_dout(indices_01_c2_dout),
    .if_full_n(indices_01_c2_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf12_readInputs_U0_indices_01_out_write),
    .if_din(tdf12_readInputs_U0_indices_01_out_din)
);

td_fused_top_fifo_w8_d7_S_x0 indices_12_c3_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(indices_12_c3_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf12_writeOutputs_unaligned_U0_indices_12_read),
    .if_dout(indices_12_c3_dout),
    .if_full_n(indices_12_c3_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf12_readInputs_U0_indices_12_out_write),
    .if_din(tdf12_readInputs_U0_indices_12_out_din)
);

td_fused_top_fifo_w16_d2_S_x9 tmp_channel_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(tmp_channel_empty_n),
    .if_read_ce(1'b1),
    .if_read(Block_entry_proc_proc446_U0_ap_ready),
    .if_dout(tmp_channel_dout),
    .if_full_n(tmp_channel_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf12_accum_2_U0_ap_done),
    .if_din(tdf12_accum_2_U0_accum_in_20)
);

td_fused_top_fifo_w16_d2_S_x9 sums_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(sums_0_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf12_adjust_U0_ap_ready),
    .if_dout(sums_0_dout),
    .if_full_n(sums_0_full_n),
    .if_write_ce(1'b1),
    .if_write(Block_entry_proc_proc446_U0_ap_done),
    .if_din(Block_entry_proc_proc446_U0_ap_return)
);

td_fused_top_fifo_w16_d2_S_x9 outputs_0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(outputs_0_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf12_writeOutputs_unaligned_U0_ap_ready),
    .if_dout(outputs_0_dout),
    .if_full_n(outputs_0_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf12_adjust_U0_ap_done),
    .if_din(tdf12_adjust_U0_ap_return)
);

td_fused_top_start_for_tdf12_readFilters78_U0 start_for_tdf12_readFilters78_U0_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .if_empty_n(start_for_tdf12_readFilters78_U0_empty_n),
    .if_read_ce(1'b1),
    .if_read(tdf12_readFilters78_U0_ap_ready),
    .if_dout(start_for_tdf12_readFilters78_U0_dout),
    .if_full_n(start_for_tdf12_readFilters78_U0_full_n),
    .if_write_ce(1'b1),
    .if_write(tdf12_get_next_ijk_U0_start_write),
    .if_din(start_for_tdf12_readFilters78_U0_din)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_sync_reg_tdf12_get_next_ijk_U0_ap_ready <= 1'b0;
    end else begin
        if (((ap_sync_ready & ap_start) == 1'b1)) begin
            ap_sync_reg_tdf12_get_next_ijk_U0_ap_ready <= 1'b0;
        end else begin
            ap_sync_reg_tdf12_get_next_ijk_U0_ap_ready <= ap_sync_tdf12_get_next_ijk_U0_ap_ready;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_sync_reg_tdf12_readInputs_U0_ap_ready <= 1'b0;
    end else begin
        if (((ap_sync_ready & ap_start) == 1'b1)) begin
            ap_sync_reg_tdf12_readInputs_U0_ap_ready <= 1'b0;
        end else begin
            ap_sync_reg_tdf12_readInputs_U0_ap_ready <= ap_sync_tdf12_readInputs_U0_ap_ready;
        end
    end
end

assign Block_entry_proc_proc446_U0_ap_continue = sums_0_full_n;

assign Block_entry_proc_proc446_U0_ap_start = tmp_channel_empty_n;

assign Block_entry_proc_proc446_U0_start_full_n = 1'b1;

assign Block_entry_proc_proc446_U0_start_write = 1'b0;

assign adjustments_address0 = tdf12_adjust_U0_adjustments_address0;

assign adjustments_address1 = 10'd0;

assign adjustments_ce0 = tdf12_adjust_U0_adjustments_ce0;

assign adjustments_ce1 = 1'b0;

assign adjustments_d0 = 48'd0;

assign adjustments_d1 = 48'd0;

assign adjustments_we0 = 1'b0;

assign adjustments_we1 = 1'b0;

assign ap_channel_done_accum1_out_0 = tdf12_accum_1_U0_ap_done;

assign ap_channel_done_ifmap_vec_0_0 = tdf12_readInputs_U0_ap_done;

assign ap_channel_done_outputs_0 = tdf12_adjust_U0_ap_done;

assign ap_channel_done_products_0 = tdf12_dot_product_U0_ap_done;

assign ap_channel_done_sums_0 = Block_entry_proc_proc446_U0_ap_done;

assign ap_channel_done_tmp_channel = tdf12_accum_2_U0_ap_done;

assign ap_channel_done_weight_vecs_0_0_0 = tdf12_readFilters78_U0_ap_done;

assign ap_done = tdf12_writeOutputs_unaligned_U0_ap_done;

assign ap_idle = (tdf12_writeOutputs_unaligned_U0_ap_idle & tdf12_readInputs_U0_ap_idle & tdf12_readFilters78_U0_ap_idle & tdf12_get_next_ijk_U0_ap_idle & tdf12_dot_product_U0_ap_idle & tdf12_adjust_U0_ap_idle & tdf12_accum_2_U0_ap_idle & tdf12_accum_1_U0_ap_idle & (outputs_0_empty_n ^ 1'b1) & (sums_0_empty_n ^ 1'b1) & (tmp_channel_empty_n ^ 1'b1) & (products_0_t_empty_n ^ 1'b1) & (weight_vecs_0_0_0_t_empty_n ^ 1'b1) & (ifmap_vec_0_0_t_empty_n ^ 1'b1) & (1'b1 ^ accum1_out_0_t_empty_n) & Block_entry_proc_proc446_U0_ap_idle);

assign ap_ready = ap_sync_ready;

assign ap_sync_continue = ap_continue;

assign ap_sync_done = tdf12_writeOutputs_unaligned_U0_ap_done;

assign ap_sync_ready = (ap_sync_tdf12_readInputs_U0_ap_ready & ap_sync_tdf12_get_next_ijk_U0_ap_ready);

assign ap_sync_tdf12_get_next_ijk_U0_ap_ready = (tdf12_get_next_ijk_U0_ap_ready | ap_sync_reg_tdf12_get_next_ijk_U0_ap_ready);

assign ap_sync_tdf12_readInputs_U0_ap_ready = (tdf12_readInputs_U0_ap_ready | ap_sync_reg_tdf12_readInputs_U0_ap_ready);

assign filter_data_address0 = tdf12_readFilters78_U0_filter_data_address0;

assign filter_data_address1 = 17'd0;

assign filter_data_ce0 = tdf12_readFilters78_U0_filter_data_ce0;

assign filter_data_ce1 = 1'b0;

assign filter_data_d0 = 16'd0;

assign filter_data_d1 = 16'd0;

assign filter_data_we0 = 1'b0;

assign filter_data_we1 = 1'b0;

assign in_data_address0 = tdf12_readInputs_U0_in_data_address0;

assign in_data_address1 = 13'd0;

assign in_data_ce0 = tdf12_readInputs_U0_in_data_ce0;

assign in_data_ce1 = 1'b0;

assign in_data_d0 = 64'd0;

assign in_data_d1 = 64'd0;

assign in_data_read = tdf12_readInputs_U0_in_data_write;

assign in_data_we0 = 1'b0;

assign in_data_we1 = 1'b0;

assign out_data_address0 = 16'd0;

assign out_data_address1 = tdf12_writeOutputs_unaligned_U0_out_data_address1;

assign out_data_ce0 = 1'b0;

assign out_data_ce1 = tdf12_writeOutputs_unaligned_U0_out_data_ce1;

assign out_data_d0 = 64'd0;

assign out_data_d1 = tdf12_writeOutputs_unaligned_U0_out_data_d1;

assign out_data_we0 = 1'b0;

assign out_data_we1 = tdf12_writeOutputs_unaligned_U0_out_data_we1;

assign out_data_write = tdf12_writeOutputs_unaligned_U0_out_data_write;

assign products_0_t_d1 = 16'd0;

assign products_0_t_we1 = 1'b0;

assign start_for_tdf12_readFilters78_U0_din = 1'b1;

assign tdf12_accum_1_U0_accum_out_full_n = accum1_out_0_i_full_n;

assign tdf12_accum_1_U0_ap_continue = accum1_out_0_i_full_n;

assign tdf12_accum_1_U0_ap_start = products_0_t_empty_n;

assign tdf12_accum_1_U0_start_full_n = 1'b1;

assign tdf12_accum_1_U0_start_write = 1'b0;

assign tdf12_accum_2_U0_ap_continue = tmp_channel_full_n;

assign tdf12_accum_2_U0_ap_start = accum1_out_0_t_empty_n;

assign tdf12_accum_2_U0_start_full_n = 1'b1;

assign tdf12_accum_2_U0_start_write = 1'b0;

assign tdf12_adjust_U0_ap_continue = outputs_0_full_n;

assign tdf12_adjust_U0_ap_start = sums_0_empty_n;

assign tdf12_adjust_U0_start_full_n = 1'b1;

assign tdf12_adjust_U0_start_write = 1'b0;

assign tdf12_dot_product_U0_ap_continue = products_0_i_full_n;

assign tdf12_dot_product_U0_ap_start = (weight_vecs_0_0_0_t_empty_n & ifmap_vec_0_0_t_empty_n);

assign tdf12_dot_product_U0_products_0_full_n = products_0_i_full_n;

assign tdf12_dot_product_U0_start_full_n = 1'b1;

assign tdf12_dot_product_U0_start_write = 1'b0;

assign tdf12_get_next_ijk_U0_ap_continue = 1'b1;

assign tdf12_get_next_ijk_U0_ap_start = ((ap_sync_reg_tdf12_get_next_ijk_U0_ap_ready ^ 1'b1) & ap_start);

assign tdf12_readFilters78_U0_ap_continue = weight_vecs_0_0_0_i_full_n;

assign tdf12_readFilters78_U0_ap_start = start_for_tdf12_readFilters78_U0_empty_n;

assign tdf12_readFilters78_U0_start_full_n = 1'b1;

assign tdf12_readFilters78_U0_start_write = 1'b0;

assign tdf12_readFilters78_U0_weight_vecs_0_0_0_full_n = weight_vecs_0_0_0_i_full_n;

assign tdf12_readInputs_U0_ap_continue = ifmap_vec_0_0_i_full_n;

assign tdf12_readInputs_U0_ap_start = ((ap_sync_reg_tdf12_readInputs_U0_ap_ready ^ 1'b1) & ap_start);

assign tdf12_readInputs_U0_ifmap_vec_0_0_full_n = ifmap_vec_0_0_i_full_n;

assign tdf12_readInputs_U0_in_data_full_n = in_data_empty_n;

assign tdf12_readInputs_U0_in_data_write = 1'b0;

assign tdf12_readInputs_U0_start_full_n = 1'b1;

assign tdf12_readInputs_U0_start_write = 1'b0;

assign tdf12_writeOutputs_unaligned_U0_ap_continue = ap_continue;

assign tdf12_writeOutputs_unaligned_U0_ap_start = outputs_0_empty_n;

assign tdf12_writeOutputs_unaligned_U0_out_data_full_n = out_data_full_n;

assign tdf12_writeOutputs_unaligned_U0_out_data_write = 1'b0;

assign tdf12_writeOutputs_unaligned_U0_start_full_n = 1'b1;

assign tdf12_writeOutputs_unaligned_U0_start_write = 1'b0;

endmodule //td_fused_top_dataflow_in_loop_TOP_LOOP76
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP76_weight_vecs_0_0_0_memcore_ram (addr0, ce0, d0, we0, q0, addr1, ce1, d1, we1, q1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 8;
parameter MEM_SIZE = 256;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
output reg[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
output reg[DWIDTH-1:0] q1;
input clk;

reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];




always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
        q0 <= ram[addr0];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1) 
            ram[addr1] <= d1; 
        q1 <= ram[addr1];
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_dataflow_in_loop_TOP_LOOP76_weight_vecs_0_0_0_memcore(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    q0,
    address1,
    ce1,
    we1,
    d1,
    q1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd256;
parameter AddressWidth = 32'd8;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;
output[DataWidth - 1:0] q1;



td_fused_top_dataflow_in_loop_TOP_LOOP76_weight_vecs_0_0_0_memcore_ram td_fused_top_dataflow_in_loop_TOP_LOOP76_weight_vecs_0_0_0_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 ),
    .q1( q1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_dataflow_in_loop_TOP_LOOP76_weight_vecs_0_0_0
#(parameter
    DataWidth    = 16,
    AddressRange = 32,
    AddressWidth = 7,
    BufferCount  = 2,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire                    i_we0,
    input  wire [AddressWidth-1:0] i_address0,
    input  wire [DataWidth-1:0]    i_d0,
    output wire [DataWidth-1:0]    i_q0,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire                    t_we0,
    input  wire [AddressWidth-1:0] t_address0,
    input  wire [DataWidth-1:0]    t_d0,
    output wire [DataWidth-1:0]    t_q0
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
wire [AddressWidth+IndexWidth-1:0]   memcore_iaddr;
wire [AddressWidth+IndexWidth-1:0]   memcore_taddr;

//------------------------Instantiation------------------
assign memcore_iaddr = {i_address0, iptr};
assign memcore_taddr = {t_address0, tptr};
td_fused_top_dataflow_in_loop_TOP_LOOP76_weight_vecs_0_0_0_memcore td_fused_top_dataflow_in_loop_TOP_LOOP76_weight_vecs_0_0_0_memcore_U (
    .reset    ( reset ),
    .clk      ( clk ),
    .address0 ( memcore_iaddr ),
    .ce0      ( i_ce0 ),
    .we0      ( i_we0),
    .d0       ( i_d0 ),
    .q0       ( i_q0 ),
    .address1 ( memcore_taddr ),
    .ce1      ( t_ce0 ),
    .we1      ( t_we0),
    .d1       ( t_d0 ),
    .q1       ( t_q0 )

);

//------------------------Body---------------------------

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w10_d2_S_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd10;
parameter ADDR_WIDTH = 32'd1;
parameter DEPTH = 2'd2;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;


        end
    end

always @( sr_0, sr_1, a) begin
   case (a)
      1'd0: q = sr_0;
      1'd1: q = sr_1;
      default: q = sr_1;
   endcase
end

endmodule

module td_fused_top_fifo_w10_d2_S (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd10;
parameter ADDR_WIDTH  = 32'd1;
parameter DEPTH       = 2'd2;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 2'd1;
            if (mOutPtr == 2'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 2'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 2'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w10_d2_S_shiftReg 
U_td_fused_top_fifo_w10_d2_S_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w10_d7_S_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd10;
parameter ADDR_WIDTH = 32'd3;
parameter DEPTH = 4'd7;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;
            sr_2 <= sr_1;
            sr_3 <= sr_2;
            sr_4 <= sr_3;
            sr_5 <= sr_4;
            sr_6 <= sr_5;


        end
    end

always @( sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, a) begin
   case (a)
      3'd0: q = sr_0;
      3'd1: q = sr_1;
      3'd2: q = sr_2;
      3'd3: q = sr_3;
      3'd4: q = sr_4;
      3'd5: q = sr_5;
      3'd6: q = sr_6;
      default: q = sr_6;
   endcase
end

endmodule

module td_fused_top_fifo_w10_d7_S (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd10;
parameter ADDR_WIDTH  = 32'd3;
parameter DEPTH       = 4'd7;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 4'd1;
            if (mOutPtr == 4'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 4'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 4'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w10_d7_S_shiftReg 
U_td_fused_top_fifo_w10_d7_S_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w10_d7_S_x_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd10;
parameter ADDR_WIDTH = 32'd3;
parameter DEPTH = 4'd7;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;
            sr_2 <= sr_1;
            sr_3 <= sr_2;
            sr_4 <= sr_3;
            sr_5 <= sr_4;
            sr_6 <= sr_5;


        end
    end

always @( sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, a) begin
   case (a)
      3'd0: q = sr_0;
      3'd1: q = sr_1;
      3'd2: q = sr_2;
      3'd3: q = sr_3;
      3'd4: q = sr_4;
      3'd5: q = sr_5;
      3'd6: q = sr_6;
      default: q = sr_6;
   endcase
end

endmodule

module td_fused_top_fifo_w10_d7_S_x (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd10;
parameter ADDR_WIDTH  = 32'd3;
parameter DEPTH       = 4'd7;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 4'd1;
            if (mOutPtr == 4'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 4'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 4'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w10_d7_S_x_shiftReg 
U_td_fused_top_fifo_w10_d7_S_x_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w10_d8_S_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd10;
parameter ADDR_WIDTH = 32'd3;
parameter DEPTH = 4'd8;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, sr_7;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;
            sr_2 <= sr_1;
            sr_3 <= sr_2;
            sr_4 <= sr_3;
            sr_5 <= sr_4;
            sr_6 <= sr_5;
            sr_7 <= sr_6;


        end
    end

always @( sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, sr_7, a) begin
   case (a)
      3'd0: q = sr_0;
      3'd1: q = sr_1;
      3'd2: q = sr_2;
      3'd3: q = sr_3;
      3'd4: q = sr_4;
      3'd5: q = sr_5;
      3'd6: q = sr_6;
      3'd7: q = sr_7;
      default: q = sr_7;
   endcase
end

endmodule

module td_fused_top_fifo_w10_d8_S (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd10;
parameter ADDR_WIDTH  = 32'd3;
parameter DEPTH       = 4'd8;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 4'd1;
            if (mOutPtr == 4'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 4'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 4'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w10_d8_S_shiftReg 
U_td_fused_top_fifo_w10_d8_S_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w10_d8_S_x_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd10;
parameter ADDR_WIDTH = 32'd3;
parameter DEPTH = 4'd8;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, sr_7;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;
            sr_2 <= sr_1;
            sr_3 <= sr_2;
            sr_4 <= sr_3;
            sr_5 <= sr_4;
            sr_6 <= sr_5;
            sr_7 <= sr_6;


        end
    end

always @( sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, sr_7, a) begin
   case (a)
      3'd0: q = sr_0;
      3'd1: q = sr_1;
      3'd2: q = sr_2;
      3'd3: q = sr_3;
      3'd4: q = sr_4;
      3'd5: q = sr_5;
      3'd6: q = sr_6;
      3'd7: q = sr_7;
      default: q = sr_7;
   endcase
end

endmodule

module td_fused_top_fifo_w10_d8_S_x (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd10;
parameter ADDR_WIDTH  = 32'd3;
parameter DEPTH       = 4'd8;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 4'd1;
            if (mOutPtr == 4'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 4'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 4'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w10_d8_S_x_shiftReg 
U_td_fused_top_fifo_w10_d8_S_x_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w11_d2_S_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd11;
parameter ADDR_WIDTH = 32'd1;
parameter DEPTH = 2'd2;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;


        end
    end

always @( sr_0, sr_1, a) begin
   case (a)
      1'd0: q = sr_0;
      1'd1: q = sr_1;
      default: q = sr_1;
   endcase
end

endmodule

module td_fused_top_fifo_w11_d2_S (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd11;
parameter ADDR_WIDTH  = 32'd1;
parameter DEPTH       = 2'd2;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 2'd1;
            if (mOutPtr == 2'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 2'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 2'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w11_d2_S_shiftReg 
U_td_fused_top_fifo_w11_d2_S_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w11_d7_S_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd11;
parameter ADDR_WIDTH = 32'd3;
parameter DEPTH = 4'd7;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;
            sr_2 <= sr_1;
            sr_3 <= sr_2;
            sr_4 <= sr_3;
            sr_5 <= sr_4;
            sr_6 <= sr_5;


        end
    end

always @( sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, a) begin
   case (a)
      3'd0: q = sr_0;
      3'd1: q = sr_1;
      3'd2: q = sr_2;
      3'd3: q = sr_3;
      3'd4: q = sr_4;
      3'd5: q = sr_5;
      3'd6: q = sr_6;
      default: q = sr_6;
   endcase
end

endmodule

module td_fused_top_fifo_w11_d7_S (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd11;
parameter ADDR_WIDTH  = 32'd3;
parameter DEPTH       = 4'd7;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 4'd1;
            if (mOutPtr == 4'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 4'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 4'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w11_d7_S_shiftReg 
U_td_fused_top_fifo_w11_d7_S_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w12_d7_S_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd12;
parameter ADDR_WIDTH = 32'd3;
parameter DEPTH = 4'd7;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;
            sr_2 <= sr_1;
            sr_3 <= sr_2;
            sr_4 <= sr_3;
            sr_5 <= sr_4;
            sr_6 <= sr_5;


        end
    end

always @( sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, a) begin
   case (a)
      3'd0: q = sr_0;
      3'd1: q = sr_1;
      3'd2: q = sr_2;
      3'd3: q = sr_3;
      3'd4: q = sr_4;
      3'd5: q = sr_5;
      3'd6: q = sr_6;
      default: q = sr_6;
   endcase
end

endmodule

module td_fused_top_fifo_w12_d7_S (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd12;
parameter ADDR_WIDTH  = 32'd3;
parameter DEPTH       = 4'd7;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 4'd1;
            if (mOutPtr == 4'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 4'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 4'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w12_d7_S_shiftReg 
U_td_fused_top_fifo_w12_d7_S_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w12_d8_S_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd12;
parameter ADDR_WIDTH = 32'd3;
parameter DEPTH = 4'd8;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, sr_7;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;
            sr_2 <= sr_1;
            sr_3 <= sr_2;
            sr_4 <= sr_3;
            sr_5 <= sr_4;
            sr_6 <= sr_5;
            sr_7 <= sr_6;


        end
    end

always @( sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, sr_7, a) begin
   case (a)
      3'd0: q = sr_0;
      3'd1: q = sr_1;
      3'd2: q = sr_2;
      3'd3: q = sr_3;
      3'd4: q = sr_4;
      3'd5: q = sr_5;
      3'd6: q = sr_6;
      3'd7: q = sr_7;
      default: q = sr_7;
   endcase
end

endmodule

module td_fused_top_fifo_w12_d8_S (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd12;
parameter ADDR_WIDTH  = 32'd3;
parameter DEPTH       = 4'd8;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 4'd1;
            if (mOutPtr == 4'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 4'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 4'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w12_d8_S_shiftReg 
U_td_fused_top_fifo_w12_d8_S_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w12_d8_S_x_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd12;
parameter ADDR_WIDTH = 32'd3;
parameter DEPTH = 4'd8;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, sr_7;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;
            sr_2 <= sr_1;
            sr_3 <= sr_2;
            sr_4 <= sr_3;
            sr_5 <= sr_4;
            sr_6 <= sr_5;
            sr_7 <= sr_6;


        end
    end

always @( sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, sr_7, a) begin
   case (a)
      3'd0: q = sr_0;
      3'd1: q = sr_1;
      3'd2: q = sr_2;
      3'd3: q = sr_3;
      3'd4: q = sr_4;
      3'd5: q = sr_5;
      3'd6: q = sr_6;
      3'd7: q = sr_7;
      default: q = sr_7;
   endcase
end

endmodule

module td_fused_top_fifo_w12_d8_S_x (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd12;
parameter ADDR_WIDTH  = 32'd3;
parameter DEPTH       = 4'd8;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 4'd1;
            if (mOutPtr == 4'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 4'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 4'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w12_d8_S_x_shiftReg 
U_td_fused_top_fifo_w12_d8_S_x_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w13_d2_S_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd13;
parameter ADDR_WIDTH = 32'd1;
parameter DEPTH = 2'd2;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;


        end
    end

always @( sr_0, sr_1, a) begin
   case (a)
      1'd0: q = sr_0;
      1'd1: q = sr_1;
      default: q = sr_1;
   endcase
end

endmodule

module td_fused_top_fifo_w13_d2_S (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd13;
parameter ADDR_WIDTH  = 32'd1;
parameter DEPTH       = 2'd2;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 2'd1;
            if (mOutPtr == 2'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 2'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 2'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w13_d2_S_shiftReg 
U_td_fused_top_fifo_w13_d2_S_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w13_d7_S_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd13;
parameter ADDR_WIDTH = 32'd3;
parameter DEPTH = 4'd7;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;
            sr_2 <= sr_1;
            sr_3 <= sr_2;
            sr_4 <= sr_3;
            sr_5 <= sr_4;
            sr_6 <= sr_5;


        end
    end

always @( sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, a) begin
   case (a)
      3'd0: q = sr_0;
      3'd1: q = sr_1;
      3'd2: q = sr_2;
      3'd3: q = sr_3;
      3'd4: q = sr_4;
      3'd5: q = sr_5;
      3'd6: q = sr_6;
      default: q = sr_6;
   endcase
end

endmodule

module td_fused_top_fifo_w13_d7_S (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd13;
parameter ADDR_WIDTH  = 32'd3;
parameter DEPTH       = 4'd7;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 4'd1;
            if (mOutPtr == 4'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 4'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 4'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w13_d7_S_shiftReg 
U_td_fused_top_fifo_w13_d7_S_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w14_d9_S_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd14;
parameter ADDR_WIDTH = 32'd4;
parameter DEPTH = 5'd9;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, sr_7, sr_8;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;
            sr_2 <= sr_1;
            sr_3 <= sr_2;
            sr_4 <= sr_3;
            sr_5 <= sr_4;
            sr_6 <= sr_5;
            sr_7 <= sr_6;
            sr_8 <= sr_7;


        end
    end

always @( sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, sr_7, sr_8, a) begin
   case (a)
      4'd0: q = sr_0;
      4'd1: q = sr_1;
      4'd2: q = sr_2;
      4'd3: q = sr_3;
      4'd4: q = sr_4;
      4'd5: q = sr_5;
      4'd6: q = sr_6;
      4'd7: q = sr_7;
      4'd8: q = sr_8;
      default: q = sr_8;
   endcase
end

endmodule

module td_fused_top_fifo_w14_d9_S (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd14;
parameter ADDR_WIDTH  = 32'd4;
parameter DEPTH       = 5'd9;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 5'd1;
            if (mOutPtr == 5'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 5'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 5'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w14_d9_S_shiftReg 
U_td_fused_top_fifo_w14_d9_S_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w15_d2_S_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd15;
parameter ADDR_WIDTH = 32'd1;
parameter DEPTH = 2'd2;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;


        end
    end

always @( sr_0, sr_1, a) begin
   case (a)
      1'd0: q = sr_0;
      1'd1: q = sr_1;
      default: q = sr_1;
   endcase
end

endmodule

module td_fused_top_fifo_w15_d2_S (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd15;
parameter ADDR_WIDTH  = 32'd1;
parameter DEPTH       = 2'd2;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 2'd1;
            if (mOutPtr == 2'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 2'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 2'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w15_d2_S_shiftReg 
U_td_fused_top_fifo_w15_d2_S_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w15_d7_S_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd15;
parameter ADDR_WIDTH = 32'd3;
parameter DEPTH = 4'd7;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;
            sr_2 <= sr_1;
            sr_3 <= sr_2;
            sr_4 <= sr_3;
            sr_5 <= sr_4;
            sr_6 <= sr_5;


        end
    end

always @( sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, a) begin
   case (a)
      3'd0: q = sr_0;
      3'd1: q = sr_1;
      3'd2: q = sr_2;
      3'd3: q = sr_3;
      3'd4: q = sr_4;
      3'd5: q = sr_5;
      3'd6: q = sr_6;
      default: q = sr_6;
   endcase
end

endmodule

module td_fused_top_fifo_w15_d7_S (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd15;
parameter ADDR_WIDTH  = 32'd3;
parameter DEPTH       = 4'd7;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 4'd1;
            if (mOutPtr == 4'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 4'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 4'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w15_d7_S_shiftReg 
U_td_fused_top_fifo_w15_d7_S_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w16_d2_S_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd16;
parameter ADDR_WIDTH = 32'd1;
parameter DEPTH = 2'd2;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;


        end
    end

always @( sr_0, sr_1, a) begin
   case (a)
      1'd0: q = sr_0;
      1'd1: q = sr_1;
      default: q = sr_1;
   endcase
end

endmodule

module td_fused_top_fifo_w16_d2_S (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd16;
parameter ADDR_WIDTH  = 32'd1;
parameter DEPTH       = 2'd2;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 2'd1;
            if (mOutPtr == 2'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 2'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 2'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w16_d2_S_shiftReg 
U_td_fused_top_fifo_w16_d2_S_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w16_d2_S_x0_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd16;
parameter ADDR_WIDTH = 32'd1;
parameter DEPTH = 2'd2;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;


        end
    end

always @( sr_0, sr_1, a) begin
   case (a)
      1'd0: q = sr_0;
      1'd1: q = sr_1;
      default: q = sr_1;
   endcase
end

endmodule

module td_fused_top_fifo_w16_d2_S_x0 (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd16;
parameter ADDR_WIDTH  = 32'd1;
parameter DEPTH       = 2'd2;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 2'd1;
            if (mOutPtr == 2'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 2'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 2'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w16_d2_S_x0_shiftReg 
U_td_fused_top_fifo_w16_d2_S_x0_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w16_d2_S_x1_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd16;
parameter ADDR_WIDTH = 32'd1;
parameter DEPTH = 2'd2;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;


        end
    end

always @( sr_0, sr_1, a) begin
   case (a)
      1'd0: q = sr_0;
      1'd1: q = sr_1;
      default: q = sr_1;
   endcase
end

endmodule

module td_fused_top_fifo_w16_d2_S_x1 (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd16;
parameter ADDR_WIDTH  = 32'd1;
parameter DEPTH       = 2'd2;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 2'd1;
            if (mOutPtr == 2'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 2'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 2'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w16_d2_S_x1_shiftReg 
U_td_fused_top_fifo_w16_d2_S_x1_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w16_d2_S_x2_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd16;
parameter ADDR_WIDTH = 32'd1;
parameter DEPTH = 2'd2;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;


        end
    end

always @( sr_0, sr_1, a) begin
   case (a)
      1'd0: q = sr_0;
      1'd1: q = sr_1;
      default: q = sr_1;
   endcase
end

endmodule

module td_fused_top_fifo_w16_d2_S_x2 (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd16;
parameter ADDR_WIDTH  = 32'd1;
parameter DEPTH       = 2'd2;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 2'd1;
            if (mOutPtr == 2'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 2'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 2'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w16_d2_S_x2_shiftReg 
U_td_fused_top_fifo_w16_d2_S_x2_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w16_d2_S_x3_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd16;
parameter ADDR_WIDTH = 32'd1;
parameter DEPTH = 2'd2;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;


        end
    end

always @( sr_0, sr_1, a) begin
   case (a)
      1'd0: q = sr_0;
      1'd1: q = sr_1;
      default: q = sr_1;
   endcase
end

endmodule

module td_fused_top_fifo_w16_d2_S_x3 (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd16;
parameter ADDR_WIDTH  = 32'd1;
parameter DEPTH       = 2'd2;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 2'd1;
            if (mOutPtr == 2'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 2'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 2'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w16_d2_S_x3_shiftReg 
U_td_fused_top_fifo_w16_d2_S_x3_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w16_d2_S_x4_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd16;
parameter ADDR_WIDTH = 32'd1;
parameter DEPTH = 2'd2;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;


        end
    end

always @( sr_0, sr_1, a) begin
   case (a)
      1'd0: q = sr_0;
      1'd1: q = sr_1;
      default: q = sr_1;
   endcase
end

endmodule

module td_fused_top_fifo_w16_d2_S_x4 (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd16;
parameter ADDR_WIDTH  = 32'd1;
parameter DEPTH       = 2'd2;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 2'd1;
            if (mOutPtr == 2'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 2'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 2'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w16_d2_S_x4_shiftReg 
U_td_fused_top_fifo_w16_d2_S_x4_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w16_d2_S_x5_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd16;
parameter ADDR_WIDTH = 32'd1;
parameter DEPTH = 2'd2;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;


        end
    end

always @( sr_0, sr_1, a) begin
   case (a)
      1'd0: q = sr_0;
      1'd1: q = sr_1;
      default: q = sr_1;
   endcase
end

endmodule

module td_fused_top_fifo_w16_d2_S_x5 (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd16;
parameter ADDR_WIDTH  = 32'd1;
parameter DEPTH       = 2'd2;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 2'd1;
            if (mOutPtr == 2'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 2'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 2'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w16_d2_S_x5_shiftReg 
U_td_fused_top_fifo_w16_d2_S_x5_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w16_d2_S_x6_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd16;
parameter ADDR_WIDTH = 32'd1;
parameter DEPTH = 2'd2;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;


        end
    end

always @( sr_0, sr_1, a) begin
   case (a)
      1'd0: q = sr_0;
      1'd1: q = sr_1;
      default: q = sr_1;
   endcase
end

endmodule

module td_fused_top_fifo_w16_d2_S_x6 (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd16;
parameter ADDR_WIDTH  = 32'd1;
parameter DEPTH       = 2'd2;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 2'd1;
            if (mOutPtr == 2'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 2'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 2'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w16_d2_S_x6_shiftReg 
U_td_fused_top_fifo_w16_d2_S_x6_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w16_d2_S_x7_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd16;
parameter ADDR_WIDTH = 32'd1;
parameter DEPTH = 2'd2;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;


        end
    end

always @( sr_0, sr_1, a) begin
   case (a)
      1'd0: q = sr_0;
      1'd1: q = sr_1;
      default: q = sr_1;
   endcase
end

endmodule

module td_fused_top_fifo_w16_d2_S_x7 (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd16;
parameter ADDR_WIDTH  = 32'd1;
parameter DEPTH       = 2'd2;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 2'd1;
            if (mOutPtr == 2'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 2'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 2'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w16_d2_S_x7_shiftReg 
U_td_fused_top_fifo_w16_d2_S_x7_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w16_d2_S_x8_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd16;
parameter ADDR_WIDTH = 32'd1;
parameter DEPTH = 2'd2;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;


        end
    end

always @( sr_0, sr_1, a) begin
   case (a)
      1'd0: q = sr_0;
      1'd1: q = sr_1;
      default: q = sr_1;
   endcase
end

endmodule

module td_fused_top_fifo_w16_d2_S_x8 (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd16;
parameter ADDR_WIDTH  = 32'd1;
parameter DEPTH       = 2'd2;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 2'd1;
            if (mOutPtr == 2'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 2'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 2'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w16_d2_S_x8_shiftReg 
U_td_fused_top_fifo_w16_d2_S_x8_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w16_d2_S_x9_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd16;
parameter ADDR_WIDTH = 32'd1;
parameter DEPTH = 2'd2;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;


        end
    end

always @( sr_0, sr_1, a) begin
   case (a)
      1'd0: q = sr_0;
      1'd1: q = sr_1;
      default: q = sr_1;
   endcase
end

endmodule

module td_fused_top_fifo_w16_d2_S_x9 (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd16;
parameter ADDR_WIDTH  = 32'd1;
parameter DEPTH       = 2'd2;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 2'd1;
            if (mOutPtr == 2'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 2'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 2'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w16_d2_S_x9_shiftReg 
U_td_fused_top_fifo_w16_d2_S_x9_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w16_d2_S_x_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd16;
parameter ADDR_WIDTH = 32'd1;
parameter DEPTH = 2'd2;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;


        end
    end

always @( sr_0, sr_1, a) begin
   case (a)
      1'd0: q = sr_0;
      1'd1: q = sr_1;
      default: q = sr_1;
   endcase
end

endmodule

module td_fused_top_fifo_w16_d2_S_x (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd16;
parameter ADDR_WIDTH  = 32'd1;
parameter DEPTH       = 2'd2;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 2'd1;
            if (mOutPtr == 2'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 2'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 2'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w16_d2_S_x_shiftReg 
U_td_fused_top_fifo_w16_d2_S_x_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w1_d8_S_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd1;
parameter ADDR_WIDTH = 32'd3;
parameter DEPTH = 4'd8;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, sr_7;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;
            sr_2 <= sr_1;
            sr_3 <= sr_2;
            sr_4 <= sr_3;
            sr_5 <= sr_4;
            sr_6 <= sr_5;
            sr_7 <= sr_6;


        end
    end

always @( sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, sr_7, a) begin
   case (a)
      3'd0: q = sr_0;
      3'd1: q = sr_1;
      3'd2: q = sr_2;
      3'd3: q = sr_3;
      3'd4: q = sr_4;
      3'd5: q = sr_5;
      3'd6: q = sr_6;
      3'd7: q = sr_7;
      default: q = sr_7;
   endcase
end

endmodule

module td_fused_top_fifo_w1_d8_S (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd1;
parameter ADDR_WIDTH  = 32'd3;
parameter DEPTH       = 4'd8;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 4'd1;
            if (mOutPtr == 4'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 4'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 4'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w1_d8_S_shiftReg 
U_td_fused_top_fifo_w1_d8_S_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w1_d8_S_x0_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd1;
parameter ADDR_WIDTH = 32'd3;
parameter DEPTH = 4'd8;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, sr_7;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;
            sr_2 <= sr_1;
            sr_3 <= sr_2;
            sr_4 <= sr_3;
            sr_5 <= sr_4;
            sr_6 <= sr_5;
            sr_7 <= sr_6;


        end
    end

always @( sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, sr_7, a) begin
   case (a)
      3'd0: q = sr_0;
      3'd1: q = sr_1;
      3'd2: q = sr_2;
      3'd3: q = sr_3;
      3'd4: q = sr_4;
      3'd5: q = sr_5;
      3'd6: q = sr_6;
      3'd7: q = sr_7;
      default: q = sr_7;
   endcase
end

endmodule

module td_fused_top_fifo_w1_d8_S_x0 (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd1;
parameter ADDR_WIDTH  = 32'd3;
parameter DEPTH       = 4'd8;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 4'd1;
            if (mOutPtr == 4'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 4'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 4'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w1_d8_S_x0_shiftReg 
U_td_fused_top_fifo_w1_d8_S_x0_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w1_d8_S_x_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd1;
parameter ADDR_WIDTH = 32'd3;
parameter DEPTH = 4'd8;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, sr_7;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;
            sr_2 <= sr_1;
            sr_3 <= sr_2;
            sr_4 <= sr_3;
            sr_5 <= sr_4;
            sr_6 <= sr_5;
            sr_7 <= sr_6;


        end
    end

always @( sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, sr_7, a) begin
   case (a)
      3'd0: q = sr_0;
      3'd1: q = sr_1;
      3'd2: q = sr_2;
      3'd3: q = sr_3;
      3'd4: q = sr_4;
      3'd5: q = sr_5;
      3'd6: q = sr_6;
      3'd7: q = sr_7;
      default: q = sr_7;
   endcase
end

endmodule

module td_fused_top_fifo_w1_d8_S_x (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd1;
parameter ADDR_WIDTH  = 32'd3;
parameter DEPTH       = 4'd8;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 4'd1;
            if (mOutPtr == 4'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 4'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 4'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w1_d8_S_x_shiftReg 
U_td_fused_top_fifo_w1_d8_S_x_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w1_d9_S_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd1;
parameter ADDR_WIDTH = 32'd4;
parameter DEPTH = 5'd9;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, sr_7, sr_8;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;
            sr_2 <= sr_1;
            sr_3 <= sr_2;
            sr_4 <= sr_3;
            sr_5 <= sr_4;
            sr_6 <= sr_5;
            sr_7 <= sr_6;
            sr_8 <= sr_7;


        end
    end

always @( sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, sr_7, sr_8, a) begin
   case (a)
      4'd0: q = sr_0;
      4'd1: q = sr_1;
      4'd2: q = sr_2;
      4'd3: q = sr_3;
      4'd4: q = sr_4;
      4'd5: q = sr_5;
      4'd6: q = sr_6;
      4'd7: q = sr_7;
      4'd8: q = sr_8;
      default: q = sr_8;
   endcase
end

endmodule

module td_fused_top_fifo_w1_d9_S (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd1;
parameter ADDR_WIDTH  = 32'd4;
parameter DEPTH       = 5'd9;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 5'd1;
            if (mOutPtr == 5'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 5'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 5'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w1_d9_S_shiftReg 
U_td_fused_top_fifo_w1_d9_S_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w1_d9_S_x0_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd1;
parameter ADDR_WIDTH = 32'd4;
parameter DEPTH = 5'd9;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, sr_7, sr_8;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;
            sr_2 <= sr_1;
            sr_3 <= sr_2;
            sr_4 <= sr_3;
            sr_5 <= sr_4;
            sr_6 <= sr_5;
            sr_7 <= sr_6;
            sr_8 <= sr_7;


        end
    end

always @( sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, sr_7, sr_8, a) begin
   case (a)
      4'd0: q = sr_0;
      4'd1: q = sr_1;
      4'd2: q = sr_2;
      4'd3: q = sr_3;
      4'd4: q = sr_4;
      4'd5: q = sr_5;
      4'd6: q = sr_6;
      4'd7: q = sr_7;
      4'd8: q = sr_8;
      default: q = sr_8;
   endcase
end

endmodule

module td_fused_top_fifo_w1_d9_S_x0 (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd1;
parameter ADDR_WIDTH  = 32'd4;
parameter DEPTH       = 5'd9;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 5'd1;
            if (mOutPtr == 5'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 5'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 5'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w1_d9_S_x0_shiftReg 
U_td_fused_top_fifo_w1_d9_S_x0_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w1_d9_S_x1_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd1;
parameter ADDR_WIDTH = 32'd4;
parameter DEPTH = 5'd9;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, sr_7, sr_8;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;
            sr_2 <= sr_1;
            sr_3 <= sr_2;
            sr_4 <= sr_3;
            sr_5 <= sr_4;
            sr_6 <= sr_5;
            sr_7 <= sr_6;
            sr_8 <= sr_7;


        end
    end

always @( sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, sr_7, sr_8, a) begin
   case (a)
      4'd0: q = sr_0;
      4'd1: q = sr_1;
      4'd2: q = sr_2;
      4'd3: q = sr_3;
      4'd4: q = sr_4;
      4'd5: q = sr_5;
      4'd6: q = sr_6;
      4'd7: q = sr_7;
      4'd8: q = sr_8;
      default: q = sr_8;
   endcase
end

endmodule

module td_fused_top_fifo_w1_d9_S_x1 (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd1;
parameter ADDR_WIDTH  = 32'd4;
parameter DEPTH       = 5'd9;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 5'd1;
            if (mOutPtr == 5'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 5'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 5'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w1_d9_S_x1_shiftReg 
U_td_fused_top_fifo_w1_d9_S_x1_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w1_d9_S_x2_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd1;
parameter ADDR_WIDTH = 32'd4;
parameter DEPTH = 5'd9;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, sr_7, sr_8;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;
            sr_2 <= sr_1;
            sr_3 <= sr_2;
            sr_4 <= sr_3;
            sr_5 <= sr_4;
            sr_6 <= sr_5;
            sr_7 <= sr_6;
            sr_8 <= sr_7;


        end
    end

always @( sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, sr_7, sr_8, a) begin
   case (a)
      4'd0: q = sr_0;
      4'd1: q = sr_1;
      4'd2: q = sr_2;
      4'd3: q = sr_3;
      4'd4: q = sr_4;
      4'd5: q = sr_5;
      4'd6: q = sr_6;
      4'd7: q = sr_7;
      4'd8: q = sr_8;
      default: q = sr_8;
   endcase
end

endmodule

module td_fused_top_fifo_w1_d9_S_x2 (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd1;
parameter ADDR_WIDTH  = 32'd4;
parameter DEPTH       = 5'd9;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 5'd1;
            if (mOutPtr == 5'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 5'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 5'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w1_d9_S_x2_shiftReg 
U_td_fused_top_fifo_w1_d9_S_x2_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w1_d9_S_x_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd1;
parameter ADDR_WIDTH = 32'd4;
parameter DEPTH = 5'd9;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, sr_7, sr_8;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;
            sr_2 <= sr_1;
            sr_3 <= sr_2;
            sr_4 <= sr_3;
            sr_5 <= sr_4;
            sr_6 <= sr_5;
            sr_7 <= sr_6;
            sr_8 <= sr_7;


        end
    end

always @( sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, sr_7, sr_8, a) begin
   case (a)
      4'd0: q = sr_0;
      4'd1: q = sr_1;
      4'd2: q = sr_2;
      4'd3: q = sr_3;
      4'd4: q = sr_4;
      4'd5: q = sr_5;
      4'd6: q = sr_6;
      4'd7: q = sr_7;
      4'd8: q = sr_8;
      default: q = sr_8;
   endcase
end

endmodule

module td_fused_top_fifo_w1_d9_S_x (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd1;
parameter ADDR_WIDTH  = 32'd4;
parameter DEPTH       = 5'd9;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 5'd1;
            if (mOutPtr == 5'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 5'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 5'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w1_d9_S_x_shiftReg 
U_td_fused_top_fifo_w1_d9_S_x_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w4_d2_S_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd4;
parameter ADDR_WIDTH = 32'd1;
parameter DEPTH = 2'd2;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;


        end
    end

always @( sr_0, sr_1, a) begin
   case (a)
      1'd0: q = sr_0;
      1'd1: q = sr_1;
      default: q = sr_1;
   endcase
end

endmodule

module td_fused_top_fifo_w4_d2_S (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd4;
parameter ADDR_WIDTH  = 32'd1;
parameter DEPTH       = 2'd2;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 2'd1;
            if (mOutPtr == 2'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 2'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 2'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w4_d2_S_shiftReg 
U_td_fused_top_fifo_w4_d2_S_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w4_d2_S_x_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd4;
parameter ADDR_WIDTH = 32'd1;
parameter DEPTH = 2'd2;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;


        end
    end

always @( sr_0, sr_1, a) begin
   case (a)
      1'd0: q = sr_0;
      1'd1: q = sr_1;
      default: q = sr_1;
   endcase
end

endmodule

module td_fused_top_fifo_w4_d2_S_x (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd4;
parameter ADDR_WIDTH  = 32'd1;
parameter DEPTH       = 2'd2;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 2'd1;
            if (mOutPtr == 2'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 2'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 2'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w4_d2_S_x_shiftReg 
U_td_fused_top_fifo_w4_d2_S_x_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w4_d7_S_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd4;
parameter ADDR_WIDTH = 32'd3;
parameter DEPTH = 4'd7;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;
            sr_2 <= sr_1;
            sr_3 <= sr_2;
            sr_4 <= sr_3;
            sr_5 <= sr_4;
            sr_6 <= sr_5;


        end
    end

always @( sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, a) begin
   case (a)
      3'd0: q = sr_0;
      3'd1: q = sr_1;
      3'd2: q = sr_2;
      3'd3: q = sr_3;
      3'd4: q = sr_4;
      3'd5: q = sr_5;
      3'd6: q = sr_6;
      default: q = sr_6;
   endcase
end

endmodule

module td_fused_top_fifo_w4_d7_S (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd4;
parameter ADDR_WIDTH  = 32'd3;
parameter DEPTH       = 4'd7;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 4'd1;
            if (mOutPtr == 4'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 4'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 4'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w4_d7_S_shiftReg 
U_td_fused_top_fifo_w4_d7_S_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w4_d7_S_x0_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd4;
parameter ADDR_WIDTH = 32'd3;
parameter DEPTH = 4'd7;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;
            sr_2 <= sr_1;
            sr_3 <= sr_2;
            sr_4 <= sr_3;
            sr_5 <= sr_4;
            sr_6 <= sr_5;


        end
    end

always @( sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, a) begin
   case (a)
      3'd0: q = sr_0;
      3'd1: q = sr_1;
      3'd2: q = sr_2;
      3'd3: q = sr_3;
      3'd4: q = sr_4;
      3'd5: q = sr_5;
      3'd6: q = sr_6;
      default: q = sr_6;
   endcase
end

endmodule

module td_fused_top_fifo_w4_d7_S_x0 (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd4;
parameter ADDR_WIDTH  = 32'd3;
parameter DEPTH       = 4'd7;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 4'd1;
            if (mOutPtr == 4'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 4'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 4'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w4_d7_S_x0_shiftReg 
U_td_fused_top_fifo_w4_d7_S_x0_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w4_d7_S_x_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd4;
parameter ADDR_WIDTH = 32'd3;
parameter DEPTH = 4'd7;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;
            sr_2 <= sr_1;
            sr_3 <= sr_2;
            sr_4 <= sr_3;
            sr_5 <= sr_4;
            sr_6 <= sr_5;


        end
    end

always @( sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, a) begin
   case (a)
      3'd0: q = sr_0;
      3'd1: q = sr_1;
      3'd2: q = sr_2;
      3'd3: q = sr_3;
      3'd4: q = sr_4;
      3'd5: q = sr_5;
      3'd6: q = sr_6;
      default: q = sr_6;
   endcase
end

endmodule

module td_fused_top_fifo_w4_d7_S_x (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd4;
parameter ADDR_WIDTH  = 32'd3;
parameter DEPTH       = 4'd7;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 4'd1;
            if (mOutPtr == 4'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 4'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 4'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w4_d7_S_x_shiftReg 
U_td_fused_top_fifo_w4_d7_S_x_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w4_d8_S_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd4;
parameter ADDR_WIDTH = 32'd3;
parameter DEPTH = 4'd8;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, sr_7;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;
            sr_2 <= sr_1;
            sr_3 <= sr_2;
            sr_4 <= sr_3;
            sr_5 <= sr_4;
            sr_6 <= sr_5;
            sr_7 <= sr_6;


        end
    end

always @( sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, sr_7, a) begin
   case (a)
      3'd0: q = sr_0;
      3'd1: q = sr_1;
      3'd2: q = sr_2;
      3'd3: q = sr_3;
      3'd4: q = sr_4;
      3'd5: q = sr_5;
      3'd6: q = sr_6;
      3'd7: q = sr_7;
      default: q = sr_7;
   endcase
end

endmodule

module td_fused_top_fifo_w4_d8_S (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd4;
parameter ADDR_WIDTH  = 32'd3;
parameter DEPTH       = 4'd8;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 4'd1;
            if (mOutPtr == 4'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 4'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 4'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w4_d8_S_shiftReg 
U_td_fused_top_fifo_w4_d8_S_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w4_d8_S_x0_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd4;
parameter ADDR_WIDTH = 32'd3;
parameter DEPTH = 4'd8;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, sr_7;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;
            sr_2 <= sr_1;
            sr_3 <= sr_2;
            sr_4 <= sr_3;
            sr_5 <= sr_4;
            sr_6 <= sr_5;
            sr_7 <= sr_6;


        end
    end

always @( sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, sr_7, a) begin
   case (a)
      3'd0: q = sr_0;
      3'd1: q = sr_1;
      3'd2: q = sr_2;
      3'd3: q = sr_3;
      3'd4: q = sr_4;
      3'd5: q = sr_5;
      3'd6: q = sr_6;
      3'd7: q = sr_7;
      default: q = sr_7;
   endcase
end

endmodule

module td_fused_top_fifo_w4_d8_S_x0 (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd4;
parameter ADDR_WIDTH  = 32'd3;
parameter DEPTH       = 4'd8;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 4'd1;
            if (mOutPtr == 4'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 4'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 4'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w4_d8_S_x0_shiftReg 
U_td_fused_top_fifo_w4_d8_S_x0_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w4_d8_S_x1_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd4;
parameter ADDR_WIDTH = 32'd3;
parameter DEPTH = 4'd8;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, sr_7;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;
            sr_2 <= sr_1;
            sr_3 <= sr_2;
            sr_4 <= sr_3;
            sr_5 <= sr_4;
            sr_6 <= sr_5;
            sr_7 <= sr_6;


        end
    end

always @( sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, sr_7, a) begin
   case (a)
      3'd0: q = sr_0;
      3'd1: q = sr_1;
      3'd2: q = sr_2;
      3'd3: q = sr_3;
      3'd4: q = sr_4;
      3'd5: q = sr_5;
      3'd6: q = sr_6;
      3'd7: q = sr_7;
      default: q = sr_7;
   endcase
end

endmodule

module td_fused_top_fifo_w4_d8_S_x1 (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd4;
parameter ADDR_WIDTH  = 32'd3;
parameter DEPTH       = 4'd8;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 4'd1;
            if (mOutPtr == 4'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 4'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 4'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w4_d8_S_x1_shiftReg 
U_td_fused_top_fifo_w4_d8_S_x1_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w4_d8_S_x_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd4;
parameter ADDR_WIDTH = 32'd3;
parameter DEPTH = 4'd8;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, sr_7;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;
            sr_2 <= sr_1;
            sr_3 <= sr_2;
            sr_4 <= sr_3;
            sr_5 <= sr_4;
            sr_6 <= sr_5;
            sr_7 <= sr_6;


        end
    end

always @( sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, sr_7, a) begin
   case (a)
      3'd0: q = sr_0;
      3'd1: q = sr_1;
      3'd2: q = sr_2;
      3'd3: q = sr_3;
      3'd4: q = sr_4;
      3'd5: q = sr_5;
      3'd6: q = sr_6;
      3'd7: q = sr_7;
      default: q = sr_7;
   endcase
end

endmodule

module td_fused_top_fifo_w4_d8_S_x (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd4;
parameter ADDR_WIDTH  = 32'd3;
parameter DEPTH       = 4'd8;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 4'd1;
            if (mOutPtr == 4'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 4'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 4'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w4_d8_S_x_shiftReg 
U_td_fused_top_fifo_w4_d8_S_x_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w5_d2_S_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd5;
parameter ADDR_WIDTH = 32'd1;
parameter DEPTH = 2'd2;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;


        end
    end

always @( sr_0, sr_1, a) begin
   case (a)
      1'd0: q = sr_0;
      1'd1: q = sr_1;
      default: q = sr_1;
   endcase
end

endmodule

module td_fused_top_fifo_w5_d2_S (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd5;
parameter ADDR_WIDTH  = 32'd1;
parameter DEPTH       = 2'd2;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 2'd1;
            if (mOutPtr == 2'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 2'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 2'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w5_d2_S_shiftReg 
U_td_fused_top_fifo_w5_d2_S_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w5_d2_S_x_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd5;
parameter ADDR_WIDTH = 32'd1;
parameter DEPTH = 2'd2;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;


        end
    end

always @( sr_0, sr_1, a) begin
   case (a)
      1'd0: q = sr_0;
      1'd1: q = sr_1;
      default: q = sr_1;
   endcase
end

endmodule

module td_fused_top_fifo_w5_d2_S_x (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd5;
parameter ADDR_WIDTH  = 32'd1;
parameter DEPTH       = 2'd2;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 2'd1;
            if (mOutPtr == 2'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 2'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 2'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w5_d2_S_x_shiftReg 
U_td_fused_top_fifo_w5_d2_S_x_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w5_d7_S_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd5;
parameter ADDR_WIDTH = 32'd3;
parameter DEPTH = 4'd7;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;
            sr_2 <= sr_1;
            sr_3 <= sr_2;
            sr_4 <= sr_3;
            sr_5 <= sr_4;
            sr_6 <= sr_5;


        end
    end

always @( sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, a) begin
   case (a)
      3'd0: q = sr_0;
      3'd1: q = sr_1;
      3'd2: q = sr_2;
      3'd3: q = sr_3;
      3'd4: q = sr_4;
      3'd5: q = sr_5;
      3'd6: q = sr_6;
      default: q = sr_6;
   endcase
end

endmodule

module td_fused_top_fifo_w5_d7_S (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd5;
parameter ADDR_WIDTH  = 32'd3;
parameter DEPTH       = 4'd7;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 4'd1;
            if (mOutPtr == 4'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 4'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 4'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w5_d7_S_shiftReg 
U_td_fused_top_fifo_w5_d7_S_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w5_d7_S_x_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd5;
parameter ADDR_WIDTH = 32'd3;
parameter DEPTH = 4'd7;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;
            sr_2 <= sr_1;
            sr_3 <= sr_2;
            sr_4 <= sr_3;
            sr_5 <= sr_4;
            sr_6 <= sr_5;


        end
    end

always @( sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, a) begin
   case (a)
      3'd0: q = sr_0;
      3'd1: q = sr_1;
      3'd2: q = sr_2;
      3'd3: q = sr_3;
      3'd4: q = sr_4;
      3'd5: q = sr_5;
      3'd6: q = sr_6;
      default: q = sr_6;
   endcase
end

endmodule

module td_fused_top_fifo_w5_d7_S_x (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd5;
parameter ADDR_WIDTH  = 32'd3;
parameter DEPTH       = 4'd7;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 4'd1;
            if (mOutPtr == 4'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 4'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 4'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w5_d7_S_x_shiftReg 
U_td_fused_top_fifo_w5_d7_S_x_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w5_d8_S_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd5;
parameter ADDR_WIDTH = 32'd3;
parameter DEPTH = 4'd8;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, sr_7;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;
            sr_2 <= sr_1;
            sr_3 <= sr_2;
            sr_4 <= sr_3;
            sr_5 <= sr_4;
            sr_6 <= sr_5;
            sr_7 <= sr_6;


        end
    end

always @( sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, sr_7, a) begin
   case (a)
      3'd0: q = sr_0;
      3'd1: q = sr_1;
      3'd2: q = sr_2;
      3'd3: q = sr_3;
      3'd4: q = sr_4;
      3'd5: q = sr_5;
      3'd6: q = sr_6;
      3'd7: q = sr_7;
      default: q = sr_7;
   endcase
end

endmodule

module td_fused_top_fifo_w5_d8_S (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd5;
parameter ADDR_WIDTH  = 32'd3;
parameter DEPTH       = 4'd8;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 4'd1;
            if (mOutPtr == 4'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 4'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 4'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w5_d8_S_shiftReg 
U_td_fused_top_fifo_w5_d8_S_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w5_d8_S_x_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd5;
parameter ADDR_WIDTH = 32'd3;
parameter DEPTH = 4'd8;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, sr_7;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;
            sr_2 <= sr_1;
            sr_3 <= sr_2;
            sr_4 <= sr_3;
            sr_5 <= sr_4;
            sr_6 <= sr_5;
            sr_7 <= sr_6;


        end
    end

always @( sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, sr_7, a) begin
   case (a)
      3'd0: q = sr_0;
      3'd1: q = sr_1;
      3'd2: q = sr_2;
      3'd3: q = sr_3;
      3'd4: q = sr_4;
      3'd5: q = sr_5;
      3'd6: q = sr_6;
      3'd7: q = sr_7;
      default: q = sr_7;
   endcase
end

endmodule

module td_fused_top_fifo_w5_d8_S_x (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd5;
parameter ADDR_WIDTH  = 32'd3;
parameter DEPTH       = 4'd8;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 4'd1;
            if (mOutPtr == 4'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 4'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 4'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w5_d8_S_x_shiftReg 
U_td_fused_top_fifo_w5_d8_S_x_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w6_d2_S_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd6;
parameter ADDR_WIDTH = 32'd1;
parameter DEPTH = 2'd2;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;


        end
    end

always @( sr_0, sr_1, a) begin
   case (a)
      1'd0: q = sr_0;
      1'd1: q = sr_1;
      default: q = sr_1;
   endcase
end

endmodule

module td_fused_top_fifo_w6_d2_S (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd6;
parameter ADDR_WIDTH  = 32'd1;
parameter DEPTH       = 2'd2;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 2'd1;
            if (mOutPtr == 2'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 2'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 2'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w6_d2_S_shiftReg 
U_td_fused_top_fifo_w6_d2_S_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w6_d7_S_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd6;
parameter ADDR_WIDTH = 32'd3;
parameter DEPTH = 4'd7;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;
            sr_2 <= sr_1;
            sr_3 <= sr_2;
            sr_4 <= sr_3;
            sr_5 <= sr_4;
            sr_6 <= sr_5;


        end
    end

always @( sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, a) begin
   case (a)
      3'd0: q = sr_0;
      3'd1: q = sr_1;
      3'd2: q = sr_2;
      3'd3: q = sr_3;
      3'd4: q = sr_4;
      3'd5: q = sr_5;
      3'd6: q = sr_6;
      default: q = sr_6;
   endcase
end

endmodule

module td_fused_top_fifo_w6_d7_S (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd6;
parameter ADDR_WIDTH  = 32'd3;
parameter DEPTH       = 4'd7;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 4'd1;
            if (mOutPtr == 4'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 4'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 4'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w6_d7_S_shiftReg 
U_td_fused_top_fifo_w6_d7_S_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w6_d7_S_x_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd6;
parameter ADDR_WIDTH = 32'd3;
parameter DEPTH = 4'd7;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;
            sr_2 <= sr_1;
            sr_3 <= sr_2;
            sr_4 <= sr_3;
            sr_5 <= sr_4;
            sr_6 <= sr_5;


        end
    end

always @( sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, a) begin
   case (a)
      3'd0: q = sr_0;
      3'd1: q = sr_1;
      3'd2: q = sr_2;
      3'd3: q = sr_3;
      3'd4: q = sr_4;
      3'd5: q = sr_5;
      3'd6: q = sr_6;
      default: q = sr_6;
   endcase
end

endmodule

module td_fused_top_fifo_w6_d7_S_x (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd6;
parameter ADDR_WIDTH  = 32'd3;
parameter DEPTH       = 4'd7;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 4'd1;
            if (mOutPtr == 4'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 4'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 4'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w6_d7_S_x_shiftReg 
U_td_fused_top_fifo_w6_d7_S_x_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w6_d8_S_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd6;
parameter ADDR_WIDTH = 32'd3;
parameter DEPTH = 4'd8;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, sr_7;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;
            sr_2 <= sr_1;
            sr_3 <= sr_2;
            sr_4 <= sr_3;
            sr_5 <= sr_4;
            sr_6 <= sr_5;
            sr_7 <= sr_6;


        end
    end

always @( sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, sr_7, a) begin
   case (a)
      3'd0: q = sr_0;
      3'd1: q = sr_1;
      3'd2: q = sr_2;
      3'd3: q = sr_3;
      3'd4: q = sr_4;
      3'd5: q = sr_5;
      3'd6: q = sr_6;
      3'd7: q = sr_7;
      default: q = sr_7;
   endcase
end

endmodule

module td_fused_top_fifo_w6_d8_S (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd6;
parameter ADDR_WIDTH  = 32'd3;
parameter DEPTH       = 4'd8;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 4'd1;
            if (mOutPtr == 4'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 4'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 4'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w6_d8_S_shiftReg 
U_td_fused_top_fifo_w6_d8_S_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w6_d8_S_x_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd6;
parameter ADDR_WIDTH = 32'd3;
parameter DEPTH = 4'd8;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, sr_7;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;
            sr_2 <= sr_1;
            sr_3 <= sr_2;
            sr_4 <= sr_3;
            sr_5 <= sr_4;
            sr_6 <= sr_5;
            sr_7 <= sr_6;


        end
    end

always @( sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, sr_7, a) begin
   case (a)
      3'd0: q = sr_0;
      3'd1: q = sr_1;
      3'd2: q = sr_2;
      3'd3: q = sr_3;
      3'd4: q = sr_4;
      3'd5: q = sr_5;
      3'd6: q = sr_6;
      3'd7: q = sr_7;
      default: q = sr_7;
   endcase
end

endmodule

module td_fused_top_fifo_w6_d8_S_x (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd6;
parameter ADDR_WIDTH  = 32'd3;
parameter DEPTH       = 4'd8;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 4'd1;
            if (mOutPtr == 4'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 4'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 4'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w6_d8_S_x_shiftReg 
U_td_fused_top_fifo_w6_d8_S_x_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w7_d2_S_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd7;
parameter ADDR_WIDTH = 32'd1;
parameter DEPTH = 2'd2;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;


        end
    end

always @( sr_0, sr_1, a) begin
   case (a)
      1'd0: q = sr_0;
      1'd1: q = sr_1;
      default: q = sr_1;
   endcase
end

endmodule

module td_fused_top_fifo_w7_d2_S (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd7;
parameter ADDR_WIDTH  = 32'd1;
parameter DEPTH       = 2'd2;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 2'd1;
            if (mOutPtr == 2'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 2'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 2'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w7_d2_S_shiftReg 
U_td_fused_top_fifo_w7_d2_S_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w7_d2_S_x_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd7;
parameter ADDR_WIDTH = 32'd1;
parameter DEPTH = 2'd2;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;


        end
    end

always @( sr_0, sr_1, a) begin
   case (a)
      1'd0: q = sr_0;
      1'd1: q = sr_1;
      default: q = sr_1;
   endcase
end

endmodule

module td_fused_top_fifo_w7_d2_S_x (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd7;
parameter ADDR_WIDTH  = 32'd1;
parameter DEPTH       = 2'd2;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 2'd1;
            if (mOutPtr == 2'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 2'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 2'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w7_d2_S_x_shiftReg 
U_td_fused_top_fifo_w7_d2_S_x_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w7_d7_S_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd7;
parameter ADDR_WIDTH = 32'd3;
parameter DEPTH = 4'd7;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;
            sr_2 <= sr_1;
            sr_3 <= sr_2;
            sr_4 <= sr_3;
            sr_5 <= sr_4;
            sr_6 <= sr_5;


        end
    end

always @( sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, a) begin
   case (a)
      3'd0: q = sr_0;
      3'd1: q = sr_1;
      3'd2: q = sr_2;
      3'd3: q = sr_3;
      3'd4: q = sr_4;
      3'd5: q = sr_5;
      3'd6: q = sr_6;
      default: q = sr_6;
   endcase
end

endmodule

module td_fused_top_fifo_w7_d7_S (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd7;
parameter ADDR_WIDTH  = 32'd3;
parameter DEPTH       = 4'd7;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 4'd1;
            if (mOutPtr == 4'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 4'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 4'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w7_d7_S_shiftReg 
U_td_fused_top_fifo_w7_d7_S_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w7_d9_S_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd7;
parameter ADDR_WIDTH = 32'd4;
parameter DEPTH = 5'd9;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, sr_7, sr_8;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;
            sr_2 <= sr_1;
            sr_3 <= sr_2;
            sr_4 <= sr_3;
            sr_5 <= sr_4;
            sr_6 <= sr_5;
            sr_7 <= sr_6;
            sr_8 <= sr_7;


        end
    end

always @( sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, sr_7, sr_8, a) begin
   case (a)
      4'd0: q = sr_0;
      4'd1: q = sr_1;
      4'd2: q = sr_2;
      4'd3: q = sr_3;
      4'd4: q = sr_4;
      4'd5: q = sr_5;
      4'd6: q = sr_6;
      4'd7: q = sr_7;
      4'd8: q = sr_8;
      default: q = sr_8;
   endcase
end

endmodule

module td_fused_top_fifo_w7_d9_S (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd7;
parameter ADDR_WIDTH  = 32'd4;
parameter DEPTH       = 5'd9;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 5'd1;
            if (mOutPtr == 5'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 5'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 5'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w7_d9_S_shiftReg 
U_td_fused_top_fifo_w7_d9_S_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w8_d2_S_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd8;
parameter ADDR_WIDTH = 32'd1;
parameter DEPTH = 2'd2;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;


        end
    end

always @( sr_0, sr_1, a) begin
   case (a)
      1'd0: q = sr_0;
      1'd1: q = sr_1;
      default: q = sr_1;
   endcase
end

endmodule

module td_fused_top_fifo_w8_d2_S (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd8;
parameter ADDR_WIDTH  = 32'd1;
parameter DEPTH       = 2'd2;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 2'd1;
            if (mOutPtr == 2'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 2'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 2'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w8_d2_S_shiftReg 
U_td_fused_top_fifo_w8_d2_S_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w8_d2_S_x_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd8;
parameter ADDR_WIDTH = 32'd1;
parameter DEPTH = 2'd2;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;


        end
    end

always @( sr_0, sr_1, a) begin
   case (a)
      1'd0: q = sr_0;
      1'd1: q = sr_1;
      default: q = sr_1;
   endcase
end

endmodule

module td_fused_top_fifo_w8_d2_S_x (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd8;
parameter ADDR_WIDTH  = 32'd1;
parameter DEPTH       = 2'd2;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 2'd1;
            if (mOutPtr == 2'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 2'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 2'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w8_d2_S_x_shiftReg 
U_td_fused_top_fifo_w8_d2_S_x_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w8_d7_S_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd8;
parameter ADDR_WIDTH = 32'd3;
parameter DEPTH = 4'd7;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;
            sr_2 <= sr_1;
            sr_3 <= sr_2;
            sr_4 <= sr_3;
            sr_5 <= sr_4;
            sr_6 <= sr_5;


        end
    end

always @( sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, a) begin
   case (a)
      3'd0: q = sr_0;
      3'd1: q = sr_1;
      3'd2: q = sr_2;
      3'd3: q = sr_3;
      3'd4: q = sr_4;
      3'd5: q = sr_5;
      3'd6: q = sr_6;
      default: q = sr_6;
   endcase
end

endmodule

module td_fused_top_fifo_w8_d7_S (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd8;
parameter ADDR_WIDTH  = 32'd3;
parameter DEPTH       = 4'd7;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 4'd1;
            if (mOutPtr == 4'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 4'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 4'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w8_d7_S_shiftReg 
U_td_fused_top_fifo_w8_d7_S_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w8_d7_S_x0_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd8;
parameter ADDR_WIDTH = 32'd3;
parameter DEPTH = 4'd7;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;
            sr_2 <= sr_1;
            sr_3 <= sr_2;
            sr_4 <= sr_3;
            sr_5 <= sr_4;
            sr_6 <= sr_5;


        end
    end

always @( sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, a) begin
   case (a)
      3'd0: q = sr_0;
      3'd1: q = sr_1;
      3'd2: q = sr_2;
      3'd3: q = sr_3;
      3'd4: q = sr_4;
      3'd5: q = sr_5;
      3'd6: q = sr_6;
      default: q = sr_6;
   endcase
end

endmodule

module td_fused_top_fifo_w8_d7_S_x0 (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd8;
parameter ADDR_WIDTH  = 32'd3;
parameter DEPTH       = 4'd7;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 4'd1;
            if (mOutPtr == 4'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 4'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 4'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w8_d7_S_x0_shiftReg 
U_td_fused_top_fifo_w8_d7_S_x0_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w8_d7_S_x_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd8;
parameter ADDR_WIDTH = 32'd3;
parameter DEPTH = 4'd7;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;
            sr_2 <= sr_1;
            sr_3 <= sr_2;
            sr_4 <= sr_3;
            sr_5 <= sr_4;
            sr_6 <= sr_5;


        end
    end

always @( sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, a) begin
   case (a)
      3'd0: q = sr_0;
      3'd1: q = sr_1;
      3'd2: q = sr_2;
      3'd3: q = sr_3;
      3'd4: q = sr_4;
      3'd5: q = sr_5;
      3'd6: q = sr_6;
      default: q = sr_6;
   endcase
end

endmodule

module td_fused_top_fifo_w8_d7_S_x (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd8;
parameter ADDR_WIDTH  = 32'd3;
parameter DEPTH       = 4'd7;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 4'd1;
            if (mOutPtr == 4'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 4'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 4'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w8_d7_S_x_shiftReg 
U_td_fused_top_fifo_w8_d7_S_x_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w8_d8_S_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd8;
parameter ADDR_WIDTH = 32'd3;
parameter DEPTH = 4'd8;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, sr_7;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;
            sr_2 <= sr_1;
            sr_3 <= sr_2;
            sr_4 <= sr_3;
            sr_5 <= sr_4;
            sr_6 <= sr_5;
            sr_7 <= sr_6;


        end
    end

always @( sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, sr_7, a) begin
   case (a)
      3'd0: q = sr_0;
      3'd1: q = sr_1;
      3'd2: q = sr_2;
      3'd3: q = sr_3;
      3'd4: q = sr_4;
      3'd5: q = sr_5;
      3'd6: q = sr_6;
      3'd7: q = sr_7;
      default: q = sr_7;
   endcase
end

endmodule

module td_fused_top_fifo_w8_d8_S (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd8;
parameter ADDR_WIDTH  = 32'd3;
parameter DEPTH       = 4'd8;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 4'd1;
            if (mOutPtr == 4'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 4'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 4'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w8_d8_S_shiftReg 
U_td_fused_top_fifo_w8_d8_S_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w8_d8_S_x0_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd8;
parameter ADDR_WIDTH = 32'd3;
parameter DEPTH = 4'd8;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, sr_7;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;
            sr_2 <= sr_1;
            sr_3 <= sr_2;
            sr_4 <= sr_3;
            sr_5 <= sr_4;
            sr_6 <= sr_5;
            sr_7 <= sr_6;


        end
    end

always @( sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, sr_7, a) begin
   case (a)
      3'd0: q = sr_0;
      3'd1: q = sr_1;
      3'd2: q = sr_2;
      3'd3: q = sr_3;
      3'd4: q = sr_4;
      3'd5: q = sr_5;
      3'd6: q = sr_6;
      3'd7: q = sr_7;
      default: q = sr_7;
   endcase
end

endmodule

module td_fused_top_fifo_w8_d8_S_x0 (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd8;
parameter ADDR_WIDTH  = 32'd3;
parameter DEPTH       = 4'd8;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 4'd1;
            if (mOutPtr == 4'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 4'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 4'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w8_d8_S_x0_shiftReg 
U_td_fused_top_fifo_w8_d8_S_x0_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w8_d8_S_x_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd8;
parameter ADDR_WIDTH = 32'd3;
parameter DEPTH = 4'd8;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, sr_7;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;
            sr_2 <= sr_1;
            sr_3 <= sr_2;
            sr_4 <= sr_3;
            sr_5 <= sr_4;
            sr_6 <= sr_5;
            sr_7 <= sr_6;


        end
    end

always @( sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, sr_7, a) begin
   case (a)
      3'd0: q = sr_0;
      3'd1: q = sr_1;
      3'd2: q = sr_2;
      3'd3: q = sr_3;
      3'd4: q = sr_4;
      3'd5: q = sr_5;
      3'd6: q = sr_6;
      3'd7: q = sr_7;
      default: q = sr_7;
   endcase
end

endmodule

module td_fused_top_fifo_w8_d8_S_x (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd8;
parameter ADDR_WIDTH  = 32'd3;
parameter DEPTH       = 4'd8;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 4'd1;
            if (mOutPtr == 4'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 4'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 4'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w8_d8_S_x_shiftReg 
U_td_fused_top_fifo_w8_d8_S_x_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w9_d2_S_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd9;
parameter ADDR_WIDTH = 32'd1;
parameter DEPTH = 2'd2;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;


        end
    end

always @( sr_0, sr_1, a) begin
   case (a)
      1'd0: q = sr_0;
      1'd1: q = sr_1;
      default: q = sr_1;
   endcase
end

endmodule

module td_fused_top_fifo_w9_d2_S (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd9;
parameter ADDR_WIDTH  = 32'd1;
parameter DEPTH       = 2'd2;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 2'd1;
            if (mOutPtr == 2'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 2'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 2'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w9_d2_S_shiftReg 
U_td_fused_top_fifo_w9_d2_S_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w9_d2_S_x_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd9;
parameter ADDR_WIDTH = 32'd1;
parameter DEPTH = 2'd2;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;


        end
    end

always @( sr_0, sr_1, a) begin
   case (a)
      1'd0: q = sr_0;
      1'd1: q = sr_1;
      default: q = sr_1;
   endcase
end

endmodule

module td_fused_top_fifo_w9_d2_S_x (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd9;
parameter ADDR_WIDTH  = 32'd1;
parameter DEPTH       = 2'd2;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 2'd1;
            if (mOutPtr == 2'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 2'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 2'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w9_d2_S_x_shiftReg 
U_td_fused_top_fifo_w9_d2_S_x_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_fifo_w9_d7_S_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd9;
parameter ADDR_WIDTH = 32'd3;
parameter DEPTH = 4'd7;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;
            sr_2 <= sr_1;
            sr_3 <= sr_2;
            sr_4 <= sr_3;
            sr_5 <= sr_4;
            sr_6 <= sr_5;


        end
    end

always @( sr_0, sr_1, sr_2, sr_3, sr_4, sr_5, sr_6, a) begin
   case (a)
      3'd0: q = sr_0;
      3'd1: q = sr_1;
      3'd2: q = sr_2;
      3'd3: q = sr_3;
      3'd4: q = sr_4;
      3'd5: q = sr_5;
      3'd6: q = sr_6;
      default: q = sr_6;
   endcase
end

endmodule

module td_fused_top_fifo_w9_d7_S (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd9;
parameter ADDR_WIDTH  = 32'd3;
parameter DEPTH       = 4'd7;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 4'd1;
            if (mOutPtr == 4'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 4'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 4'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_fifo_w9_d7_S_shiftReg 
U_td_fused_top_fifo_w9_d7_S_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_ap_hadd_3_full_dsp_16 (
   input  wire        aclk,
   input wire         aclken,
   input  wire        s_axis_a_tvalid,
   input  wire [15:0] s_axis_a_tdata,
   input  wire        s_axis_b_tvalid,
   input  wire [15:0] s_axis_b_tdata,
   output wire        m_axis_result_tvalid,
   output wire [15:0] m_axis_result_tdata
);
    wire res;
   reg [15:0] a_reg, b_reg, res_reg;

   always @(posedge aclk) begin
      if (aclken) begin
         a_reg <= s_axis_a_tdata;     
         b_reg <= s_axis_b_tdata;     
         res_reg <= res;
      end
   end


`ifdef complex_dsp
   adder_fp u_add_fp (
      .a(a_reg), 
      .b(b_reg), 
      .out(res)
   );
`else
FPAddSub u_FPAddSub (.clk(), .rst(1'b0), .a(a_reg), .b(b_reg), .operation(1'b0), .result(res), .flags());
`endif


   assign m_axis_result_tdata = res_reg;

endmodule


module td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1
#(parameter
    ID         = 25,
    NUM_STAGE  = 5,
    din0_WIDTH = 16,
    din1_WIDTH = 16,
    dout_WIDTH = 16
)(
    input  wire                  clk,
    input  wire                  reset,
    input  wire                  ce,
    input  wire [din0_WIDTH-1:0] din0,
    input  wire [din1_WIDTH-1:0] din1,
    output wire [dout_WIDTH-1:0] dout
);
//------------------------Local signal-------------------
wire                  aclk;
wire                  aclken;
wire                  a_tvalid;
wire [15:0]           a_tdata;
wire                  b_tvalid;
wire [15:0]           b_tdata;
wire                  r_tvalid;
wire [15:0]           r_tdata;
reg  [din0_WIDTH-1:0] din0_buf1;
reg  [din1_WIDTH-1:0] din1_buf1;
reg                   ce_r;
wire [dout_WIDTH-1:0] dout_i;
reg  [dout_WIDTH-1:0] dout_r;
//------------------------Instantiation------------------
td_fused_top_ap_hadd_3_full_dsp_16 td_fused_top_ap_hadd_3_full_dsp_16_u (
    .aclk                 ( aclk ),
    .aclken               ( aclken ),
    .s_axis_a_tvalid      ( a_tvalid ),
    .s_axis_a_tdata       ( a_tdata ),
    .s_axis_b_tvalid      ( b_tvalid ),
    .s_axis_b_tdata       ( b_tdata ),
    .m_axis_result_tvalid ( r_tvalid ),
    .m_axis_result_tdata  ( r_tdata )
);
//------------------------Body---------------------------
assign aclk     = clk;
assign aclken   = ce_r;
assign a_tvalid = 1'b1;
assign a_tdata  = din0_buf1;
assign b_tvalid = 1'b1;
assign b_tdata  = din1_buf1;
assign dout_i   = r_tdata;

always @(posedge clk) begin
    if (ce) begin
        din0_buf1 <= din0;
        din1_buf1 <= din1;
    end
end

always @ (posedge clk) begin
    ce_r <= ce;
end

always @ (posedge clk) begin
    if (ce_r) begin
        dout_r <= dout_i;
    end
end

assign dout = ce_r?dout_i:dout_r;
endmodule
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_ap_hcmp_0_no_dsp_16 (
   input  wire        s_axis_a_tvalid,
   input  wire [15:0] s_axis_a_tdata,
   input  wire        s_axis_b_tvalid,
   input  wire [15:0] s_axis_b_tdata,
   input  wire        s_axis_operation_tvalid,
   input  wire [7:0]  s_axis_operation_tdata,
   output wire        m_axis_result_tvalid,
   output wire [7:0]  m_axis_result_tdata
);
   // TEMP - compare module not yet ready
   // In the meantime, negate operand B, add them
   // together, and return the sign bit of the result.
   wire [15:0] b_negative;
   wire [15:0] result;
   assign b_negative = {~s_axis_b_tdata[15], s_axis_b_tdata[14:0]};
   
`ifdef complex_dsp
adder_fp u_add_fp (
      .a(s_axis_a_tdata), 
      .b(b_negative), 
      .out(result)
   );
`else
FPAddSub u_FPAddSub_2 (.clk(), .rst(1'b0), .a(s_axis_a_tdata), .b(b_negative), .operation(1'b0), .result(result), .flags());
`endif
   
   assign m_axis_result_tdata = {7'b0, result[15]};
endmodule

module td_fused_top_hcmp_16ns_16ns_1_2_no_dsp_1
#(parameter
    ID         = 47,
    NUM_STAGE  = 2,
    din0_WIDTH = 16,
    din1_WIDTH = 16,
    dout_WIDTH = 1
)(
    input  wire                  clk,
    input  wire                  reset,
    input  wire                  ce,
    input  wire [din0_WIDTH-1:0] din0,
    input  wire [din1_WIDTH-1:0] din1,
    input  wire [4:0]            opcode,
    output wire [dout_WIDTH-1:0] dout
);
//------------------------Parameter----------------------
// AutoESL opcode
localparam [4:0]
    AP_OEQ = 5'b00001,
    AP_OGT = 5'b00010,
    AP_OGE = 5'b00011,
    AP_OLT = 5'b00100,
    AP_OLE = 5'b00101,
    AP_ONE = 5'b00110,
    AP_UNO = 5'b01000;
// FPV6 opcode
localparam [7:0]
    OP_EQ = 8'b00010100,
    OP_GT = 8'b00100100,
    OP_GE = 8'b00110100,
    OP_LT = 8'b00001100,
    OP_LE = 8'b00011100,
    OP_NE = 8'b00101100,
    OP_UO = 8'b00000100;
//------------------------Local signal-------------------
wire                  a_tvalid;
wire [15:0]           a_tdata;
wire                  b_tvalid;
wire [15:0]           b_tdata;
wire                  op_tvalid;
reg  [7:0]            op_tdata;
wire                  r_tvalid;
wire [7:0]            r_tdata;
reg  [din0_WIDTH-1:0] din0_buf1;
reg  [din1_WIDTH-1:0] din1_buf1;
reg  [4:0]            opcode_buf1;
reg                   ce_r;
wire [dout_WIDTH-1:0] dout_i;
reg  [dout_WIDTH-1:0] dout_r;
//------------------------Instantiation------------------
td_fused_top_ap_hcmp_0_no_dsp_16 td_fused_top_ap_hcmp_0_no_dsp_16_u (
    .s_axis_a_tvalid         ( a_tvalid ),
    .s_axis_a_tdata          ( a_tdata ),
    .s_axis_b_tvalid         ( b_tvalid ),
    .s_axis_b_tdata          ( b_tdata ),
    .s_axis_operation_tvalid ( op_tvalid ),
    .s_axis_operation_tdata  ( op_tdata ),
    .m_axis_result_tvalid    ( r_tvalid ),
    .m_axis_result_tdata     ( r_tdata )
);
//------------------------Body---------------------------
assign a_tvalid  = 1'b1;
assign a_tdata   = din0_buf1;
assign b_tvalid  = 1'b1;
assign b_tdata   = din1_buf1;
assign op_tvalid = 1'b1;
assign dout_i    = r_tdata[0];

always @(*) begin
    case (opcode_buf1)
        AP_OEQ  : op_tdata = OP_EQ;
        AP_OGT  : op_tdata = OP_GT;
        AP_OGE  : op_tdata = OP_GE;
        AP_OLT  : op_tdata = OP_LT;
        AP_OLE  : op_tdata = OP_LE;
        AP_ONE  : op_tdata = OP_NE;
        AP_UNO  : op_tdata = OP_UO;
        default : op_tdata = OP_EQ;
    endcase
end

always @(posedge clk) begin
    if (ce) begin
        din0_buf1   <= din0;
        din1_buf1   <= din1;
        opcode_buf1 <= opcode;
    end
end

always @ (posedge clk) begin
    ce_r <= ce;
end

always @ (posedge clk) begin
    if (ce_r) begin
        dout_r <= dout_i;
    end
end

assign dout = ce_r?dout_i:dout_r;
endmodule
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_ap_hmul_2_max_dsp_16 (
   input  wire        aclk,
   input  wire        aclken,
   input  wire        s_axis_a_tvalid,
   input  wire [15:0] s_axis_a_tdata,
   input  wire        s_axis_b_tvalid,
   input  wire [15:0] s_axis_b_tdata,
   output wire        m_axis_result_tvalid,
   output wire [15:0] m_axis_result_tdata
);
   
   wire res;
   reg [15:0] a_reg, b_reg, res_reg;

   always @(posedge aclk) begin
      if (aclken) begin
         a_reg <= s_axis_a_tdata;     
         b_reg <= s_axis_b_tdata;     
         res_reg <= res;
      end
   end

`ifdef complex_dsp
   multiply_fp u_mult_fp (
      .a(a_reg), 
      .b(b_reg), 
      .out(res)
   );
`else
FPMult_16 u_FPMult (.clk(), .rst(1'b0), .a(a_reg), .b(b_reg), .result(res), .flags());
`endif
   assign m_axis_result_tdata = res_reg;

endmodule


module td_fused_top_hmul_16ns_16ns_16_4_max_dsp_1
#(parameter
    ID         = 20,
    NUM_STAGE  = 4,
    din0_WIDTH = 16,
    din1_WIDTH = 16,
    dout_WIDTH = 16
)(
    input  wire                  clk,
    input  wire                  reset,
    input  wire                  ce,
    input  wire [din0_WIDTH-1:0] din0,
    input  wire [din1_WIDTH-1:0] din1,
    output wire [dout_WIDTH-1:0] dout
);
//------------------------Local signal-------------------
wire                  aclk;
wire                  aclken;
wire                  a_tvalid;
wire [15:0]           a_tdata;
wire                  b_tvalid;
wire [15:0]           b_tdata;
wire                  r_tvalid;
wire [15:0]           r_tdata;
reg  [din0_WIDTH-1:0] din0_buf1;
reg  [din1_WIDTH-1:0] din1_buf1;
reg                   ce_r;
wire [dout_WIDTH-1:0] dout_i;
reg  [dout_WIDTH-1:0] dout_r;
//------------------------Instantiation------------------
td_fused_top_ap_hmul_2_max_dsp_16 td_fused_top_ap_hmul_2_max_dsp_16_u (
    .aclk                 ( aclk ),
    .aclken               ( aclken ),
    .s_axis_a_tvalid      ( a_tvalid ),
    .s_axis_a_tdata       ( a_tdata ),
    .s_axis_b_tvalid      ( b_tvalid ),
    .s_axis_b_tdata       ( b_tdata ),
    .m_axis_result_tvalid ( r_tvalid ),
    .m_axis_result_tdata  ( r_tdata )
);
//------------------------Body---------------------------
assign aclk     = clk;
assign aclken   = ce_r;
assign a_tvalid = 1'b1;
assign a_tdata  = din0_buf1;
assign b_tvalid = 1'b1;
assign b_tdata  = din1_buf1;
assign dout_i   = r_tdata;

always @(posedge clk) begin
    if (ce) begin
        din0_buf1 <= din0;
        din1_buf1 <= din1;
    end
end

always @ (posedge clk) begin
    ce_r <= ce;
end

always @ (posedge clk) begin
    if (ce_r) begin
        dout_r <= dout_i;
    end
end

assign dout = ce_r?dout_i:dout_r;
endmodule
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_hsub_16ns_16ns_16_5_full_dsp_1
#(parameter
    ID         = 37,
    NUM_STAGE  = 5,
    din0_WIDTH = 16,
    din1_WIDTH = 16,
    dout_WIDTH = 16
)(
    input  wire                  clk,
    input  wire                  reset,
    input  wire                  ce,
    input  wire [din0_WIDTH-1:0] din0,
    input  wire [din1_WIDTH-1:0] din1,
    output wire [dout_WIDTH-1:0] dout
);
//------------------------Local signal-------------------
wire                  aclk;
wire                  aclken;
wire                  a_tvalid;
wire [15:0]           a_tdata;
wire                  b_tvalid;
wire [15:0]           b_tdata;
wire                  r_tvalid;
wire [15:0]           r_tdata;
reg  [din0_WIDTH-1:0] din0_buf1;
reg  [din1_WIDTH-1:0] din1_buf1;
reg                   ce_r;
wire [dout_WIDTH-1:0] dout_i;
reg  [dout_WIDTH-1:0] dout_r;
//------------------------Instantiation------------------
// Just replace with the hadd, logic is similar enough.
//td_fused_top_ap_hsub_3_full_dsp_16 td_fused_top_ap_hsub_3_full_dsp_16_u (
td_fused_top_ap_hadd_3_full_dsp_16 td_fused_top_ap_hsub_3_full_dsp_16_u (
    .aclk                 ( aclk ),
    .aclken               ( aclken ),
    .s_axis_a_tvalid      ( a_tvalid ),
    .s_axis_a_tdata       ( a_tdata ),
    .s_axis_b_tvalid      ( b_tvalid ),
    .s_axis_b_tdata       ( b_tdata ),
    .m_axis_result_tvalid ( r_tvalid ),
    .m_axis_result_tdata  ( r_tdata )
);
//------------------------Body---------------------------
assign aclk     = clk;
assign aclken   = ce_r;
assign a_tvalid = 1'b1;
assign a_tdata  = din0_buf1;
assign b_tvalid = 1'b1;
assign b_tdata  = din1_buf1;
assign dout_i   = r_tdata;

always @(posedge clk) begin
    if (ce) begin
        din0_buf1 <= din0;
        din1_buf1 <= din1;
    end
end

always @ (posedge clk) begin
    ce_r <= ce;
end

always @ (posedge clk) begin
    if (ce_r) begin
        dout_r <= dout_i;
    end
end

assign dout = ce_r?dout_i:dout_r;
endmodule
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps

  module td_fused_top_mac_muladd_10s_9ns_8ns_16_4_1_DSP48_0(
    input clk,
    input rst,
    input ce,
    input  [10 - 1:0] in0,
    input  [9 - 1:0] in1,
    input  [8 - 1:0] in2,
    output [16 - 1:0]  dout);

wire  [27 - 1:0]     a;
wire  [18 - 1:0]     b;
wire  [48 - 1:0]     c;
wire  [45 - 1:0]     m;
wire  [48 - 1:0]     p;
reg   [45 - 1:0]     m_reg;
reg   [27 - 1:0]     a_reg;
reg   [18 - 1:0]     b_reg;
reg   [48 - 1:0]     p_reg;

assign a  = (in0);
assign b  = (in1);
assign c  = (in2);

assign m  = a_reg * b_reg;
assign p  = m_reg + c;

always @(posedge clk) begin
    if (ce) begin
        m_reg  <= m;
        a_reg  <= a;
        b_reg  <= b;
        p_reg  <= p;
    end
end

assign dout = p_reg;

endmodule
`timescale 1 ns / 1 ps
module td_fused_top_mac_muladd_10s_9ns_8ns_16_4_1(
    clk,
    reset,
    ce,
    din0,
    din1,
    din2,
    dout);

parameter ID = 32'd1;
parameter NUM_STAGE = 32'd1;
parameter din0_WIDTH = 32'd1;
parameter din1_WIDTH = 32'd1;
parameter din2_WIDTH = 32'd1;
parameter dout_WIDTH = 32'd1;
input clk;
input reset;
input ce;
input[din0_WIDTH - 1:0] din0;
input[din1_WIDTH - 1:0] din1;
input[din2_WIDTH - 1:0] din2;
output[dout_WIDTH - 1:0] dout;



td_fused_top_mac_muladd_10s_9ns_8ns_16_4_1_DSP48_0 td_fused_top_mac_muladd_10s_9ns_8ns_16_4_1_DSP48_0_U(
    .clk( clk ),
    .rst( reset ),
    .ce( ce ),
    .in0( din0 ),
    .in1( din1 ),
    .in2( din2 ),
    .dout( dout )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_mul_10s_9ns_16_1_1_Multiplier_0(a, b, p);
input[10 - 1 : 0] a; 
input[9 - 1 : 0] b; 
output[16 - 1 : 0] p;

assign p = (a) * ({1'b0, b});
endmodule
`timescale 1 ns / 1 ps
module td_fused_top_mul_10s_9ns_16_1_1(
    din0,
    din1,
    dout);

parameter ID = 32'd1;
parameter NUM_STAGE = 32'd1;
parameter din0_WIDTH = 32'd1;
parameter din1_WIDTH = 32'd1;
parameter dout_WIDTH = 32'd1;
input[din0_WIDTH - 1:0] din0;
input[din1_WIDTH - 1:0] din1;
output[dout_WIDTH - 1:0] dout;



td_fused_top_mul_10s_9ns_16_1_1_Multiplier_0 td_fused_top_mul_10s_9ns_16_1_1_Multiplier_0_U(
    .a( din0 ),
    .b( din1 ),
    .p( dout )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_regslice_both
#(parameter 
    DataWidth=32
)(
    input ap_clk ,
    input ap_rst,

    input [DataWidth-1:0] data_in , 
    input vld_in , 
    output ack_in ,
    output [DataWidth-1:0] data_out, 
    output vld_out,
    input ack_out,
    output apdone_blk
);
 

reg   [1:0] B_V_data_1_state;
wire   [DataWidth-1:0] B_V_data_1_data_in;
reg   [DataWidth-1:0] B_V_data_1_data_out;
wire    B_V_data_1_vld_reg;
wire    B_V_data_1_vld_in;
wire    B_V_data_1_vld_out;
reg   [DataWidth-1:0] B_V_data_1_payload_A;
reg   [DataWidth-1:0] B_V_data_1_payload_B;
reg    B_V_data_1_sel_rd;
reg    B_V_data_1_sel_wr;
wire    B_V_data_1_sel;
wire    B_V_data_1_load_A;
wire    B_V_data_1_load_B;
wire    B_V_data_1_state_cmp_full;
wire    B_V_data_1_ack_in;
wire    B_V_data_1_ack_out;

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        B_V_data_1_sel_rd <= 1'b0;
    end else begin
        if (((1'b1 == B_V_data_1_vld_out) & (1'b1 == B_V_data_1_ack_out))) begin
            B_V_data_1_sel_rd <= ~B_V_data_1_sel_rd;
        end else begin
            B_V_data_1_sel_rd <= B_V_data_1_sel_rd;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        B_V_data_1_sel_wr <= 1'b0;
    end else begin
        if (((1'b1 == B_V_data_1_vld_in) & (1'b1 == B_V_data_1_ack_in))) begin
            B_V_data_1_sel_wr <= ~B_V_data_1_sel_wr;
        end else begin
            B_V_data_1_sel_wr <= B_V_data_1_sel_wr;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        B_V_data_1_state <= 2'd0;
    end else begin
        if ((((2'd3 == B_V_data_1_state) & (1'b0 == B_V_data_1_vld_in) & (1'b1 == B_V_data_1_ack_out)) | ((2'd2 == B_V_data_1_state) & (1'b0 == B_V_data_1_vld_in)))) begin
            B_V_data_1_state <= 2'd2;
        end else if ((((2'd1 == B_V_data_1_state) & (1'b0 == B_V_data_1_ack_out)) | ((2'd3 == B_V_data_1_state) & (1'b0 == B_V_data_1_ack_out) & (1'b1 == B_V_data_1_vld_in)))) begin
            B_V_data_1_state <= 2'd1;
        end else if ((((2'd1 == B_V_data_1_state) & (1'b1 == B_V_data_1_ack_out)) | (~((1'b0 == B_V_data_1_ack_out) & (1'b1 == B_V_data_1_vld_in)) & ~((1'b0 == B_V_data_1_vld_in) & (1'b1 == B_V_data_1_ack_out)) & (2'd3 == B_V_data_1_state)) | ((2'd2 == B_V_data_1_state) & (1'b1 == B_V_data_1_vld_in)))) begin
            B_V_data_1_state <= 2'd3;
        end else begin
            B_V_data_1_state <= 2'd2;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == B_V_data_1_load_A)) begin
        B_V_data_1_payload_A <= B_V_data_1_data_in;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == B_V_data_1_load_B)) begin
        B_V_data_1_payload_B <= B_V_data_1_data_in;
    end
end

always @ (*) begin
    if ((1'b1 == B_V_data_1_sel)) begin
        B_V_data_1_data_out = B_V_data_1_payload_B;
    end else begin
        B_V_data_1_data_out = B_V_data_1_payload_A;
    end
end

assign B_V_data_1_ack_in = B_V_data_1_state[1'd1];
assign B_V_data_1_load_A = (~B_V_data_1_sel_wr & B_V_data_1_state_cmp_full);
assign B_V_data_1_load_B = (B_V_data_1_state_cmp_full & B_V_data_1_sel_wr);
assign B_V_data_1_sel = B_V_data_1_sel_rd;
assign B_V_data_1_state_cmp_full = ((B_V_data_1_state != 2'd1) ? 1'b1 : 1'b0);
assign B_V_data_1_vld_out = B_V_data_1_state[1'd0];

assign ack_in = B_V_data_1_ack_in;
assign B_V_data_1_data_in = data_in;
assign B_V_data_1_vld_in = vld_in;

assign vld_out = B_V_data_1_vld_out;
assign data_out = B_V_data_1_data_out;
assign B_V_data_1_ack_out = ack_out;

assign apdone_blk = ((B_V_data_1_state == 2'd3 && ack_out == 1'b0) | (B_V_data_1_state == 2'd1));

endmodule // both



// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_start_for_tdf10_readFilters68_U0_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd1;
parameter ADDR_WIDTH = 32'd1;
parameter DEPTH = 2'd2;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;


        end
    end

always @( sr_0, sr_1, a) begin
   case (a)
      1'd0: q = sr_0;
      1'd1: q = sr_1;
      default: q = sr_1;
   endcase
end

endmodule

module td_fused_top_start_for_tdf10_readFilters68_U0 (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd1;
parameter ADDR_WIDTH  = 32'd1;
parameter DEPTH       = 2'd2;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 2'd1;
            if (mOutPtr == 2'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 2'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 2'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_start_for_tdf10_readFilters68_U0_shiftReg 
U_td_fused_top_start_for_tdf10_readFilters68_U0_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_start_for_tdf11_readFilters74_U0_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd1;
parameter ADDR_WIDTH = 32'd1;
parameter DEPTH = 2'd2;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;


        end
    end

always @( sr_0, sr_1, a) begin
   case (a)
      1'd0: q = sr_0;
      1'd1: q = sr_1;
      default: q = sr_1;
   endcase
end

endmodule

module td_fused_top_start_for_tdf11_readFilters74_U0 (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd1;
parameter ADDR_WIDTH  = 32'd1;
parameter DEPTH       = 2'd2;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 2'd1;
            if (mOutPtr == 2'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 2'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 2'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_start_for_tdf11_readFilters74_U0_shiftReg 
U_td_fused_top_start_for_tdf11_readFilters74_U0_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_start_for_tdf12_readFilters78_U0_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd1;
parameter ADDR_WIDTH = 32'd1;
parameter DEPTH = 2'd2;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;


        end
    end

always @( sr_0, sr_1, a) begin
   case (a)
      1'd0: q = sr_0;
      1'd1: q = sr_1;
      default: q = sr_1;
   endcase
end

endmodule

module td_fused_top_start_for_tdf12_readFilters78_U0 (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd1;
parameter ADDR_WIDTH  = 32'd1;
parameter DEPTH       = 2'd2;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 2'd1;
            if (mOutPtr == 2'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 2'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 2'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_start_for_tdf12_readFilters78_U0_shiftReg 
U_td_fused_top_start_for_tdf12_readFilters78_U0_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_start_for_tdf1_readFilters18_U0_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd1;
parameter ADDR_WIDTH = 32'd1;
parameter DEPTH = 2'd2;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;


        end
    end

always @( sr_0, sr_1, a) begin
   case (a)
      1'd0: q = sr_0;
      1'd1: q = sr_1;
      default: q = sr_1;
   endcase
end

endmodule

module td_fused_top_start_for_tdf1_readFilters18_U0 (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd1;
parameter ADDR_WIDTH  = 32'd1;
parameter DEPTH       = 2'd2;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 2'd1;
            if (mOutPtr == 2'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 2'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 2'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_start_for_tdf1_readFilters18_U0_shiftReg 
U_td_fused_top_start_for_tdf1_readFilters18_U0_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_start_for_tdf2_readFilters24_U0_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd1;
parameter ADDR_WIDTH = 32'd1;
parameter DEPTH = 2'd2;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;


        end
    end

always @( sr_0, sr_1, a) begin
   case (a)
      1'd0: q = sr_0;
      1'd1: q = sr_1;
      default: q = sr_1;
   endcase
end

endmodule

module td_fused_top_start_for_tdf2_readFilters24_U0 (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd1;
parameter ADDR_WIDTH  = 32'd1;
parameter DEPTH       = 2'd2;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 2'd1;
            if (mOutPtr == 2'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 2'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 2'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_start_for_tdf2_readFilters24_U0_shiftReg 
U_td_fused_top_start_for_tdf2_readFilters24_U0_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_start_for_tdf3_readFilters30_U0_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd1;
parameter ADDR_WIDTH = 32'd1;
parameter DEPTH = 2'd2;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;


        end
    end

always @( sr_0, sr_1, a) begin
   case (a)
      1'd0: q = sr_0;
      1'd1: q = sr_1;
      default: q = sr_1;
   endcase
end

endmodule

module td_fused_top_start_for_tdf3_readFilters30_U0 (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd1;
parameter ADDR_WIDTH  = 32'd1;
parameter DEPTH       = 2'd2;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 2'd1;
            if (mOutPtr == 2'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 2'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 2'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_start_for_tdf3_readFilters30_U0_shiftReg 
U_td_fused_top_start_for_tdf3_readFilters30_U0_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_start_for_tdf4_readFilters36_U0_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd1;
parameter ADDR_WIDTH = 32'd1;
parameter DEPTH = 2'd2;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;


        end
    end

always @( sr_0, sr_1, a) begin
   case (a)
      1'd0: q = sr_0;
      1'd1: q = sr_1;
      default: q = sr_1;
   endcase
end

endmodule

module td_fused_top_start_for_tdf4_readFilters36_U0 (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd1;
parameter ADDR_WIDTH  = 32'd1;
parameter DEPTH       = 2'd2;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 2'd1;
            if (mOutPtr == 2'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 2'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 2'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_start_for_tdf4_readFilters36_U0_shiftReg 
U_td_fused_top_start_for_tdf4_readFilters36_U0_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_start_for_tdf5_readFilters40_U0_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd1;
parameter ADDR_WIDTH = 32'd1;
parameter DEPTH = 2'd2;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;


        end
    end

always @( sr_0, sr_1, a) begin
   case (a)
      1'd0: q = sr_0;
      1'd1: q = sr_1;
      default: q = sr_1;
   endcase
end

endmodule

module td_fused_top_start_for_tdf5_readFilters40_U0 (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd1;
parameter ADDR_WIDTH  = 32'd1;
parameter DEPTH       = 2'd2;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 2'd1;
            if (mOutPtr == 2'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 2'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 2'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_start_for_tdf5_readFilters40_U0_shiftReg 
U_td_fused_top_start_for_tdf5_readFilters40_U0_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_start_for_tdf6_readFilters46_U0_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd1;
parameter ADDR_WIDTH = 32'd1;
parameter DEPTH = 2'd2;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;


        end
    end

always @( sr_0, sr_1, a) begin
   case (a)
      1'd0: q = sr_0;
      1'd1: q = sr_1;
      default: q = sr_1;
   endcase
end

endmodule

module td_fused_top_start_for_tdf6_readFilters46_U0 (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd1;
parameter ADDR_WIDTH  = 32'd1;
parameter DEPTH       = 2'd2;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 2'd1;
            if (mOutPtr == 2'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 2'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 2'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_start_for_tdf6_readFilters46_U0_shiftReg 
U_td_fused_top_start_for_tdf6_readFilters46_U0_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_start_for_tdf7_readFilters52_U0_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd1;
parameter ADDR_WIDTH = 32'd1;
parameter DEPTH = 2'd2;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;


        end
    end

always @( sr_0, sr_1, a) begin
   case (a)
      1'd0: q = sr_0;
      1'd1: q = sr_1;
      default: q = sr_1;
   endcase
end

endmodule

module td_fused_top_start_for_tdf7_readFilters52_U0 (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd1;
parameter ADDR_WIDTH  = 32'd1;
parameter DEPTH       = 2'd2;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 2'd1;
            if (mOutPtr == 2'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 2'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 2'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_start_for_tdf7_readFilters52_U0_shiftReg 
U_td_fused_top_start_for_tdf7_readFilters52_U0_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_start_for_tdf8_readFilters56_U0_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd1;
parameter ADDR_WIDTH = 32'd1;
parameter DEPTH = 2'd2;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;


        end
    end

always @( sr_0, sr_1, a) begin
   case (a)
      1'd0: q = sr_0;
      1'd1: q = sr_1;
      default: q = sr_1;
   endcase
end

endmodule

module td_fused_top_start_for_tdf8_readFilters56_U0 (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd1;
parameter ADDR_WIDTH  = 32'd1;
parameter DEPTH       = 2'd2;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 2'd1;
            if (mOutPtr == 2'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 2'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 2'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_start_for_tdf8_readFilters56_U0_shiftReg 
U_td_fused_top_start_for_tdf8_readFilters56_U0_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module td_fused_top_start_for_tdf9_readFilters62_U0_shiftReg (
    clk,
    data,
    ce,
    a,
    q);

parameter DATA_WIDTH = 32'd1;
parameter ADDR_WIDTH = 32'd1;
parameter DEPTH = 2'd2;

input clk;
input [DATA_WIDTH-1:0] data;
input ce;
input [ADDR_WIDTH-1:0] a;
output reg [DATA_WIDTH-1:0] q;

reg[DATA_WIDTH-1:0] sr_0, sr_1;
integer i;

always @ (posedge clk)
    begin
        if (ce)
        begin
            sr_0 <= data;
            sr_1 <= sr_0;


        end
    end

always @( sr_0, sr_1, a) begin
   case (a)
      1'd0: q = sr_0;
      1'd1: q = sr_1;
      default: q = sr_1;
   endcase
end

endmodule

module td_fused_top_start_for_tdf9_readFilters62_U0 (
    clk,
    reset,
    if_empty_n,
    if_read_ce,
    if_read,
    if_dout,
    if_full_n,
    if_write_ce,
    if_write,
    if_din);

parameter MEM_STYLE   = "shiftreg";
parameter DATA_WIDTH  = 32'd1;
parameter ADDR_WIDTH  = 32'd1;
parameter DEPTH       = 2'd2;

input clk;
input reset;
output if_empty_n;
input if_read_ce;
input if_read;
output[DATA_WIDTH - 1:0] if_dout;
output if_full_n;
input if_write_ce;
input if_write;
input[DATA_WIDTH - 1:0] if_din;

wire[ADDR_WIDTH - 1:0] shiftReg_addr ;
wire[DATA_WIDTH - 1:0] shiftReg_data, shiftReg_q;
wire                     shiftReg_ce;
reg[ADDR_WIDTH:0] mOutPtr = ~{(ADDR_WIDTH+1){1'b0}};
reg internal_empty_n = 0;
reg internal_full_n = 1;

assign if_full_n = internal_full_n;
assign if_empty_n = internal_empty_n;
assign shiftReg_data = if_din;
assign if_dout = shiftReg_q;

always @ (posedge clk) begin
    if (reset == 1'b1)
    begin
        mOutPtr <= ~{ADDR_WIDTH+1{1'b0}};
        internal_empty_n <= 1'b0;
        internal_full_n <= 1'b1;
    end
    else begin
        if (((if_read & if_read_ce) == 1 & internal_empty_n == 1) && 
            ((if_write & if_write_ce) == 0 | internal_full_n == 0))
        begin
            mOutPtr <= mOutPtr - 2'd1;
            if (mOutPtr == 2'd0)
                internal_empty_n <= 1'b0;
            internal_full_n <= 1'b1;
        end 
        else if (((if_read & if_read_ce) == 0 | internal_empty_n == 0) && 
            ((if_write & if_write_ce) == 1 & internal_full_n == 1))
        begin
            mOutPtr <= mOutPtr + 2'd1;
            internal_empty_n <= 1'b1;
            if (mOutPtr == DEPTH - 2'd2)
                internal_full_n <= 1'b0;
        end 
    end
end

assign shiftReg_addr = mOutPtr[ADDR_WIDTH] == 1'b0 ? mOutPtr[ADDR_WIDTH-1:0]:{ADDR_WIDTH{1'b0}};
assign shiftReg_ce = (if_write & if_write_ce) & internal_full_n;

td_fused_top_start_for_tdf9_readFilters62_U0_shiftReg 
U_td_fused_top_start_for_tdf9_readFilters62_U0_ram (
    .clk(clk),
    .data(shiftReg_data),
    .ce(shiftReg_ce),
    .a(shiftReg_addr),
    .q(shiftReg_q)
);

endmodule  

// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf10_15 (
        in_data_address0,
        in_data_ce0,
        in_data_d0,
        in_data_q0,
        in_data_we0,
        in_data_address1,
        in_data_ce1,
        in_data_d1,
        in_data_q1,
        in_data_we1,
        out_data_address0,
        out_data_ce0,
        out_data_d0,
        out_data_q0,
        out_data_we0,
        out_data_address1,
        out_data_ce1,
        out_data_d1,
        out_data_q1,
        out_data_we1,
        l1_filter_data_address0,
        l1_filter_data_ce0,
        l1_filter_data_d0,
        l1_filter_data_q0,
        l1_filter_data_we0,
        l1_filter_data_address1,
        l1_filter_data_ce1,
        l1_filter_data_d1,
        l1_filter_data_q1,
        l1_filter_data_we1,
        l2_filter_data_address0,
        l2_filter_data_ce0,
        l2_filter_data_d0,
        l2_filter_data_q0,
        l2_filter_data_we0,
        l2_filter_data_address1,
        l2_filter_data_ce1,
        l2_filter_data_d1,
        l2_filter_data_q1,
        l2_filter_data_we1,
        l1_adjustments_address0,
        l1_adjustments_ce0,
        l1_adjustments_d0,
        l1_adjustments_q0,
        l1_adjustments_we0,
        l1_adjustments_address1,
        l1_adjustments_ce1,
        l1_adjustments_d1,
        l1_adjustments_q1,
        l1_adjustments_we1,
        l2_adjustments_address0,
        l2_adjustments_ce0,
        l2_adjustments_d0,
        l2_adjustments_q0,
        l2_adjustments_we0,
        l2_adjustments_address1,
        l2_adjustments_ce1,
        l2_adjustments_d1,
        l2_adjustments_q1,
        l2_adjustments_we1,
        ap_clk,
        ap_rst,
        in_data_empty_n,
        in_data_read,
        out_data_full_n,
        out_data_write,
        ap_start,
        ap_done,
        ap_ready,
        ap_idle,
        ap_continue
);


output  [11:0] in_data_address0;
output   in_data_ce0;
output  [63:0] in_data_d0;
input  [63:0] in_data_q0;
output   in_data_we0;
output  [11:0] in_data_address1;
output   in_data_ce1;
output  [63:0] in_data_d1;
input  [63:0] in_data_q1;
output   in_data_we1;
output  [11:0] out_data_address0;
output   out_data_ce0;
output  [63:0] out_data_d0;
input  [63:0] out_data_q0;
output   out_data_we0;
output  [11:0] out_data_address1;
output   out_data_ce1;
output  [63:0] out_data_d1;
input  [63:0] out_data_q1;
output   out_data_we1;
output  [16:0] l1_filter_data_address0;
output   l1_filter_data_ce0;
output  [63:0] l1_filter_data_d0;
input  [63:0] l1_filter_data_q0;
output   l1_filter_data_we0;
output  [16:0] l1_filter_data_address1;
output   l1_filter_data_ce1;
output  [63:0] l1_filter_data_d1;
input  [63:0] l1_filter_data_q1;
output   l1_filter_data_we1;
output  [14:0] l2_filter_data_address0;
output   l2_filter_data_ce0;
output  [15:0] l2_filter_data_d0;
input  [15:0] l2_filter_data_q0;
output   l2_filter_data_we0;
output  [14:0] l2_filter_data_address1;
output   l2_filter_data_ce1;
output  [15:0] l2_filter_data_d1;
input  [15:0] l2_filter_data_q1;
output   l2_filter_data_we1;
output  [8:0] l1_adjustments_address0;
output   l1_adjustments_ce0;
output  [47:0] l1_adjustments_d0;
input  [47:0] l1_adjustments_q0;
output   l1_adjustments_we0;
output  [8:0] l1_adjustments_address1;
output   l1_adjustments_ce1;
output  [47:0] l1_adjustments_d1;
input  [47:0] l1_adjustments_q1;
output   l1_adjustments_we1;
output  [5:0] l2_adjustments_address0;
output   l2_adjustments_ce0;
output  [47:0] l2_adjustments_d0;
input  [47:0] l2_adjustments_q0;
output   l2_adjustments_we0;
output  [5:0] l2_adjustments_address1;
output   l2_adjustments_ce1;
output  [47:0] l2_adjustments_d1;
input  [47:0] l2_adjustments_q1;
output   l2_adjustments_we1;
input   ap_clk;
input   ap_rst;
input   in_data_empty_n;
output   in_data_read;
input   out_data_full_n;
output   out_data_write;
input   ap_start;
output   ap_done;
output   ap_ready;
output   ap_idle;
input   ap_continue;

reg ap_done;
reg ap_ready;
reg ap_idle;

wire   [11:0] dataflow_in_loop_TOP_LOOP38364_U0_in_data_address0;
wire    dataflow_in_loop_TOP_LOOP38364_U0_in_data_ce0;
wire   [63:0] dataflow_in_loop_TOP_LOOP38364_U0_in_data_d0;
wire    dataflow_in_loop_TOP_LOOP38364_U0_in_data_we0;
wire   [11:0] dataflow_in_loop_TOP_LOOP38364_U0_in_data_address1;
wire    dataflow_in_loop_TOP_LOOP38364_U0_in_data_ce1;
wire   [63:0] dataflow_in_loop_TOP_LOOP38364_U0_in_data_d1;
wire    dataflow_in_loop_TOP_LOOP38364_U0_in_data_we1;
wire   [16:0] dataflow_in_loop_TOP_LOOP38364_U0_l1_filter_data_address0;
wire    dataflow_in_loop_TOP_LOOP38364_U0_l1_filter_data_ce0;
wire   [63:0] dataflow_in_loop_TOP_LOOP38364_U0_l1_filter_data_d0;
wire    dataflow_in_loop_TOP_LOOP38364_U0_l1_filter_data_we0;
wire   [16:0] dataflow_in_loop_TOP_LOOP38364_U0_l1_filter_data_address1;
wire    dataflow_in_loop_TOP_LOOP38364_U0_l1_filter_data_ce1;
wire   [63:0] dataflow_in_loop_TOP_LOOP38364_U0_l1_filter_data_d1;
wire    dataflow_in_loop_TOP_LOOP38364_U0_l1_filter_data_we1;
wire   [8:0] dataflow_in_loop_TOP_LOOP38364_U0_l1_adjustments_address0;
wire    dataflow_in_loop_TOP_LOOP38364_U0_l1_adjustments_ce0;
wire   [47:0] dataflow_in_loop_TOP_LOOP38364_U0_l1_adjustments_d0;
wire    dataflow_in_loop_TOP_LOOP38364_U0_l1_adjustments_we0;
wire   [8:0] dataflow_in_loop_TOP_LOOP38364_U0_l1_adjustments_address1;
wire    dataflow_in_loop_TOP_LOOP38364_U0_l1_adjustments_ce1;
wire   [47:0] dataflow_in_loop_TOP_LOOP38364_U0_l1_adjustments_d1;
wire    dataflow_in_loop_TOP_LOOP38364_U0_l1_adjustments_we1;
wire   [14:0] dataflow_in_loop_TOP_LOOP38364_U0_l2_filter_data_address0;
wire    dataflow_in_loop_TOP_LOOP38364_U0_l2_filter_data_ce0;
wire   [15:0] dataflow_in_loop_TOP_LOOP38364_U0_l2_filter_data_d0;
wire    dataflow_in_loop_TOP_LOOP38364_U0_l2_filter_data_we0;
wire   [14:0] dataflow_in_loop_TOP_LOOP38364_U0_l2_filter_data_address1;
wire    dataflow_in_loop_TOP_LOOP38364_U0_l2_filter_data_ce1;
wire   [15:0] dataflow_in_loop_TOP_LOOP38364_U0_l2_filter_data_d1;
wire    dataflow_in_loop_TOP_LOOP38364_U0_l2_filter_data_we1;
wire   [11:0] dataflow_in_loop_TOP_LOOP38364_U0_out_data_address0;
wire    dataflow_in_loop_TOP_LOOP38364_U0_out_data_ce0;
wire   [63:0] dataflow_in_loop_TOP_LOOP38364_U0_out_data_d0;
wire    dataflow_in_loop_TOP_LOOP38364_U0_out_data_we0;
wire   [11:0] dataflow_in_loop_TOP_LOOP38364_U0_out_data_address1;
wire    dataflow_in_loop_TOP_LOOP38364_U0_out_data_ce1;
wire   [63:0] dataflow_in_loop_TOP_LOOP38364_U0_out_data_d1;
wire    dataflow_in_loop_TOP_LOOP38364_U0_out_data_we1;
wire   [5:0] dataflow_in_loop_TOP_LOOP38364_U0_l2_adjustments_address0;
wire    dataflow_in_loop_TOP_LOOP38364_U0_l2_adjustments_ce0;
wire   [47:0] dataflow_in_loop_TOP_LOOP38364_U0_l2_adjustments_d0;
wire    dataflow_in_loop_TOP_LOOP38364_U0_l2_adjustments_we0;
wire   [5:0] dataflow_in_loop_TOP_LOOP38364_U0_l2_adjustments_address1;
wire    dataflow_in_loop_TOP_LOOP38364_U0_l2_adjustments_ce1;
wire   [47:0] dataflow_in_loop_TOP_LOOP38364_U0_l2_adjustments_d1;
wire    dataflow_in_loop_TOP_LOOP38364_U0_l2_adjustments_we1;
wire    dataflow_in_loop_TOP_LOOP38364_U0_ap_start;
wire    dataflow_in_loop_TOP_LOOP38364_U0_in_data_read;
wire    dataflow_in_loop_TOP_LOOP38364_U0_out_data_write;
wire    dataflow_in_loop_TOP_LOOP38364_U0_ap_done;
wire    dataflow_in_loop_TOP_LOOP38364_U0_ap_ready;
wire    dataflow_in_loop_TOP_LOOP38364_U0_ap_idle;
reg    dataflow_in_loop_TOP_LOOP38364_U0_ap_continue;
wire    dataflow_in_loop_TOP_LOOP38364_U0_in_data_full_n;
wire    dataflow_in_loop_TOP_LOOP38364_U0_in_data_write;
wire    ap_sync_continue;
wire    ap_sync_done;
wire    ap_sync_ready;
reg   [16:0] loop_dataflow_input_count;
reg   [16:0] loop_dataflow_output_count;
wire   [16:0] bound_minus_1;
wire    dataflow_in_loop_TOP_LOOP38364_U0_start_full_n;
wire    dataflow_in_loop_TOP_LOOP38364_U0_start_write;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 loop_dataflow_input_count = 17'd0;
#0 loop_dataflow_output_count = 17'd0;
end

td_fused_top_dataflow_in_loop_TOP_LOOP38364 dataflow_in_loop_TOP_LOOP38364_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .in_data_address0(dataflow_in_loop_TOP_LOOP38364_U0_in_data_address0),
    .in_data_ce0(dataflow_in_loop_TOP_LOOP38364_U0_in_data_ce0),
    .in_data_d0(dataflow_in_loop_TOP_LOOP38364_U0_in_data_d0),
    .in_data_q0(in_data_q0),
    .in_data_we0(dataflow_in_loop_TOP_LOOP38364_U0_in_data_we0),
    .in_data_address1(dataflow_in_loop_TOP_LOOP38364_U0_in_data_address1),
    .in_data_ce1(dataflow_in_loop_TOP_LOOP38364_U0_in_data_ce1),
    .in_data_d1(dataflow_in_loop_TOP_LOOP38364_U0_in_data_d1),
    .in_data_q1(64'd0),
    .in_data_we1(dataflow_in_loop_TOP_LOOP38364_U0_in_data_we1),
    .l1_filter_data_address0(dataflow_in_loop_TOP_LOOP38364_U0_l1_filter_data_address0),
    .l1_filter_data_ce0(dataflow_in_loop_TOP_LOOP38364_U0_l1_filter_data_ce0),
    .l1_filter_data_d0(dataflow_in_loop_TOP_LOOP38364_U0_l1_filter_data_d0),
    .l1_filter_data_q0(l1_filter_data_q0),
    .l1_filter_data_we0(dataflow_in_loop_TOP_LOOP38364_U0_l1_filter_data_we0),
    .l1_filter_data_address1(dataflow_in_loop_TOP_LOOP38364_U0_l1_filter_data_address1),
    .l1_filter_data_ce1(dataflow_in_loop_TOP_LOOP38364_U0_l1_filter_data_ce1),
    .l1_filter_data_d1(dataflow_in_loop_TOP_LOOP38364_U0_l1_filter_data_d1),
    .l1_filter_data_q1(64'd0),
    .l1_filter_data_we1(dataflow_in_loop_TOP_LOOP38364_U0_l1_filter_data_we1),
    .l1_adjustments_address0(dataflow_in_loop_TOP_LOOP38364_U0_l1_adjustments_address0),
    .l1_adjustments_ce0(dataflow_in_loop_TOP_LOOP38364_U0_l1_adjustments_ce0),
    .l1_adjustments_d0(dataflow_in_loop_TOP_LOOP38364_U0_l1_adjustments_d0),
    .l1_adjustments_q0(l1_adjustments_q0),
    .l1_adjustments_we0(dataflow_in_loop_TOP_LOOP38364_U0_l1_adjustments_we0),
    .l1_adjustments_address1(dataflow_in_loop_TOP_LOOP38364_U0_l1_adjustments_address1),
    .l1_adjustments_ce1(dataflow_in_loop_TOP_LOOP38364_U0_l1_adjustments_ce1),
    .l1_adjustments_d1(dataflow_in_loop_TOP_LOOP38364_U0_l1_adjustments_d1),
    .l1_adjustments_q1(48'd0),
    .l1_adjustments_we1(dataflow_in_loop_TOP_LOOP38364_U0_l1_adjustments_we1),
    .l2_filter_data_address0(dataflow_in_loop_TOP_LOOP38364_U0_l2_filter_data_address0),
    .l2_filter_data_ce0(dataflow_in_loop_TOP_LOOP38364_U0_l2_filter_data_ce0),
    .l2_filter_data_d0(dataflow_in_loop_TOP_LOOP38364_U0_l2_filter_data_d0),
    .l2_filter_data_q0(l2_filter_data_q0),
    .l2_filter_data_we0(dataflow_in_loop_TOP_LOOP38364_U0_l2_filter_data_we0),
    .l2_filter_data_address1(dataflow_in_loop_TOP_LOOP38364_U0_l2_filter_data_address1),
    .l2_filter_data_ce1(dataflow_in_loop_TOP_LOOP38364_U0_l2_filter_data_ce1),
    .l2_filter_data_d1(dataflow_in_loop_TOP_LOOP38364_U0_l2_filter_data_d1),
    .l2_filter_data_q1(16'd0),
    .l2_filter_data_we1(dataflow_in_loop_TOP_LOOP38364_U0_l2_filter_data_we1),
    .out_data_address0(dataflow_in_loop_TOP_LOOP38364_U0_out_data_address0),
    .out_data_ce0(dataflow_in_loop_TOP_LOOP38364_U0_out_data_ce0),
    .out_data_d0(dataflow_in_loop_TOP_LOOP38364_U0_out_data_d0),
    .out_data_q0(64'd0),
    .out_data_we0(dataflow_in_loop_TOP_LOOP38364_U0_out_data_we0),
    .out_data_address1(dataflow_in_loop_TOP_LOOP38364_U0_out_data_address1),
    .out_data_ce1(dataflow_in_loop_TOP_LOOP38364_U0_out_data_ce1),
    .out_data_d1(dataflow_in_loop_TOP_LOOP38364_U0_out_data_d1),
    .out_data_q1(64'd0),
    .out_data_we1(dataflow_in_loop_TOP_LOOP38364_U0_out_data_we1),
    .l2_adjustments_address0(dataflow_in_loop_TOP_LOOP38364_U0_l2_adjustments_address0),
    .l2_adjustments_ce0(dataflow_in_loop_TOP_LOOP38364_U0_l2_adjustments_ce0),
    .l2_adjustments_d0(dataflow_in_loop_TOP_LOOP38364_U0_l2_adjustments_d0),
    .l2_adjustments_q0(l2_adjustments_q0),
    .l2_adjustments_we0(dataflow_in_loop_TOP_LOOP38364_U0_l2_adjustments_we0),
    .l2_adjustments_address1(dataflow_in_loop_TOP_LOOP38364_U0_l2_adjustments_address1),
    .l2_adjustments_ce1(dataflow_in_loop_TOP_LOOP38364_U0_l2_adjustments_ce1),
    .l2_adjustments_d1(dataflow_in_loop_TOP_LOOP38364_U0_l2_adjustments_d1),
    .l2_adjustments_q1(48'd0),
    .l2_adjustments_we1(dataflow_in_loop_TOP_LOOP38364_U0_l2_adjustments_we1),
    .ap_start(dataflow_in_loop_TOP_LOOP38364_U0_ap_start),
    .in_data_empty_n(1'b0),
    .in_data_read(dataflow_in_loop_TOP_LOOP38364_U0_in_data_read),
    .out_data_full_n(out_data_full_n),
    .out_data_write(dataflow_in_loop_TOP_LOOP38364_U0_out_data_write),
    .ap_done(dataflow_in_loop_TOP_LOOP38364_U0_ap_done),
    .ap_ready(dataflow_in_loop_TOP_LOOP38364_U0_ap_ready),
    .ap_idle(dataflow_in_loop_TOP_LOOP38364_U0_ap_idle),
    .ap_continue(dataflow_in_loop_TOP_LOOP38364_U0_ap_continue)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        loop_dataflow_input_count <= 17'd0;
    end else begin
        if ((~(loop_dataflow_input_count == bound_minus_1) & (ap_start == 1'b1) & (dataflow_in_loop_TOP_LOOP38364_U0_ap_ready == 1'b1))) begin
            loop_dataflow_input_count <= (loop_dataflow_input_count + 17'd1);
        end else if (((loop_dataflow_input_count == bound_minus_1) & (ap_start == 1'b1) & (dataflow_in_loop_TOP_LOOP38364_U0_ap_ready == 1'b1))) begin
            loop_dataflow_input_count <= 17'd0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        loop_dataflow_output_count <= 17'd0;
    end else begin
        if ((~(loop_dataflow_output_count == bound_minus_1) & (dataflow_in_loop_TOP_LOOP38364_U0_ap_continue == 1'b1) & (dataflow_in_loop_TOP_LOOP38364_U0_ap_done == 1'b1))) begin
            loop_dataflow_output_count <= (loop_dataflow_output_count + 17'd1);
        end else if (((loop_dataflow_output_count == bound_minus_1) & (dataflow_in_loop_TOP_LOOP38364_U0_ap_continue == 1'b1) & (dataflow_in_loop_TOP_LOOP38364_U0_ap_done == 1'b1))) begin
            loop_dataflow_output_count <= 17'd0;
        end
    end
end

always @ (*) begin
    if (((loop_dataflow_output_count == bound_minus_1) & (dataflow_in_loop_TOP_LOOP38364_U0_ap_done == 1'b1))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = 1'b0;
    end
end

always @ (*) begin
    if (((loop_dataflow_output_count == 17'd0) & (ap_start == 1'b0) & (dataflow_in_loop_TOP_LOOP38364_U0_ap_idle == 1'b1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((loop_dataflow_input_count == bound_minus_1) & (ap_start == 1'b1) & (dataflow_in_loop_TOP_LOOP38364_U0_ap_ready == 1'b1))) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((~(loop_dataflow_output_count == bound_minus_1) | (ap_continue == 1'b1))) begin
        dataflow_in_loop_TOP_LOOP38364_U0_ap_continue = 1'b1;
    end else begin
        dataflow_in_loop_TOP_LOOP38364_U0_ap_continue = 1'b0;
    end
end

assign ap_sync_continue = ap_continue;

assign ap_sync_done = dataflow_in_loop_TOP_LOOP38364_U0_ap_done;

assign ap_sync_ready = dataflow_in_loop_TOP_LOOP38364_U0_ap_ready;

assign bound_minus_1 = (17'd100352 - 17'd1);

assign dataflow_in_loop_TOP_LOOP38364_U0_ap_start = ap_start;

assign dataflow_in_loop_TOP_LOOP38364_U0_in_data_full_n = in_data_empty_n;

assign dataflow_in_loop_TOP_LOOP38364_U0_in_data_write = 1'b0;

assign dataflow_in_loop_TOP_LOOP38364_U0_start_full_n = 1'b1;

assign dataflow_in_loop_TOP_LOOP38364_U0_start_write = 1'b0;

assign in_data_address0 = dataflow_in_loop_TOP_LOOP38364_U0_in_data_address0;

assign in_data_address1 = 12'd0;

assign in_data_ce0 = dataflow_in_loop_TOP_LOOP38364_U0_in_data_ce0;

assign in_data_ce1 = 1'b0;

assign in_data_d0 = 64'd0;

assign in_data_d1 = 64'd0;

assign in_data_read = dataflow_in_loop_TOP_LOOP38364_U0_in_data_write;

assign in_data_we0 = 1'b0;

assign in_data_we1 = 1'b0;

assign l1_adjustments_address0 = dataflow_in_loop_TOP_LOOP38364_U0_l1_adjustments_address0;

assign l1_adjustments_address1 = 9'd0;

assign l1_adjustments_ce0 = dataflow_in_loop_TOP_LOOP38364_U0_l1_adjustments_ce0;

assign l1_adjustments_ce1 = 1'b0;

assign l1_adjustments_d0 = 48'd0;

assign l1_adjustments_d1 = 48'd0;

assign l1_adjustments_we0 = 1'b0;

assign l1_adjustments_we1 = 1'b0;

assign l1_filter_data_address0 = dataflow_in_loop_TOP_LOOP38364_U0_l1_filter_data_address0;

assign l1_filter_data_address1 = 17'd0;

assign l1_filter_data_ce0 = dataflow_in_loop_TOP_LOOP38364_U0_l1_filter_data_ce0;

assign l1_filter_data_ce1 = 1'b0;

assign l1_filter_data_d0 = 64'd0;

assign l1_filter_data_d1 = 64'd0;

assign l1_filter_data_we0 = 1'b0;

assign l1_filter_data_we1 = 1'b0;

assign l2_adjustments_address0 = dataflow_in_loop_TOP_LOOP38364_U0_l2_adjustments_address0;

assign l2_adjustments_address1 = 6'd0;

assign l2_adjustments_ce0 = dataflow_in_loop_TOP_LOOP38364_U0_l2_adjustments_ce0;

assign l2_adjustments_ce1 = 1'b0;

assign l2_adjustments_d0 = 48'd0;

assign l2_adjustments_d1 = 48'd0;

assign l2_adjustments_we0 = 1'b0;

assign l2_adjustments_we1 = 1'b0;

assign l2_filter_data_address0 = dataflow_in_loop_TOP_LOOP38364_U0_l2_filter_data_address0;

assign l2_filter_data_address1 = 15'd0;

assign l2_filter_data_ce0 = dataflow_in_loop_TOP_LOOP38364_U0_l2_filter_data_ce0;

assign l2_filter_data_ce1 = 1'b0;

assign l2_filter_data_d0 = 16'd0;

assign l2_filter_data_d1 = 16'd0;

assign l2_filter_data_we0 = 1'b0;

assign l2_filter_data_we1 = 1'b0;

assign out_data_address0 = 12'd0;

assign out_data_address1 = dataflow_in_loop_TOP_LOOP38364_U0_out_data_address1;

assign out_data_ce0 = 1'b0;

assign out_data_ce1 = dataflow_in_loop_TOP_LOOP38364_U0_out_data_ce1;

assign out_data_d0 = 64'd0;

assign out_data_d1 = dataflow_in_loop_TOP_LOOP38364_U0_out_data_d1;

assign out_data_we0 = 1'b0;

assign out_data_we1 = dataflow_in_loop_TOP_LOOP38364_U0_out_data_we1;

assign out_data_write = dataflow_in_loop_TOP_LOOP38364_U0_out_data_write;

endmodule //td_fused_top_tdf10_15
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf10_accum_1 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        accum_in_0_address0,
        accum_in_0_ce0,
        accum_in_0_q0,
        accum_in_0_address1,
        accum_in_0_ce1,
        accum_in_0_q1,
        accum_out_address0,
        accum_out_ce0,
        accum_out_we0,
        accum_out_d0,
        accum_out_address1,
        accum_out_ce1,
        accum_out_we1,
        accum_out_d1
);

parameter    ap_ST_fsm_state1 = 8'd1;
parameter    ap_ST_fsm_pp0_stage0 = 8'd2;
parameter    ap_ST_fsm_pp0_stage1 = 8'd4;
parameter    ap_ST_fsm_pp0_stage2 = 8'd8;
parameter    ap_ST_fsm_pp0_stage3 = 8'd16;
parameter    ap_ST_fsm_state12 = 8'd32;
parameter    ap_ST_fsm_state13 = 8'd64;
parameter    ap_ST_fsm_state14 = 8'd128;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [9:0] accum_in_0_address0;
output   accum_in_0_ce0;
input  [15:0] accum_in_0_q0;
output  [9:0] accum_in_0_address1;
output   accum_in_0_ce1;
input  [15:0] accum_in_0_q1;
output  [2:0] accum_out_address0;
output   accum_out_ce0;
output   accum_out_we0;
output  [15:0] accum_out_d0;
output  [2:0] accum_out_address1;
output   accum_out_ce1;
output   accum_out_we1;
output  [15:0] accum_out_d1;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg[9:0] accum_in_0_address0;
reg accum_in_0_ce0;
reg[9:0] accum_in_0_address1;
reg accum_in_0_ce1;
reg accum_out_ce0;
reg accum_out_we0;
reg accum_out_ce1;
reg accum_out_we1;

reg    ap_done_reg;
  reg   [7:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg   [9:0] x_reg_168;
reg   [15:0] psum_7_08_reg_180;
reg   [15:0] psum_6_07_reg_192;
reg   [15:0] psum_5_06_reg_204;
reg   [15:0] psum_4_05_reg_216;
reg   [15:0] psum_3_04_reg_228;
reg   [15:0] psum_2_03_reg_240;
reg   [15:0] psum_1_02_reg_252;
reg   [15:0] psum_0_01_reg_264;
wire   [0:0] icmp_ln132_fu_321_p2;
reg   [0:0] icmp_ln132_reg_492;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state6_pp0_stage0_iter1;
wire    ap_block_state10_pp0_stage0_iter2;
wire    ap_block_pp0_stage0_11001;
reg   [0:0] icmp_ln132_reg_492_pp0_iter1_reg;
reg   [0:0] icmp_ln132_reg_492_pp0_iter2_reg;
reg   [15:0] accum_in_0_load_reg_506;
wire    ap_CS_fsm_pp0_stage1;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_state3_pp0_stage1_iter0;
wire    ap_block_state7_pp0_stage1_iter1;
wire    ap_block_state11_pp0_stage1_iter2;
wire    ap_block_pp0_stage1_11001;
reg   [15:0] accum_in_0_load_72_reg_511;
reg   [15:0] accum_in_0_load_73_reg_526;
wire    ap_CS_fsm_pp0_stage2;
wire    ap_block_state4_pp0_stage2_iter0;
wire    ap_block_state8_pp0_stage2_iter1;
wire    ap_block_pp0_stage2_11001;
reg   [15:0] accum_in_0_load_74_reg_531;
wire   [9:0] add_ln132_fu_387_p2;
reg   [9:0] add_ln132_reg_546;
wire    ap_CS_fsm_pp0_stage3;
wire    ap_block_state5_pp0_stage3_iter0;
wire    ap_block_state9_pp0_stage3_iter1;
wire    ap_block_pp0_stage3_11001;
reg   [15:0] accum_in_0_load_75_reg_551;
reg   [15:0] accum_in_0_load_76_reg_556;
reg   [15:0] accum_in_0_load_77_reg_571;
reg    ap_enable_reg_pp0_iter1;
reg   [15:0] accum_in_0_load_78_reg_576;
wire   [15:0] grp_fu_305_p2;
wire   [15:0] grp_fu_310_p2;
reg    ap_enable_reg_pp0_iter2;
wire   [3:0] add_ln140_fu_432_p2;
wire    ap_CS_fsm_state13;
wire   [0:0] tmp_fu_415_p3;
reg    ap_block_state1;
wire    ap_block_pp0_stage2_subdone;
reg    ap_condition_pp0_exit_iter0_state4;
wire    ap_block_pp0_stage3_subdone;
wire    ap_block_pp0_stage1_subdone;
reg   [9:0] ap_phi_mux_x_phi_fu_172_p4;
wire    ap_block_pp0_stage0;
wire   [15:0] ap_phi_mux_psum_7_08_phi_fu_184_p4;
wire    ap_block_pp0_stage1;
wire   [15:0] ap_phi_mux_psum_6_07_phi_fu_196_p4;
wire   [15:0] ap_phi_mux_psum_5_06_phi_fu_208_p4;
wire   [15:0] ap_phi_mux_psum_4_05_phi_fu_220_p4;
wire   [15:0] ap_phi_mux_psum_3_04_phi_fu_232_p4;
wire    ap_block_pp0_stage3;
wire   [15:0] ap_phi_mux_psum_2_03_phi_fu_244_p4;
wire    ap_block_pp0_stage2;
reg   [3:0] q_reg_276;
wire    ap_CS_fsm_state12;
reg   [15:0] ap_phi_mux_phi_ln152_phi_fu_290_p8;
wire   [2:0] trunc_ln140_fu_428_p1;
wire   [63:0] zext_ln132_fu_327_p1;
wire   [63:0] zext_ln136_fu_338_p1;
wire   [63:0] zext_ln136_19_fu_349_p1;
wire   [63:0] zext_ln136_20_fu_360_p1;
wire   [63:0] zext_ln136_21_fu_371_p1;
wire   [63:0] zext_ln136_22_fu_382_p1;
wire   [63:0] zext_ln136_23_fu_399_p1;
wire   [63:0] zext_ln136_24_fu_410_p1;
wire   [63:0] zext_ln140_fu_423_p1;
wire   [63:0] zext_ln140_4_fu_444_p1;
reg   [15:0] grp_fu_305_p0;
reg   [15:0] grp_fu_305_p1;
reg   [15:0] grp_fu_310_p0;
reg   [15:0] grp_fu_310_p1;
wire   [9:0] or_ln136_fu_332_p2;
wire   [9:0] or_ln136_19_fu_343_p2;
wire   [9:0] or_ln136_20_fu_354_p2;
wire   [9:0] or_ln136_21_fu_365_p2;
wire   [9:0] or_ln136_22_fu_376_p2;
wire   [9:0] or_ln136_23_fu_393_p2;
wire   [9:0] or_ln136_24_fu_404_p2;
wire   [2:0] or_ln140_fu_438_p2;
wire   [0:0] icmp_ln152_fu_449_p2;
wire   [0:0] icmp_ln152_7_fu_463_p2;
wire   [15:0] select_ln152_fu_455_p3;
wire   [0:0] icmp_ln152_8_fu_477_p2;
wire   [15:0] select_ln152_7_fu_469_p3;
wire    ap_CS_fsm_state14;
reg   [7:0] ap_NS_fsm;
wire    ap_block_pp0_stage0_subdone;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
reg    ap_condition_514;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 8'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
end

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U622(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(grp_fu_305_p0),
    .din1(grp_fu_305_p1),
    .dout(grp_fu_305_p2)
);

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U623(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(grp_fu_310_p0),
    .din1(grp_fu_310_p1),
    .dout(grp_fu_310_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state14)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage2_subdone) & (1'b1 == ap_condition_pp0_exit_iter0_state4) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage3_subdone) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b0)) | ((1'b0 == ap_block_pp0_stage3_subdone) & (1'b1 == ap_CS_fsm_pp0_stage3)))) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end else if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter2 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state12)) begin
        q_reg_276 <= 4'd0;
    end else if (((tmp_fu_415_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state13))) begin
        q_reg_276 <= add_ln140_fu_432_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln132_reg_492 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        x_reg_168 <= add_ln132_reg_546;
    end else if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        x_reg_168 <= 10'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage1_11001) & (icmp_ln132_reg_492 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
        accum_in_0_load_72_reg_511 <= accum_in_0_q0;
        accum_in_0_load_reg_506 <= accum_in_0_q1;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2_11001) & (icmp_ln132_reg_492 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
        accum_in_0_load_73_reg_526 <= accum_in_0_q1;
        accum_in_0_load_74_reg_531 <= accum_in_0_q0;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage3_11001) & (icmp_ln132_reg_492 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
        accum_in_0_load_75_reg_551 <= accum_in_0_q1;
        accum_in_0_load_76_reg_556 <= accum_in_0_q0;
        add_ln132_reg_546 <= add_ln132_fu_387_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln132_reg_492 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        accum_in_0_load_77_reg_571 <= accum_in_0_q1;
        accum_in_0_load_78_reg_576 <= accum_in_0_q0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln132_reg_492 <= icmp_ln132_fu_321_p2;
        icmp_ln132_reg_492_pp0_iter1_reg <= icmp_ln132_reg_492;
        icmp_ln132_reg_492_pp0_iter2_reg <= icmp_ln132_reg_492_pp0_iter1_reg;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln132_reg_492_pp0_iter1_reg == 1'd1) & (1'b0 == ap_block_pp0_stage2_11001) & (1'b1 == ap_CS_fsm_pp0_stage2) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        psum_0_01_reg_264 <= grp_fu_305_p2;
        psum_1_02_reg_252 <= grp_fu_310_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln132_reg_492_pp0_iter1_reg == 1'd1) & (1'b0 == ap_block_pp0_stage3_11001) & (1'b1 == ap_CS_fsm_pp0_stage3) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        psum_2_03_reg_240 <= grp_fu_305_p2;
        psum_3_04_reg_228 <= grp_fu_310_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln132_reg_492_pp0_iter1_reg == 1'd1) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        psum_4_05_reg_216 <= grp_fu_305_p2;
        psum_5_06_reg_204 <= grp_fu_310_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln132_reg_492_pp0_iter2_reg == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        psum_6_07_reg_192 <= grp_fu_305_p2;
        psum_7_08_reg_180 <= grp_fu_310_p2;
    end
end

always @ (*) begin
    if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
        if (((1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            accum_in_0_address0 = zext_ln136_24_fu_410_p1;
        end else if (((1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            accum_in_0_address0 = zext_ln136_22_fu_382_p1;
        end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            accum_in_0_address0 = zext_ln136_20_fu_360_p1;
        end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            accum_in_0_address0 = zext_ln136_fu_338_p1;
        end else begin
            accum_in_0_address0 = 'bx;
        end
    end else begin
        accum_in_0_address0 = 'bx;
    end
end

always @ (*) begin
    if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
        if (((1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            accum_in_0_address1 = zext_ln136_23_fu_399_p1;
        end else if (((1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            accum_in_0_address1 = zext_ln136_21_fu_371_p1;
        end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            accum_in_0_address1 = zext_ln136_19_fu_349_p1;
        end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            accum_in_0_address1 = zext_ln132_fu_327_p1;
        end else begin
            accum_in_0_address1 = 'bx;
        end
    end else begin
        accum_in_0_address1 = 'bx;
    end
end

always @ (*) begin
    if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage3_11001) & (1'b1 == ap_CS_fsm_pp0_stage3)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2_11001) & (1'b1 == ap_CS_fsm_pp0_stage2)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1)))) begin
        accum_in_0_ce0 = 1'b1;
    end else begin
        accum_in_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage3_11001) & (1'b1 == ap_CS_fsm_pp0_stage3)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2_11001) & (1'b1 == ap_CS_fsm_pp0_stage2)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1)))) begin
        accum_in_0_ce1 = 1'b1;
    end else begin
        accum_in_0_ce1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state13)) begin
        accum_out_ce0 = 1'b1;
    end else begin
        accum_out_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state13)) begin
        accum_out_ce1 = 1'b1;
    end else begin
        accum_out_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((tmp_fu_415_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state13))) begin
        accum_out_we0 = 1'b1;
    end else begin
        accum_out_we0 = 1'b0;
    end
end

always @ (*) begin
    if (((tmp_fu_415_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state13))) begin
        accum_out_we1 = 1'b1;
    end else begin
        accum_out_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((icmp_ln132_reg_492 == 1'd0)) begin
        ap_condition_pp0_exit_iter0_state4 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state4 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state14)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((tmp_fu_415_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state13))) begin
        if ((trunc_ln140_fu_428_p1 == 3'd0)) begin
            ap_phi_mux_phi_ln152_phi_fu_290_p8 = psum_0_01_reg_264;
        end else if ((1'b1 == ap_condition_514)) begin
            ap_phi_mux_phi_ln152_phi_fu_290_p8 = psum_6_07_reg_192;
        end else if ((trunc_ln140_fu_428_p1 == 3'd4)) begin
            ap_phi_mux_phi_ln152_phi_fu_290_p8 = psum_4_05_reg_216;
        end else if ((trunc_ln140_fu_428_p1 == 3'd2)) begin
            ap_phi_mux_phi_ln152_phi_fu_290_p8 = psum_2_03_reg_240;
        end else begin
            ap_phi_mux_phi_ln152_phi_fu_290_p8 = 'bx;
        end
    end else begin
        ap_phi_mux_phi_ln152_phi_fu_290_p8 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0) & (icmp_ln132_reg_492 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_x_phi_fu_172_p4 = add_ln132_reg_546;
    end else begin
        ap_phi_mux_x_phi_fu_172_p4 = x_reg_168;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state14)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_305_p0 = ap_phi_mux_psum_6_07_phi_fu_196_p4;
    end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_305_p0 = ap_phi_mux_psum_4_05_phi_fu_220_p4;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
        grp_fu_305_p0 = ap_phi_mux_psum_2_03_phi_fu_244_p4;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
        grp_fu_305_p0 = grp_fu_305_p2;
    end else begin
        grp_fu_305_p0 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_305_p1 = accum_in_0_load_77_reg_571;
    end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_305_p1 = accum_in_0_load_75_reg_551;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
        grp_fu_305_p1 = accum_in_0_load_73_reg_526;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
        grp_fu_305_p1 = accum_in_0_load_reg_506;
    end else begin
        grp_fu_305_p1 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_310_p0 = ap_phi_mux_psum_7_08_phi_fu_184_p4;
    end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_310_p0 = ap_phi_mux_psum_5_06_phi_fu_208_p4;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
        grp_fu_310_p0 = ap_phi_mux_psum_3_04_phi_fu_232_p4;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
        grp_fu_310_p0 = grp_fu_310_p2;
    end else begin
        grp_fu_310_p0 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_310_p1 = accum_in_0_load_78_reg_576;
    end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_310_p1 = accum_in_0_load_76_reg_556;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
        grp_fu_310_p1 = accum_in_0_load_74_reg_531;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
        grp_fu_310_p1 = accum_in_0_load_72_reg_511;
    end else begin
        grp_fu_310_p1 = 'bx;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_pp0_stage1 : begin
            if ((~((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter2 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0)) & (1'b0 == ap_block_pp0_stage1_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage2;
            end else if (((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter2 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
                ap_NS_fsm = ap_ST_fsm_state12;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end
        end
        ap_ST_fsm_pp0_stage2 : begin
            if ((~((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2_subdone) & (icmp_ln132_reg_492 == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b0)) & (1'b0 == ap_block_pp0_stage2_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage3;
            end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2_subdone) & (icmp_ln132_reg_492 == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
                ap_NS_fsm = ap_ST_fsm_state12;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage2;
            end
        end
        ap_ST_fsm_pp0_stage3 : begin
            if ((1'b0 == ap_block_pp0_stage3_subdone)) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage3;
            end
        end
        ap_ST_fsm_state12 : begin
            ap_NS_fsm = ap_ST_fsm_state13;
        end
        ap_ST_fsm_state13 : begin
            if (((tmp_fu_415_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state13))) begin
                ap_NS_fsm = ap_ST_fsm_state13;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state14;
            end
        end
        ap_ST_fsm_state14 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign accum_out_address0 = zext_ln140_4_fu_444_p1;

assign accum_out_address1 = zext_ln140_fu_423_p1;

assign accum_out_d0 = ((icmp_ln152_8_fu_477_p2[0:0] == 1'b1) ? psum_5_06_reg_204 : select_ln152_7_fu_469_p3);

assign accum_out_d1 = ap_phi_mux_phi_ln152_phi_fu_290_p8;

assign add_ln132_fu_387_p2 = (x_reg_168 + 10'd8);

assign add_ln140_fu_432_p2 = (q_reg_276 + 4'd2);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_pp0_stage1 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_pp0_stage2 = ap_CS_fsm[32'd3];

assign ap_CS_fsm_pp0_stage3 = ap_CS_fsm[32'd4];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state12 = ap_CS_fsm[32'd5];

assign ap_CS_fsm_state13 = ap_CS_fsm[32'd6];

assign ap_CS_fsm_state14 = ap_CS_fsm[32'd7];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1_subdone = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage2 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage2_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage2_subdone = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage3 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage3_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage3_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((ap_done_reg == 1'b1) | (ap_start == 1'b0));
end

assign ap_block_state10_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state11_pp0_stage1_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage1_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage2_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage3_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage1_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage2_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state9_pp0_stage3_iter1 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_condition_514 = (~(trunc_ln140_fu_428_p1 == 3'd0) & ~(trunc_ln140_fu_428_p1 == 3'd4) & ~(trunc_ln140_fu_428_p1 == 3'd2));
end

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign ap_phi_mux_psum_2_03_phi_fu_244_p4 = grp_fu_305_p2;

assign ap_phi_mux_psum_3_04_phi_fu_232_p4 = grp_fu_310_p2;

assign ap_phi_mux_psum_4_05_phi_fu_220_p4 = grp_fu_305_p2;

assign ap_phi_mux_psum_5_06_phi_fu_208_p4 = grp_fu_310_p2;

assign ap_phi_mux_psum_6_07_phi_fu_196_p4 = grp_fu_305_p2;

assign ap_phi_mux_psum_7_08_phi_fu_184_p4 = grp_fu_310_p2;

assign icmp_ln132_fu_321_p2 = ((ap_phi_mux_x_phi_fu_172_p4 < 10'd576) ? 1'b1 : 1'b0);

assign icmp_ln152_7_fu_463_p2 = ((or_ln140_fu_438_p2 == 3'd3) ? 1'b1 : 1'b0);

assign icmp_ln152_8_fu_477_p2 = ((or_ln140_fu_438_p2 == 3'd5) ? 1'b1 : 1'b0);

assign icmp_ln152_fu_449_p2 = ((or_ln140_fu_438_p2 == 3'd1) ? 1'b1 : 1'b0);

assign or_ln136_19_fu_343_p2 = (x_reg_168 | 10'd2);

assign or_ln136_20_fu_354_p2 = (x_reg_168 | 10'd3);

assign or_ln136_21_fu_365_p2 = (x_reg_168 | 10'd4);

assign or_ln136_22_fu_376_p2 = (x_reg_168 | 10'd5);

assign or_ln136_23_fu_393_p2 = (x_reg_168 | 10'd6);

assign or_ln136_24_fu_404_p2 = (x_reg_168 | 10'd7);

assign or_ln136_fu_332_p2 = (ap_phi_mux_x_phi_fu_172_p4 | 10'd1);

assign or_ln140_fu_438_p2 = (trunc_ln140_fu_428_p1 | 3'd1);

assign select_ln152_7_fu_469_p3 = ((icmp_ln152_7_fu_463_p2[0:0] == 1'b1) ? psum_3_04_reg_228 : select_ln152_fu_455_p3);

assign select_ln152_fu_455_p3 = ((icmp_ln152_fu_449_p2[0:0] == 1'b1) ? psum_1_02_reg_252 : psum_7_08_reg_180);

assign tmp_fu_415_p3 = q_reg_276[32'd3];

assign trunc_ln140_fu_428_p1 = q_reg_276[2:0];

assign zext_ln132_fu_327_p1 = ap_phi_mux_x_phi_fu_172_p4;

assign zext_ln136_19_fu_349_p1 = or_ln136_19_fu_343_p2;

assign zext_ln136_20_fu_360_p1 = or_ln136_20_fu_354_p2;

assign zext_ln136_21_fu_371_p1 = or_ln136_21_fu_365_p2;

assign zext_ln136_22_fu_382_p1 = or_ln136_22_fu_376_p2;

assign zext_ln136_23_fu_399_p1 = or_ln136_23_fu_393_p2;

assign zext_ln136_24_fu_410_p1 = or_ln136_24_fu_404_p2;

assign zext_ln136_fu_338_p1 = or_ln136_fu_332_p2;

assign zext_ln140_4_fu_444_p1 = or_ln140_fu_438_p2;

assign zext_ln140_fu_423_p1 = q_reg_276;

endmodule //td_fused_top_tdf10_accum_1
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf10_accum_2 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        accum_in_24,
        accum_in_24_ap_vld,
        accum_in_address0,
        accum_in_ce0,
        accum_in_q0
);

parameter    ap_ST_fsm_state1 = 7'd1;
parameter    ap_ST_fsm_state2 = 7'd2;
parameter    ap_ST_fsm_state3 = 7'd4;
parameter    ap_ST_fsm_state4 = 7'd8;
parameter    ap_ST_fsm_state5 = 7'd16;
parameter    ap_ST_fsm_state6 = 7'd32;
parameter    ap_ST_fsm_state7 = 7'd64;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [15:0] accum_in_24;
output   accum_in_24_ap_vld;
output  [2:0] accum_in_address0;
output   accum_in_ce0;
input  [15:0] accum_in_q0;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg[15:0] accum_in_24;
reg accum_in_24_ap_vld;
reg accum_in_ce0;

reg    ap_done_reg;
  reg   [6:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
wire   [3:0] add_ln164_fu_74_p2;
reg   [3:0] add_ln164_reg_91;
wire    ap_CS_fsm_state2;
wire   [0:0] icmp_ln164_fu_85_p2;
wire    ap_CS_fsm_state3;
wire   [15:0] grp_fu_68_p2;
wire    ap_CS_fsm_state7;
reg   [3:0] i_1_1_reg_44;
reg    ap_block_state1;
reg   [15:0] sum_01_reg_55;
wire   [63:0] zext_ln164_fu_80_p1;
reg   [15:0] accum_in_24_preg;
reg   [6:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 7'd1;
#0 accum_in_24_preg = 16'd0;
end

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U626(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(sum_01_reg_55),
    .din1(accum_in_q0),
    .dout(grp_fu_68_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        accum_in_24_preg <= 16'd0;
    end else begin
        if (((icmp_ln164_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
            accum_in_24_preg <= sum_01_reg_55;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if (((icmp_ln164_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        i_1_1_reg_44 <= 4'd0;
    end else if ((1'b1 == ap_CS_fsm_state7)) begin
        i_1_1_reg_44 <= add_ln164_reg_91;
    end
end

always @ (posedge ap_clk) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        sum_01_reg_55 <= 16'd0;
    end else if ((1'b1 == ap_CS_fsm_state7)) begin
        sum_01_reg_55 <= grp_fu_68_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        add_ln164_reg_91 <= add_ln164_fu_74_p2;
    end
end

always @ (*) begin
    if (((icmp_ln164_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        accum_in_24 = sum_01_reg_55;
    end else begin
        accum_in_24 = accum_in_24_preg;
    end
end

always @ (*) begin
    if (((icmp_ln164_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        accum_in_24_ap_vld = 1'b1;
    end else begin
        accum_in_24_ap_vld = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        accum_in_ce0 = 1'b1;
    end else begin
        accum_in_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln164_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln164_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_state2 : begin
            if (((icmp_ln164_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end
        end
        ap_ST_fsm_state3 : begin
            ap_NS_fsm = ap_ST_fsm_state4;
        end
        ap_ST_fsm_state4 : begin
            ap_NS_fsm = ap_ST_fsm_state5;
        end
        ap_ST_fsm_state5 : begin
            ap_NS_fsm = ap_ST_fsm_state6;
        end
        ap_ST_fsm_state6 : begin
            ap_NS_fsm = ap_ST_fsm_state7;
        end
        ap_ST_fsm_state7 : begin
            ap_NS_fsm = ap_ST_fsm_state2;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign accum_in_address0 = zext_ln164_fu_80_p1;

assign add_ln164_fu_74_p2 = (i_1_1_reg_44 + 4'd1);

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state7 = ap_CS_fsm[32'd6];

always @ (*) begin
    ap_block_state1 = ((ap_done_reg == 1'b1) | (ap_start == 1'b0));
end

assign icmp_ln164_fu_85_p2 = ((i_1_1_reg_44 == 4'd8) ? 1'b1 : 1'b0);

assign zext_ln164_fu_80_p1 = i_1_1_reg_44;

endmodule //td_fused_top_tdf10_accum_2
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_tdf10_adjustments_ram (addr0, ce0, q0, addr1, ce1, d1, we1,  clk);

parameter DWIDTH = 48;
parameter AWIDTH = 9;
parameter MEM_SIZE = 512;

input[AWIDTH-1:0] addr0;
input ce0;
output wire[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
input clk;

 reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];
wire [AWIDTH-1:0] addr0_t0; 
reg [AWIDTH-1:0] addr0_t1; 
reg [DWIDTH-1:0] q0_t0;
reg [DWIDTH-1:0] q0_t1;
wire [AWIDTH-1:0] addr1_t0; 
reg [AWIDTH-1:0] addr1_t1; 
wire [DWIDTH-1:0] d1_t0; 
wire we1_t0; 
reg [DWIDTH-1:0] d1_t1; 
reg we1_t1; 


assign addr0_t0 = addr0;
assign q0 = q0_t1;
assign addr1_t0 = addr1;
assign d1_t0 = d1;
assign we1_t0 = we1;

always @(posedge clk)  
begin
    if (ce0) 
    begin
        addr0_t1 <= addr0_t0; 
        q0_t1 <= q0_t0;
    end
    if (ce1) 
    begin
        addr1_t1 <= addr1_t0; 
        d1_t1 <= d1_t0;
        we1_t1 <= we1_t0;
    end
end


always @(posedge clk)  
begin 
    if (ce0) begin
        q0_t0 <= ram[addr0_t1];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1_t1) 
            ram[addr1_t1] <= d1_t1; 
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_tdf10_adjustments(
    reset,
    clk,
    address0,
    ce0,
    q0,
    address1,
    ce1,
    we1,
    d1);

parameter DataWidth = 32'd48;
parameter AddressRange = 32'd512;
parameter AddressWidth = 32'd9;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;



td_fused_top_tdf10_adjustments_ram td_fused_top_tdf10_adjustments_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 )
);

endmodule

// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf10_adjust (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        sums_read,
        adjustments_address0,
        adjustments_ce0,
        adjustments_q0,
        indices_23_dout,
        indices_23_empty_n,
        indices_23_read,
        indices_23_out_din,
        indices_23_out_full_n,
        indices_23_out_write,
        ap_return
);

parameter    ap_ST_fsm_state1 = 17'd1;
parameter    ap_ST_fsm_state2 = 17'd2;
parameter    ap_ST_fsm_state3 = 17'd4;
parameter    ap_ST_fsm_state4 = 17'd8;
parameter    ap_ST_fsm_state5 = 17'd16;
parameter    ap_ST_fsm_state6 = 17'd32;
parameter    ap_ST_fsm_state7 = 17'd64;
parameter    ap_ST_fsm_state8 = 17'd128;
parameter    ap_ST_fsm_state9 = 17'd256;
parameter    ap_ST_fsm_state10 = 17'd512;
parameter    ap_ST_fsm_state11 = 17'd1024;
parameter    ap_ST_fsm_state12 = 17'd2048;
parameter    ap_ST_fsm_state13 = 17'd4096;
parameter    ap_ST_fsm_state14 = 17'd8192;
parameter    ap_ST_fsm_state15 = 17'd16384;
parameter    ap_ST_fsm_state16 = 17'd32768;
parameter    ap_ST_fsm_state17 = 17'd65536;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
input  [15:0] sums_read;
output  [8:0] adjustments_address0;
output   adjustments_ce0;
input  [47:0] adjustments_q0;
input  [14:0] indices_23_dout;
input   indices_23_empty_n;
output   indices_23_read;
output  [14:0] indices_23_out_din;
input   indices_23_out_full_n;
output   indices_23_out_write;
output  [15:0] ap_return;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg adjustments_ce0;
reg indices_23_read;
reg indices_23_out_write;

reg    ap_done_reg;
  reg   [16:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    indices_23_blk_n;
reg    indices_23_out_blk_n;
wire    ap_CS_fsm_state4;
reg   [15:0] tmp_110_i_i_reg_183;
reg   [15:0] tmp_111_i_i_reg_188;
wire   [15:0] grp_fu_93_p2;
reg   [15:0] sub_i_i_i_reg_193;
wire    ap_CS_fsm_state8;
wire    ap_CS_fsm_state9;
wire   [15:0] grp_fu_98_p2;
reg   [15:0] mul_i_i_i_reg_203;
wire    ap_CS_fsm_state12;
wire    ap_CS_fsm_state13;
wire   [63:0] zext_ln220_fu_106_p1;
reg    ap_block_state1;
wire    ap_CS_fsm_state2;
wire    ap_CS_fsm_state3;
wire   [15:0] grp_fu_89_p1;
wire   [15:0] grp_fu_93_p1;
wire   [15:0] grp_fu_98_p1;
wire   [8:0] trunc_ln251_fu_102_p1;
wire   [15:0] trunc_ln220_fu_111_p1;
wire   [15:0] grp_fu_89_p2;
wire    ap_CS_fsm_state17;
wire   [15:0] bitcast_ln648_fu_148_p1;
wire   [0:0] tmp_fu_152_p3;
reg   [16:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 17'd1;
end

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U630(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(mul_i_i_i_reg_203),
    .din1(grp_fu_89_p1),
    .dout(grp_fu_89_p2)
);

td_fused_top_hsub_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hsub_16ns_16ns_16_5_full_dsp_1_U631(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(sums_read),
    .din1(grp_fu_93_p1),
    .dout(grp_fu_93_p2)
);

td_fused_top_hmul_16ns_16ns_16_4_max_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hmul_16ns_16ns_16_4_max_dsp_1_U632(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(sub_i_i_i_reg_193),
    .din1(grp_fu_98_p1),
    .dout(grp_fu_98_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state17)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state12)) begin
        mul_i_i_i_reg_203 <= grp_fu_98_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state8)) begin
        sub_i_i_i_reg_193 <= grp_fu_93_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        tmp_110_i_i_reg_183 <= {{adjustments_q0[31:16]}};
        tmp_111_i_i_reg_188 <= {{adjustments_q0[47:32]}};
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state2) | (~((indices_23_out_full_n == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1)))) begin
        adjustments_ce0 = 1'b1;
    end else begin
        adjustments_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state17)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state17)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_23_blk_n = indices_23_empty_n;
    end else begin
        indices_23_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_23_out_blk_n = indices_23_out_full_n;
    end else begin
        indices_23_out_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((indices_23_out_full_n == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_23_out_write = 1'b1;
    end else begin
        indices_23_out_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((indices_23_out_full_n == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_23_read = 1'b1;
    end else begin
        indices_23_read = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((indices_23_out_full_n == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_state2 : begin
            ap_NS_fsm = ap_ST_fsm_state3;
        end
        ap_ST_fsm_state3 : begin
            ap_NS_fsm = ap_ST_fsm_state4;
        end
        ap_ST_fsm_state4 : begin
            ap_NS_fsm = ap_ST_fsm_state5;
        end
        ap_ST_fsm_state5 : begin
            ap_NS_fsm = ap_ST_fsm_state6;
        end
        ap_ST_fsm_state6 : begin
            ap_NS_fsm = ap_ST_fsm_state7;
        end
        ap_ST_fsm_state7 : begin
            ap_NS_fsm = ap_ST_fsm_state8;
        end
        ap_ST_fsm_state8 : begin
            ap_NS_fsm = ap_ST_fsm_state9;
        end
        ap_ST_fsm_state9 : begin
            ap_NS_fsm = ap_ST_fsm_state10;
        end
        ap_ST_fsm_state10 : begin
            ap_NS_fsm = ap_ST_fsm_state11;
        end
        ap_ST_fsm_state11 : begin
            ap_NS_fsm = ap_ST_fsm_state12;
        end
        ap_ST_fsm_state12 : begin
            ap_NS_fsm = ap_ST_fsm_state13;
        end
        ap_ST_fsm_state13 : begin
            ap_NS_fsm = ap_ST_fsm_state14;
        end
        ap_ST_fsm_state14 : begin
            ap_NS_fsm = ap_ST_fsm_state15;
        end
        ap_ST_fsm_state15 : begin
            ap_NS_fsm = ap_ST_fsm_state16;
        end
        ap_ST_fsm_state16 : begin
            ap_NS_fsm = ap_ST_fsm_state17;
        end
        ap_ST_fsm_state17 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign adjustments_address0 = zext_ln220_fu_106_p1;

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state12 = ap_CS_fsm[32'd11];

assign ap_CS_fsm_state13 = ap_CS_fsm[32'd12];

assign ap_CS_fsm_state17 = ap_CS_fsm[32'd16];

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

assign ap_CS_fsm_state8 = ap_CS_fsm[32'd7];

assign ap_CS_fsm_state9 = ap_CS_fsm[32'd8];

always @ (*) begin
    ap_block_state1 = ((indices_23_out_full_n == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0));
end

assign ap_return = ((tmp_fu_152_p3[0:0] == 1'b1) ? 16'd0 : grp_fu_89_p2);

assign bitcast_ln648_fu_148_p1 = grp_fu_89_p2;

assign grp_fu_89_p1 = tmp_111_i_i_reg_188;

assign grp_fu_93_p1 = trunc_ln220_fu_111_p1;

assign grp_fu_98_p1 = tmp_110_i_i_reg_183;

assign indices_23_out_din = indices_23_dout;

assign tmp_fu_152_p3 = bitcast_ln648_fu_148_p1[32'd15];

assign trunc_ln220_fu_111_p1 = adjustments_q0[15:0];

assign trunc_ln251_fu_102_p1 = indices_23_dout[8:0];

assign zext_ln220_fu_106_p1 = trunc_ln251_fu_102_p1;

endmodule //td_fused_top_tdf10_adjust
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf10_dot_product (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        ifmap_vec_address0,
        ifmap_vec_ce0,
        ifmap_vec_q0,
        weight_vecs_0_address0,
        weight_vecs_0_ce0,
        weight_vecs_0_q0,
        products_0_address0,
        products_0_ce0,
        products_0_we0,
        products_0_d0
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state10 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [9:0] ifmap_vec_address0;
output   ifmap_vec_ce0;
input  [15:0] ifmap_vec_q0;
output  [9:0] weight_vecs_0_address0;
output   weight_vecs_0_ce0;
input  [15:0] weight_vecs_0_q0;
output  [9:0] products_0_address0;
output   products_0_ce0;
output   products_0_we0;
output  [15:0] products_0_d0;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg ifmap_vec_ce0;
reg weight_vecs_0_ce0;
reg products_0_ce0;
reg products_0_we0;

reg    ap_done_reg;
  reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg   [9:0] indvar_flatten17_reg_97;
reg   [8:0] indvar_flatten_reg_108;
reg   [1:0] jj_reg_119;
reg   [6:0] ic_reg_131;
reg   [1:0] ii_reg_142;
wire   [9:0] add_ln147_8_fu_157_p2;
wire    ap_CS_fsm_pp0_stage0;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
wire    ap_block_state4_pp0_stage0_iter2;
wire    ap_block_state5_pp0_stage0_iter3;
wire    ap_block_state6_pp0_stage0_iter4;
wire    ap_block_state7_pp0_stage0_iter5;
wire    ap_block_state8_pp0_stage0_iter6;
wire    ap_block_state9_pp0_stage0_iter7;
wire    ap_block_pp0_stage0_11001;
wire   [0:0] icmp_ln147_fu_163_p2;
reg   [0:0] icmp_ln147_reg_408;
reg   [0:0] icmp_ln147_reg_408_pp0_iter1_reg;
reg   [0:0] icmp_ln147_reg_408_pp0_iter2_reg;
reg   [0:0] icmp_ln147_reg_408_pp0_iter3_reg;
reg   [0:0] icmp_ln147_reg_408_pp0_iter4_reg;
reg   [0:0] icmp_ln147_reg_408_pp0_iter5_reg;
reg   [0:0] icmp_ln147_reg_408_pp0_iter6_reg;
wire   [0:0] icmp_ln148_fu_169_p2;
reg   [0:0] icmp_ln148_reg_412;
wire   [0:0] and_ln147_fu_195_p2;
reg   [0:0] and_ln147_reg_419;
wire   [1:0] add_ln148_fu_201_p2;
reg   [1:0] add_ln148_reg_424;
wire   [6:0] select_ln148_fu_213_p3;
reg   [6:0] select_ln148_reg_429;
wire   [1:0] select_ln148_22_fu_221_p3;
reg   [1:0] select_ln148_22_reg_434;
wire   [5:0] trunc_ln150_fu_229_p1;
reg   [5:0] trunc_ln150_reg_440;
reg   [5:0] trunc_ln150_reg_440_pp0_iter1_reg;
reg   [5:0] trunc_ln150_reg_440_pp0_iter2_reg;
reg   [5:0] trunc_ln150_reg_440_pp0_iter3_reg;
reg   [5:0] trunc_ln150_reg_440_pp0_iter4_reg;
reg   [5:0] trunc_ln150_reg_440_pp0_iter5_reg;
reg   [5:0] trunc_ln150_reg_440_pp0_iter6_reg;
wire   [6:0] add_ln149_fu_233_p2;
wire   [8:0] select_ln148_24_fu_245_p3;
wire   [1:0] select_ln147_23_fu_287_p3;
reg   [1:0] select_ln147_23_reg_455;
reg    ap_enable_reg_pp0_iter1;
wire   [3:0] select_ln148_23_fu_370_p3;
reg   [3:0] select_ln148_23_reg_460;
reg   [3:0] select_ln148_23_reg_460_pp0_iter2_reg;
reg   [3:0] select_ln148_23_reg_460_pp0_iter3_reg;
reg   [3:0] select_ln148_23_reg_460_pp0_iter4_reg;
reg   [3:0] select_ln148_23_reg_460_pp0_iter5_reg;
reg   [3:0] select_ln148_23_reg_460_pp0_iter6_reg;
reg   [15:0] ifmap_vec_load_reg_475;
reg   [15:0] weight_vecs_0_load_reg_480;
wire   [15:0] grp_fu_153_p2;
reg   [15:0] mul_reg_485;
reg    ap_block_state1;
wire    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_flush_enable;
reg    ap_enable_reg_pp0_iter2;
reg    ap_condition_pp0_exit_iter1_state3;
reg    ap_enable_reg_pp0_iter3;
reg    ap_enable_reg_pp0_iter4;
reg    ap_enable_reg_pp0_iter5;
reg    ap_enable_reg_pp0_iter6;
reg    ap_enable_reg_pp0_iter7;
reg   [1:0] ap_phi_mux_jj_phi_fu_123_p4;
wire    ap_block_pp0_stage0;
reg   [1:0] ap_phi_mux_ii_phi_fu_146_p4;
wire   [63:0] p_cast25_fu_386_p1;
wire   [63:0] idxprom30_fu_398_p1;
wire   [0:0] icmp_ln149_fu_189_p2;
wire   [0:0] xor_ln147_fu_183_p2;
wire   [1:0] select_ln147_fu_175_p3;
wire   [0:0] or_ln148_fu_207_p2;
wire   [8:0] add_ln148_8_fu_239_p2;
wire   [3:0] shl_ln_fu_257_p3;
wire   [3:0] zext_ln150_fu_253_p1;
wire   [3:0] sub_ln150_fu_265_p2;
wire   [3:0] zext_ln150_11_fu_271_p1;
wire   [1:0] add_ln147_fu_281_p2;
wire   [3:0] tmp_fu_298_p3;
wire   [3:0] select_ln147_30_cast_fu_294_p1;
wire   [3:0] shl_ln150_mid1_fu_316_p3;
wire   [3:0] zext_ln150_17_fu_312_p1;
wire   [3:0] sub_ln150_10_fu_324_p2;
wire   [3:0] add_ln150_fu_275_p2;
wire   [3:0] empty_150_fu_306_p2;
wire   [3:0] select_ln148_29_cast_fu_344_p1;
wire   [3:0] empty_151_fu_347_p2;
wire   [3:0] select_ln147_24_fu_330_p3;
wire   [3:0] zext_ln150_18_fu_361_p1;
wire   [3:0] add_ln150_9_fu_364_p2;
wire   [3:0] select_ln147_25_fu_337_p3;
wire   [9:0] tmp_203_cast_fu_353_p3;
wire   [9:0] select_ln148_cast_fu_377_p1;
wire   [9:0] empty_152_fu_380_p2;
wire   [9:0] p_fu_392_p3;
wire    ap_CS_fsm_state10;
reg   [2:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
#0 ap_enable_reg_pp0_iter4 = 1'b0;
#0 ap_enable_reg_pp0_iter5 = 1'b0;
#0 ap_enable_reg_pp0_iter6 = 1'b0;
#0 ap_enable_reg_pp0_iter7 = 1'b0;
end

td_fused_top_hmul_16ns_16ns_16_4_max_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hmul_16ns_16ns_16_4_max_dsp_1_U618(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(ifmap_vec_load_reg_475),
    .din1(weight_vecs_0_load_reg_480),
    .dout(grp_fu_153_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state10)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if ((1'b1 == ap_condition_pp0_flush_enable)) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            if ((1'b1 == ap_condition_pp0_exit_iter1_state3)) begin
                ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter0;
            end else if ((1'b1 == 1'b1)) begin
                ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
            end
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter4 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter5 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter5 <= ap_enable_reg_pp0_iter4;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter6 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter6 <= ap_enable_reg_pp0_iter5;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter7 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter7 <= ap_enable_reg_pp0_iter6;
        end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter7 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_fu_163_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ic_reg_131 <= add_ln149_fu_233_p2;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ic_reg_131 <= 7'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_reg_408_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        ii_reg_142 <= select_ln147_23_reg_455;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ii_reg_142 <= 2'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_fu_163_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        indvar_flatten17_reg_97 <= add_ln147_8_fu_157_p2;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indvar_flatten17_reg_97 <= 10'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_fu_163_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        indvar_flatten_reg_108 <= select_ln148_24_fu_245_p3;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indvar_flatten_reg_108 <= 9'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_reg_408 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        jj_reg_119 <= select_ln148_22_reg_434;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        jj_reg_119 <= 2'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_fu_163_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        add_ln148_reg_424 <= add_ln148_fu_201_p2;
        and_ln147_reg_419 <= and_ln147_fu_195_p2;
        icmp_ln148_reg_412 <= icmp_ln148_fu_169_p2;
        select_ln148_reg_429 <= select_ln148_fu_213_p3;
        trunc_ln150_reg_440 <= trunc_ln150_fu_229_p1;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln147_reg_408 <= icmp_ln147_fu_163_p2;
        icmp_ln147_reg_408_pp0_iter1_reg <= icmp_ln147_reg_408;
        trunc_ln150_reg_440_pp0_iter1_reg <= trunc_ln150_reg_440;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        icmp_ln147_reg_408_pp0_iter2_reg <= icmp_ln147_reg_408_pp0_iter1_reg;
        icmp_ln147_reg_408_pp0_iter3_reg <= icmp_ln147_reg_408_pp0_iter2_reg;
        icmp_ln147_reg_408_pp0_iter4_reg <= icmp_ln147_reg_408_pp0_iter3_reg;
        icmp_ln147_reg_408_pp0_iter5_reg <= icmp_ln147_reg_408_pp0_iter4_reg;
        icmp_ln147_reg_408_pp0_iter6_reg <= icmp_ln147_reg_408_pp0_iter5_reg;
        select_ln148_23_reg_460_pp0_iter2_reg <= select_ln148_23_reg_460;
        select_ln148_23_reg_460_pp0_iter3_reg <= select_ln148_23_reg_460_pp0_iter2_reg;
        select_ln148_23_reg_460_pp0_iter4_reg <= select_ln148_23_reg_460_pp0_iter3_reg;
        select_ln148_23_reg_460_pp0_iter5_reg <= select_ln148_23_reg_460_pp0_iter4_reg;
        select_ln148_23_reg_460_pp0_iter6_reg <= select_ln148_23_reg_460_pp0_iter5_reg;
        trunc_ln150_reg_440_pp0_iter2_reg <= trunc_ln150_reg_440_pp0_iter1_reg;
        trunc_ln150_reg_440_pp0_iter3_reg <= trunc_ln150_reg_440_pp0_iter2_reg;
        trunc_ln150_reg_440_pp0_iter4_reg <= trunc_ln150_reg_440_pp0_iter3_reg;
        trunc_ln150_reg_440_pp0_iter5_reg <= trunc_ln150_reg_440_pp0_iter4_reg;
        trunc_ln150_reg_440_pp0_iter6_reg <= trunc_ln150_reg_440_pp0_iter5_reg;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_reg_408_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        ifmap_vec_load_reg_475 <= ifmap_vec_q0;
        weight_vecs_0_load_reg_480 <= weight_vecs_0_q0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_reg_408_pp0_iter5_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        mul_reg_485 <= grp_fu_153_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_reg_408 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        select_ln147_23_reg_455 <= select_ln147_23_fu_287_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_fu_163_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        select_ln148_22_reg_434 <= select_ln148_22_fu_221_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_reg_408 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        select_ln148_23_reg_460 <= select_ln148_23_fu_370_p3;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_condition_pp0_exit_iter1_state3 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter1_state3 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln147_fu_163_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_condition_pp0_flush_enable = 1'b1;
    end else begin
        ap_condition_pp0_flush_enable = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state10)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter7 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln147_reg_408_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        ap_phi_mux_ii_phi_fu_146_p4 = select_ln147_23_reg_455;
    end else begin
        ap_phi_mux_ii_phi_fu_146_p4 = ii_reg_142;
    end
end

always @ (*) begin
    if (((icmp_ln147_reg_408 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_jj_phi_fu_123_p4 = select_ln148_22_reg_434;
    end else begin
        ap_phi_mux_jj_phi_fu_123_p4 = jj_reg_119;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state10)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ifmap_vec_ce0 = 1'b1;
    end else begin
        ifmap_vec_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter7 == 1'b1))) begin
        products_0_ce0 = 1'b1;
    end else begin
        products_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln147_reg_408_pp0_iter6_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter7 == 1'b1))) begin
        products_0_we0 = 1'b1;
    end else begin
        products_0_we0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        weight_vecs_0_ce0 = 1'b1;
    end else begin
        weight_vecs_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((~((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b1)) & ~((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter7 == 1'b1) & (ap_enable_reg_pp0_iter6 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if ((((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter7 == 1'b1) & (ap_enable_reg_pp0_iter6 == 1'b0)) | ((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b1)))) begin
                ap_NS_fsm = ap_ST_fsm_state10;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state10 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln147_8_fu_157_p2 = (indvar_flatten17_reg_97 + 10'd1);

assign add_ln147_fu_281_p2 = (ap_phi_mux_ii_phi_fu_146_p4 + 2'd1);

assign add_ln148_8_fu_239_p2 = (indvar_flatten_reg_108 + 9'd1);

assign add_ln148_fu_201_p2 = (select_ln147_fu_175_p3 + 2'd1);

assign add_ln149_fu_233_p2 = (select_ln148_fu_213_p3 + 7'd1);

assign add_ln150_9_fu_364_p2 = (select_ln147_24_fu_330_p3 + zext_ln150_18_fu_361_p1);

assign add_ln150_fu_275_p2 = (sub_ln150_fu_265_p2 + zext_ln150_11_fu_271_p1);

assign and_ln147_fu_195_p2 = (xor_ln147_fu_183_p2 & icmp_ln149_fu_189_p2);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state10 = ap_CS_fsm[32'd2];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (ap_done_reg == 1'b1));
end

assign ap_block_state2_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter4 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage0_iter5 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage0_iter6 = ~(1'b1 == 1'b1);

assign ap_block_state9_pp0_stage0_iter7 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign empty_150_fu_306_p2 = (tmp_fu_298_p3 - select_ln147_30_cast_fu_294_p1);

assign empty_151_fu_347_p2 = (empty_150_fu_306_p2 + select_ln148_29_cast_fu_344_p1);

assign empty_152_fu_380_p2 = (tmp_203_cast_fu_353_p3 + select_ln148_cast_fu_377_p1);

assign icmp_ln147_fu_163_p2 = ((indvar_flatten17_reg_97 == 10'd576) ? 1'b1 : 1'b0);

assign icmp_ln148_fu_169_p2 = ((indvar_flatten_reg_108 == 9'd192) ? 1'b1 : 1'b0);

assign icmp_ln149_fu_189_p2 = ((ic_reg_131 == 7'd64) ? 1'b1 : 1'b0);

assign idxprom30_fu_398_p1 = p_fu_392_p3;

assign ifmap_vec_address0 = p_cast25_fu_386_p1;

assign or_ln148_fu_207_p2 = (icmp_ln148_fu_169_p2 | and_ln147_fu_195_p2);

assign p_cast25_fu_386_p1 = empty_152_fu_380_p2;

assign p_fu_392_p3 = {{select_ln148_23_reg_460_pp0_iter6_reg}, {trunc_ln150_reg_440_pp0_iter6_reg}};

assign products_0_address0 = idxprom30_fu_398_p1;

assign products_0_d0 = mul_reg_485;

assign select_ln147_23_fu_287_p3 = ((icmp_ln148_reg_412[0:0] == 1'b1) ? add_ln147_fu_281_p2 : ap_phi_mux_ii_phi_fu_146_p4);

assign select_ln147_24_fu_330_p3 = ((icmp_ln148_reg_412[0:0] == 1'b1) ? sub_ln150_10_fu_324_p2 : sub_ln150_fu_265_p2);

assign select_ln147_25_fu_337_p3 = ((icmp_ln148_reg_412[0:0] == 1'b1) ? sub_ln150_10_fu_324_p2 : add_ln150_fu_275_p2);

assign select_ln147_30_cast_fu_294_p1 = select_ln147_23_fu_287_p3;

assign select_ln147_fu_175_p3 = ((icmp_ln148_fu_169_p2[0:0] == 1'b1) ? 2'd0 : ap_phi_mux_jj_phi_fu_123_p4);

assign select_ln148_22_fu_221_p3 = ((and_ln147_fu_195_p2[0:0] == 1'b1) ? add_ln148_fu_201_p2 : select_ln147_fu_175_p3);

assign select_ln148_23_fu_370_p3 = ((and_ln147_reg_419[0:0] == 1'b1) ? add_ln150_9_fu_364_p2 : select_ln147_25_fu_337_p3);

assign select_ln148_24_fu_245_p3 = ((icmp_ln148_fu_169_p2[0:0] == 1'b1) ? 9'd1 : add_ln148_8_fu_239_p2);

assign select_ln148_29_cast_fu_344_p1 = select_ln148_22_reg_434;

assign select_ln148_cast_fu_377_p1 = select_ln148_reg_429;

assign select_ln148_fu_213_p3 = ((or_ln148_fu_207_p2[0:0] == 1'b1) ? 7'd0 : ic_reg_131);

assign shl_ln150_mid1_fu_316_p3 = {{add_ln147_fu_281_p2}, {2'd0}};

assign shl_ln_fu_257_p3 = {{ap_phi_mux_ii_phi_fu_146_p4}, {2'd0}};

assign sub_ln150_10_fu_324_p2 = (shl_ln150_mid1_fu_316_p3 - zext_ln150_17_fu_312_p1);

assign sub_ln150_fu_265_p2 = (shl_ln_fu_257_p3 - zext_ln150_fu_253_p1);

assign tmp_203_cast_fu_353_p3 = {{empty_151_fu_347_p2}, {6'd0}};

assign tmp_fu_298_p3 = {{select_ln147_23_fu_287_p3}, {2'd0}};

assign trunc_ln150_fu_229_p1 = select_ln148_fu_213_p3[5:0];

assign weight_vecs_0_address0 = p_cast25_fu_386_p1;

assign xor_ln147_fu_183_p2 = (icmp_ln148_fu_169_p2 ^ 1'd1);

assign zext_ln150_11_fu_271_p1 = jj_reg_119;

assign zext_ln150_17_fu_312_p1 = add_ln147_fu_281_p2;

assign zext_ln150_18_fu_361_p1 = add_ln148_reg_424;

assign zext_ln150_fu_253_p1 = ap_phi_mux_ii_phi_fu_146_p4;

endmodule //td_fused_top_tdf10_dot_product
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_tdf10_filters_ram (addr0, ce0, q0, addr1, ce1, d1, we1,  clk);

parameter DWIDTH = 64;
parameter AWIDTH = 17;
parameter MEM_SIZE = 73728;

input[AWIDTH-1:0] addr0;
input ce0;
output wire[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
input clk;

 reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];
wire [AWIDTH-1:0] addr0_t0; 
reg [AWIDTH-1:0] addr0_t1; 
reg [DWIDTH-1:0] q0_t0;
  reg [DWIDTH-1:0] q0_t1;
wire [AWIDTH-1:0] addr1_t0; 
reg [AWIDTH-1:0] addr1_t1; 
wire [DWIDTH-1:0] d1_t0; 
wire we1_t0; 
reg [DWIDTH-1:0] d1_t1; 
reg we1_t1; 


assign addr0_t0 = addr0;
assign q0 = q0_t1;
assign addr1_t0 = addr1;
assign d1_t0 = d1;
assign we1_t0 = we1;

always @(posedge clk)  
begin
    if (ce0) 
    begin
        addr0_t1 <= addr0_t0; 
        q0_t1 <= q0_t0;
    end
    if (ce1) 
    begin
        addr1_t1 <= addr1_t0; 
        d1_t1 <= d1_t0;
        we1_t1 <= we1_t0;
    end
end


always @(posedge clk)  
begin 
    if (ce0) begin
        q0_t0 <= ram[addr0_t1];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1_t1) 
            ram[addr1_t1] <= d1_t1; 
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_tdf10_filters(
    reset,
    clk,
    address0,
    ce0,
    q0,
    address1,
    ce1,
    we1,
    d1);

parameter DataWidth = 32'd64;
parameter AddressRange = 32'd73728;
parameter AddressWidth = 32'd17;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;



td_fused_top_tdf10_filters_ram td_fused_top_tdf10_filters_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 )
);

endmodule

// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf10_get_next_ijk (
        ap_clk,
        ap_rst,
        ap_start,
        start_full_n,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        start_out,
        start_write,
        indices_0_din,
        indices_0_full_n,
        indices_0_write,
        indices_1_din,
        indices_1_full_n,
        indices_1_write,
        indices_2_out_din,
        indices_2_out_full_n,
        indices_2_out_write,
        indices_2_out1_din,
        indices_2_out1_full_n,
        indices_2_out1_write,
        write_r_din,
        write_r_full_n,
        write_r_write
);

parameter    ap_ST_fsm_state1 = 1'd1;

input   ap_clk;
input   ap_rst;
input   ap_start;
input   start_full_n;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output   start_out;
output   start_write;
output  [15:0] indices_0_din;
input   indices_0_full_n;
output   indices_0_write;
output  [15:0] indices_1_din;
input   indices_1_full_n;
output   indices_1_write;
output  [8:0] indices_2_out_din;
input   indices_2_out_full_n;
output   indices_2_out_write;
output  [14:0] indices_2_out1_din;
input   indices_2_out1_full_n;
output   indices_2_out1_write;
output   write_r_din;
input   write_r_full_n;
output   write_r_write;

reg ap_done;
reg ap_idle;
reg start_write;
reg indices_0_write;
reg indices_1_write;
reg indices_2_out_write;
reg indices_2_out1_write;
reg write_r_write;

reg    real_start;
reg    start_once_reg;
reg    ap_done_reg;
  reg   [0:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    internal_ap_ready;
reg   [15:0] i_10;
reg   [15:0] j_10;
reg   [15:0] k_10;
reg    indices_0_blk_n;
reg    indices_1_blk_n;
reg    indices_2_out_blk_n;
reg    indices_2_out1_blk_n;
reg    write_r_blk_n;
reg   [0:0] ap_phi_mux_j_19_flag_0_i_phi_fu_92_p6;
reg    ap_block_state1;
wire   [0:0] icmp_ln188_fu_167_p2;
wire   [0:0] icmp_ln191_fu_180_p2;
reg   [15:0] ap_phi_mux_j_19_new_0_i_phi_fu_106_p6;
wire   [15:0] add_ln190_fu_173_p2;
reg   [15:0] ap_phi_mux_k_19_new_0_i_phi_fu_119_p6;
wire   [15:0] add_ln187_fu_160_p2;
wire   [15:0] select_ln194_fu_198_p3;
wire   [15:0] add_ln193_fu_186_p2;
wire   [0:0] icmp_ln194_fu_192_p2;
reg   [0:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 start_once_reg = 1'b0;
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 1'd1;
#0 i_10 = 16'd0;
#0 j_10 = 16'd0;
#0 k_10 = 16'd0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((~((real_start == 1'b0) | (write_r_full_n == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        start_once_reg <= 1'b0;
    end else begin
        if (((real_start == 1'b1) & (internal_ap_ready == 1'b0))) begin
            start_once_reg <= 1'b1;
        end else if ((internal_ap_ready == 1'b1)) begin
            start_once_reg <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((~((real_start == 1'b0) | (write_r_full_n == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (icmp_ln191_fu_180_p2 == 1'd1) & (icmp_ln188_fu_167_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1))) begin
        i_10 <= select_ln194_fu_198_p3;
    end
end

always @ (posedge ap_clk) begin
    if ((~((real_start == 1'b0) | (write_r_full_n == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (ap_phi_mux_j_19_flag_0_i_phi_fu_92_p6 == 1'd1) & (1'b1 == ap_CS_fsm_state1))) begin
        j_10 <= ap_phi_mux_j_19_new_0_i_phi_fu_106_p6;
    end
end

always @ (posedge ap_clk) begin
    if ((~((real_start == 1'b0) | (write_r_full_n == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        k_10 <= ap_phi_mux_k_19_new_0_i_phi_fu_119_p6;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (write_r_full_n == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((real_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln188_fu_167_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_phi_mux_j_19_flag_0_i_phi_fu_92_p6 = 1'd0;
    end else if ((((icmp_ln191_fu_180_p2 == 1'd0) & (icmp_ln188_fu_167_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1)) | ((icmp_ln191_fu_180_p2 == 1'd1) & (icmp_ln188_fu_167_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1)))) begin
        ap_phi_mux_j_19_flag_0_i_phi_fu_92_p6 = 1'd1;
    end else begin
        ap_phi_mux_j_19_flag_0_i_phi_fu_92_p6 = 'bx;
    end
end

always @ (*) begin
    if (((icmp_ln188_fu_167_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1))) begin
        if ((icmp_ln191_fu_180_p2 == 1'd0)) begin
            ap_phi_mux_j_19_new_0_i_phi_fu_106_p6 = add_ln190_fu_173_p2;
        end else if ((icmp_ln191_fu_180_p2 == 1'd1)) begin
            ap_phi_mux_j_19_new_0_i_phi_fu_106_p6 = 16'd0;
        end else begin
            ap_phi_mux_j_19_new_0_i_phi_fu_106_p6 = 'bx;
        end
    end else begin
        ap_phi_mux_j_19_new_0_i_phi_fu_106_p6 = 'bx;
    end
end

always @ (*) begin
    if (((icmp_ln188_fu_167_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_phi_mux_k_19_new_0_i_phi_fu_119_p6 = add_ln187_fu_160_p2;
    end else if ((((icmp_ln191_fu_180_p2 == 1'd0) & (icmp_ln188_fu_167_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1)) | ((icmp_ln191_fu_180_p2 == 1'd1) & (icmp_ln188_fu_167_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1)))) begin
        ap_phi_mux_k_19_new_0_i_phi_fu_119_p6 = 16'd0;
    end else begin
        ap_phi_mux_k_19_new_0_i_phi_fu_119_p6 = 'bx;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_0_blk_n = indices_0_full_n;
    end else begin
        indices_0_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (write_r_full_n == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_0_write = 1'b1;
    end else begin
        indices_0_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_1_blk_n = indices_1_full_n;
    end else begin
        indices_1_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (write_r_full_n == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_1_write = 1'b1;
    end else begin
        indices_1_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_2_out1_blk_n = indices_2_out1_full_n;
    end else begin
        indices_2_out1_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (write_r_full_n == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_2_out1_write = 1'b1;
    end else begin
        indices_2_out1_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_2_out_blk_n = indices_2_out_full_n;
    end else begin
        indices_2_out_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (write_r_full_n == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_2_out_write = 1'b1;
    end else begin
        indices_2_out_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (write_r_full_n == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        internal_ap_ready = 1'b1;
    end else begin
        internal_ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((start_full_n == 1'b0) & (start_once_reg == 1'b0))) begin
        real_start = 1'b0;
    end else begin
        real_start = ap_start;
    end
end

always @ (*) begin
    if (((real_start == 1'b1) & (start_once_reg == 1'b0))) begin
        start_write = 1'b1;
    end else begin
        start_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        write_r_blk_n = write_r_full_n;
    end else begin
        write_r_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (write_r_full_n == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        write_r_write = 1'b1;
    end else begin
        write_r_write = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln187_fu_160_p2 = (k_10 + 16'd1);

assign add_ln190_fu_173_p2 = (j_10 + 16'd1);

assign add_ln193_fu_186_p2 = (i_10 + 16'd1);

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

always @ (*) begin
    ap_block_state1 = ((real_start == 1'b0) | (write_r_full_n == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1));
end

assign ap_ready = internal_ap_ready;

assign icmp_ln188_fu_167_p2 = ((add_ln187_fu_160_p2 == 16'd512) ? 1'b1 : 1'b0);

assign icmp_ln191_fu_180_p2 = ((add_ln190_fu_173_p2 == 16'd14) ? 1'b1 : 1'b0);

assign icmp_ln194_fu_192_p2 = ((add_ln193_fu_186_p2 == 16'd14) ? 1'b1 : 1'b0);

assign indices_0_din = i_10;

assign indices_1_din = j_10;

assign indices_2_out1_din = k_10[14:0];

assign indices_2_out_din = k_10[8:0];

assign select_ln194_fu_198_p3 = ((icmp_ln194_fu_192_p2[0:0] == 1'b1) ? 16'd0 : add_ln193_fu_186_p2);

assign start_out = real_start;

assign write_r_din = ((k_10 == 16'd511) ? 1'b1 : 1'b0);

endmodule //td_fused_top_tdf10_get_next_ijk
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_tdf10_l2_filters_ram (addr0, ce0, q0, addr1, ce1, d1, we1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 15;
parameter MEM_SIZE = 32768;

input[AWIDTH-1:0] addr0;
input ce0;
output wire[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
input clk;

 reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];
wire [AWIDTH-1:0] addr0_t0; 
reg [AWIDTH-1:0] addr0_t1; 
reg [DWIDTH-1:0] q0_t0;
reg [DWIDTH-1:0] q0_t1;
wire [AWIDTH-1:0] addr1_t0; 
reg [AWIDTH-1:0] addr1_t1; 
wire [DWIDTH-1:0] d1_t0; 
wire we1_t0; 
reg [DWIDTH-1:0] d1_t1; 
reg we1_t1; 


assign addr0_t0 = addr0;
assign q0 = q0_t1;
assign addr1_t0 = addr1;
assign d1_t0 = d1;
assign we1_t0 = we1;

always @(posedge clk)  
begin
    if (ce0) 
    begin
        addr0_t1 <= addr0_t0; 
        q0_t1 <= q0_t0;
    end
    if (ce1) 
    begin
        addr1_t1 <= addr1_t0; 
        d1_t1 <= d1_t0;
        we1_t1 <= we1_t0;
    end
end


always @(posedge clk)  
begin 
    if (ce0) begin
        q0_t0 <= ram[addr0_t1];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1_t1) 
            ram[addr1_t1] <= d1_t1; 
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_tdf10_l2_filters(
    reset,
    clk,
    address0,
    ce0,
    q0,
    address1,
    ce1,
    we1,
    d1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd32768;
parameter AddressWidth = 32'd15;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;



td_fused_top_tdf10_l2_filters_ram td_fused_top_tdf10_l2_filters_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 )
);

endmodule

// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf10_l2_multiply66 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        intermediate_fmaps_read,
        l2_filter_data_address0,
        l2_filter_data_ce0,
        l2_filter_data_q0,
        l2_products_address0,
        l2_products_ce0,
        l2_products_we0,
        l2_products_d0,
        indices_23_dout,
        indices_23_empty_n,
        indices_23_read
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state10 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
input  [15:0] intermediate_fmaps_read;
output  [14:0] l2_filter_data_address0;
output   l2_filter_data_ce0;
input  [15:0] l2_filter_data_q0;
output  [5:0] l2_products_address0;
output   l2_products_ce0;
output   l2_products_we0;
output  [15:0] l2_products_d0;
input  [14:0] indices_23_dout;
input   indices_23_empty_n;
output   indices_23_read;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg l2_filter_data_ce0;
reg l2_products_ce0;
reg l2_products_we0;
reg indices_23_read;

reg    ap_done_reg;
  reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    indices_23_blk_n;
reg   [6:0] i_1_1_reg_106;
reg   [14:0] l2_ichan_reg_165;
wire   [6:0] add_ln20_fu_122_p2;
wire    ap_CS_fsm_pp0_stage0;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
wire    ap_block_state4_pp0_stage0_iter2;
wire    ap_block_state5_pp0_stage0_iter3;
wire    ap_block_state6_pp0_stage0_iter4;
wire    ap_block_state7_pp0_stage0_iter5;
wire    ap_block_state8_pp0_stage0_iter6;
wire    ap_block_state9_pp0_stage0_iter7;
wire    ap_block_pp0_stage0_11001;
wire   [0:0] icmp_ln20_fu_128_p2;
reg   [0:0] icmp_ln20_reg_175;
reg   [0:0] icmp_ln20_reg_175_pp0_iter1_reg;
reg   [0:0] icmp_ln20_reg_175_pp0_iter2_reg;
reg   [0:0] icmp_ln20_reg_175_pp0_iter3_reg;
reg   [0:0] icmp_ln20_reg_175_pp0_iter4_reg;
reg   [0:0] icmp_ln20_reg_175_pp0_iter5_reg;
reg   [0:0] icmp_ln20_reg_175_pp0_iter6_reg;
wire   [5:0] l2_o_fu_134_p1;
reg   [5:0] l2_o_reg_179;
reg   [5:0] l2_o_reg_179_pp0_iter1_reg;
reg   [5:0] l2_o_reg_179_pp0_iter2_reg;
reg   [5:0] l2_o_reg_179_pp0_iter3_reg;
reg   [5:0] l2_o_reg_179_pp0_iter4_reg;
reg   [5:0] l2_o_reg_179_pp0_iter5_reg;
reg   [5:0] l2_o_reg_179_pp0_iter6_reg;
wire   [15:0] grp_fu_117_p2;
reg   [15:0] mul_i_i_reg_194;
reg    ap_block_state1;
wire    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_exit_iter0_state2;
reg    ap_enable_reg_pp0_iter1;
reg    ap_enable_reg_pp0_iter2;
reg    ap_enable_reg_pp0_iter3;
reg    ap_enable_reg_pp0_iter4;
reg    ap_enable_reg_pp0_iter5;
reg    ap_enable_reg_pp0_iter6;
reg    ap_enable_reg_pp0_iter7;
wire   [63:0] zext_ln29_26_fu_151_p1;
wire    ap_block_pp0_stage0;
wire   [63:0] zext_ln29_fu_156_p1;
wire   [14:0] tmp_s_fu_138_p3;
wire   [14:0] add_ln29_fu_146_p2;
wire    ap_CS_fsm_state10;
reg   [2:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
#0 ap_enable_reg_pp0_iter4 = 1'b0;
#0 ap_enable_reg_pp0_iter5 = 1'b0;
#0 ap_enable_reg_pp0_iter6 = 1'b0;
#0 ap_enable_reg_pp0_iter7 = 1'b0;
end

td_fused_top_hmul_16ns_16ns_16_4_max_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hmul_16ns_16ns_16_4_max_dsp_1_U637(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(l2_filter_data_q0),
    .din1(intermediate_fmaps_read),
    .dout(grp_fu_117_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state10)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b1 == ap_condition_pp0_exit_iter0_state2))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            if ((1'b1 == ap_condition_pp0_exit_iter0_state2)) begin
                ap_enable_reg_pp0_iter1 <= (1'b1 ^ ap_condition_pp0_exit_iter0_state2);
            end else if ((1'b1 == 1'b1)) begin
                ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
            end
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter4 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter5 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter5 <= ap_enable_reg_pp0_iter4;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter6 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter6 <= ap_enable_reg_pp0_iter5;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter7 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter7 <= ap_enable_reg_pp0_iter6;
        end else if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter7 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        i_1_1_reg_106 <= 7'd0;
    end else if (((icmp_ln20_fu_128_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        i_1_1_reg_106 <= add_ln20_fu_122_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln20_reg_175 <= icmp_ln20_fu_128_p2;
        icmp_ln20_reg_175_pp0_iter1_reg <= icmp_ln20_reg_175;
        l2_o_reg_179_pp0_iter1_reg <= l2_o_reg_179;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        icmp_ln20_reg_175_pp0_iter2_reg <= icmp_ln20_reg_175_pp0_iter1_reg;
        icmp_ln20_reg_175_pp0_iter3_reg <= icmp_ln20_reg_175_pp0_iter2_reg;
        icmp_ln20_reg_175_pp0_iter4_reg <= icmp_ln20_reg_175_pp0_iter3_reg;
        icmp_ln20_reg_175_pp0_iter5_reg <= icmp_ln20_reg_175_pp0_iter4_reg;
        icmp_ln20_reg_175_pp0_iter6_reg <= icmp_ln20_reg_175_pp0_iter5_reg;
        l2_o_reg_179_pp0_iter2_reg <= l2_o_reg_179_pp0_iter1_reg;
        l2_o_reg_179_pp0_iter3_reg <= l2_o_reg_179_pp0_iter2_reg;
        l2_o_reg_179_pp0_iter4_reg <= l2_o_reg_179_pp0_iter3_reg;
        l2_o_reg_179_pp0_iter5_reg <= l2_o_reg_179_pp0_iter4_reg;
        l2_o_reg_179_pp0_iter6_reg <= l2_o_reg_179_pp0_iter5_reg;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state1)) begin
        l2_ichan_reg_165 <= indices_23_dout;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln20_fu_128_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        l2_o_reg_179 <= l2_o_fu_134_p1;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln20_reg_175_pp0_iter5_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        mul_i_i_reg_194 <= grp_fu_117_p2;
    end
end

always @ (*) begin
    if ((icmp_ln20_fu_128_p2 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state2 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state2 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state10)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter7 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state10)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_23_blk_n = indices_23_empty_n;
    end else begin
        indices_23_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_23_read = 1'b1;
    end else begin
        indices_23_read = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter3 == 1'b1)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1)))) begin
        l2_filter_data_ce0 = 1'b1;
    end else begin
        l2_filter_data_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter7 == 1'b1))) begin
        l2_products_ce0 = 1'b1;
    end else begin
        l2_products_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln20_reg_175_pp0_iter6_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter7 == 1'b1))) begin
        l2_products_we0 = 1'b1;
    end else begin
        l2_products_we0 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((~((icmp_ln20_fu_128_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0)) & ~((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter7 == 1'b1) & (ap_enable_reg_pp0_iter6 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if ((((icmp_ln20_fu_128_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0)) | ((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter7 == 1'b1) & (ap_enable_reg_pp0_iter6 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_state10;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state10 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln20_fu_122_p2 = (i_1_1_reg_106 + 7'd1);

assign add_ln29_fu_146_p2 = (tmp_s_fu_138_p3 + l2_ichan_reg_165);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state10 = ap_CS_fsm[32'd2];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1));
end

assign ap_block_state2_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter4 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage0_iter5 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage0_iter6 = ~(1'b1 == 1'b1);

assign ap_block_state9_pp0_stage0_iter7 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign icmp_ln20_fu_128_p2 = ((i_1_1_reg_106 == 7'd64) ? 1'b1 : 1'b0);

assign l2_filter_data_address0 = zext_ln29_26_fu_151_p1;

assign l2_o_fu_134_p1 = i_1_1_reg_106[5:0];

assign l2_products_address0 = zext_ln29_fu_156_p1;

assign l2_products_d0 = mul_i_i_reg_194;

assign tmp_s_fu_138_p3 = {{l2_o_fu_134_p1}, {9'd0}};

assign zext_ln29_26_fu_151_p1 = add_ln29_fu_146_p2;

assign zext_ln29_fu_156_p1 = l2_o_reg_179_pp0_iter6_reg;

endmodule //td_fused_top_tdf10_l2_multiply66
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_tdf10_l2_writeOutputs_165_running_sums_3_ram (addr0, ce0, d0, we0, addr1, ce1, q1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
input[AWIDTH-1:0] addr1;
input ce1;
output reg[DWIDTH-1:0] q1;
input clk;

 reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];

//initial begin
//    $readmemh("./td_fused_top_tdf10_l2_writeOutputs_165_running_sums_3_ram.dat", ram);
//end



always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        q1 <= ram[addr1];
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_tdf10_l2_writeOutputs_165_running_sums_3(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    address1,
    ce1,
    q1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
input[AddressWidth - 1:0] address1;
input ce1;
output[DataWidth - 1:0] q1;



td_fused_top_tdf10_l2_writeOutputs_165_running_sums_3_ram td_fused_top_tdf10_l2_writeOutputs_165_running_sums_3_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .q1( q1 )
);

endmodule

// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf10_l2_writeOutputs_165 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        indices_01_dout,
        indices_01_empty_n,
        indices_01_read,
        indices_12_dout,
        indices_12_empty_n,
        indices_12_read,
        write4_dout,
        write4_empty_n,
        write4_read,
        l2_partial_sums_address0,
        l2_partial_sums_ce0,
        l2_partial_sums_q0,
        out_data_address1,
        out_data_ce1,
        out_data_we1,
        out_data_d1,
        l2_adjustments_address0,
        l2_adjustments_ce0,
        l2_adjustments_q0
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state25 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
input  [3:0] indices_01_dout;
input   indices_01_empty_n;
output   indices_01_read;
input  [7:0] indices_12_dout;
input   indices_12_empty_n;
output   indices_12_read;
input  [0:0] write4_dout;
input   write4_empty_n;
output   write4_read;
output  [5:0] l2_partial_sums_address0;
output   l2_partial_sums_ce0;
input  [15:0] l2_partial_sums_q0;
output  [11:0] out_data_address1;
output   out_data_ce1;
output   out_data_we1;
output  [63:0] out_data_d1;
output  [5:0] l2_adjustments_address0;
output   l2_adjustments_ce0;
input  [47:0] l2_adjustments_q0;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg indices_01_read;
reg indices_12_read;
reg write4_read;
reg l2_partial_sums_ce0;
reg out_data_ce1;
reg out_data_we1;
reg l2_adjustments_ce0;

reg    ap_done_reg;
  reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    running_sums_3_ce0;
reg    running_sums_3_we0;
wire   [15:0] running_sums_3_d0;
wire   [5:0] running_sums_3_address1;
reg    running_sums_3_ce1;
wire   [15:0] running_sums_3_q1;
reg    indices_01_blk_n;
reg    indices_12_blk_n;
reg    write4_blk_n;
reg   [6:0] ochan_reg_208;
reg   [0:0] write4_read_reg_567;
wire   [9:0] add_ln109_fu_273_p2;
reg   [9:0] add_ln109_reg_573;
wire   [6:0] add_ln86_fu_279_p2;
wire    ap_CS_fsm_pp0_stage0;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
wire    ap_block_state4_pp0_stage0_iter2;
wire    ap_block_state5_pp0_stage0_iter3;
wire    ap_block_state6_pp0_stage0_iter4;
wire    ap_block_state7_pp0_stage0_iter5;
wire    ap_block_state8_pp0_stage0_iter6;
wire    ap_block_state9_pp0_stage0_iter7;
wire    ap_block_state10_pp0_stage0_iter8;
wire    ap_block_state11_pp0_stage0_iter9;
wire    ap_block_state12_pp0_stage0_iter10;
wire    ap_block_state13_pp0_stage0_iter11;
wire    ap_block_state14_pp0_stage0_iter12;
wire    ap_block_state15_pp0_stage0_iter13;
wire    ap_block_state16_pp0_stage0_iter14;
wire    ap_block_state17_pp0_stage0_iter15;
wire    ap_block_state18_pp0_stage0_iter16;
wire    ap_block_state19_pp0_stage0_iter17;
wire    ap_block_state20_pp0_stage0_iter18;
wire    ap_block_state21_pp0_stage0_iter19;
wire    ap_block_state22_pp0_stage0_iter20;
wire    ap_block_state23_pp0_stage0_iter21;
wire    ap_block_state24_pp0_stage0_iter22;
wire    ap_block_pp0_stage0_11001;
wire   [0:0] icmp_ln86_fu_285_p2;
wire   [63:0] zext_ln86_fu_291_p1;
reg   [63:0] zext_ln86_reg_587;
reg   [63:0] zext_ln86_reg_587_pp0_iter1_reg;
reg   [63:0] zext_ln86_reg_587_pp0_iter2_reg;
reg   [63:0] zext_ln86_reg_587_pp0_iter3_reg;
reg   [5:0] running_sums_3_addr_reg_597;
reg   [5:0] running_sums_3_addr_reg_597_pp0_iter1_reg;
reg   [5:0] running_sums_3_addr_reg_597_pp0_iter2_reg;
reg   [5:0] running_sums_3_addr_reg_597_pp0_iter3_reg;
reg   [5:0] running_sums_3_addr_reg_597_pp0_iter4_reg;
reg   [5:0] running_sums_3_addr_reg_597_pp0_iter5_reg;
reg   [5:0] running_sums_3_addr_reg_597_pp0_iter6_reg;
wire   [1:0] trunc_ln99_fu_297_p1;
reg   [1:0] trunc_ln99_reg_603;
reg   [1:0] trunc_ln99_reg_603_pp0_iter1_reg;
reg   [1:0] trunc_ln99_reg_603_pp0_iter2_reg;
reg   [1:0] trunc_ln99_reg_603_pp0_iter3_reg;
reg   [1:0] trunc_ln99_reg_603_pp0_iter4_reg;
reg   [1:0] trunc_ln99_reg_603_pp0_iter5_reg;
reg   [1:0] trunc_ln99_reg_603_pp0_iter6_reg;
reg   [1:0] trunc_ln99_reg_603_pp0_iter7_reg;
reg   [1:0] trunc_ln99_reg_603_pp0_iter8_reg;
reg   [1:0] trunc_ln99_reg_603_pp0_iter9_reg;
reg   [1:0] trunc_ln99_reg_603_pp0_iter10_reg;
reg   [1:0] trunc_ln99_reg_603_pp0_iter11_reg;
reg   [1:0] trunc_ln99_reg_603_pp0_iter12_reg;
reg   [1:0] trunc_ln99_reg_603_pp0_iter13_reg;
reg   [1:0] trunc_ln99_reg_603_pp0_iter14_reg;
reg   [1:0] trunc_ln99_reg_603_pp0_iter15_reg;
reg   [1:0] trunc_ln99_reg_603_pp0_iter16_reg;
reg   [1:0] trunc_ln99_reg_603_pp0_iter17_reg;
reg   [1:0] trunc_ln99_reg_603_pp0_iter18_reg;
reg   [1:0] trunc_ln99_reg_603_pp0_iter19_reg;
reg   [1:0] trunc_ln99_reg_603_pp0_iter20_reg;
wire   [0:0] and_ln103_fu_307_p2;
reg   [0:0] and_ln103_reg_610;
reg   [0:0] and_ln103_reg_610_pp0_iter1_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter2_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter3_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter4_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter5_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter6_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter7_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter8_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter9_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter10_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter11_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter12_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter13_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter14_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter15_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter16_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter17_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter18_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter19_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter20_reg;
reg   [3:0] lshr_ln_reg_614;
reg   [3:0] lshr_ln_reg_614_pp0_iter1_reg;
reg   [3:0] lshr_ln_reg_614_pp0_iter2_reg;
reg   [3:0] lshr_ln_reg_614_pp0_iter3_reg;
reg   [3:0] lshr_ln_reg_614_pp0_iter4_reg;
reg   [3:0] lshr_ln_reg_614_pp0_iter5_reg;
reg   [3:0] lshr_ln_reg_614_pp0_iter6_reg;
reg   [3:0] lshr_ln_reg_614_pp0_iter7_reg;
reg   [3:0] lshr_ln_reg_614_pp0_iter8_reg;
reg   [3:0] lshr_ln_reg_614_pp0_iter9_reg;
reg   [3:0] lshr_ln_reg_614_pp0_iter10_reg;
reg   [3:0] lshr_ln_reg_614_pp0_iter11_reg;
reg   [3:0] lshr_ln_reg_614_pp0_iter12_reg;
reg   [3:0] lshr_ln_reg_614_pp0_iter13_reg;
reg   [3:0] lshr_ln_reg_614_pp0_iter14_reg;
reg   [3:0] lshr_ln_reg_614_pp0_iter15_reg;
reg   [3:0] lshr_ln_reg_614_pp0_iter16_reg;
reg   [3:0] lshr_ln_reg_614_pp0_iter17_reg;
reg   [3:0] lshr_ln_reg_614_pp0_iter18_reg;
reg   [3:0] lshr_ln_reg_614_pp0_iter19_reg;
reg   [3:0] lshr_ln_reg_614_pp0_iter20_reg;
reg   [15:0] val_reg_619;
reg   [15:0] running_sums_3_load_reg_624;
reg    ap_enable_reg_pp0_iter1;
wire   [15:0] grp_fu_219_p2;
reg   [15:0] sum_reg_634;
reg   [15:0] tmp_104_i_i_reg_645;
reg   [15:0] tmp_104_i_i_reg_645_pp0_iter8_reg;
reg   [15:0] tmp_104_i_i_reg_645_pp0_iter9_reg;
reg   [15:0] tmp_104_i_i_reg_645_pp0_iter10_reg;
reg   [15:0] tmp_104_i_i_reg_645_pp0_iter11_reg;
reg   [15:0] tmp_105_i_i_reg_650;
reg   [15:0] tmp_105_i_i_reg_650_pp0_iter8_reg;
reg   [15:0] tmp_105_i_i_reg_650_pp0_iter9_reg;
reg   [15:0] tmp_105_i_i_reg_650_pp0_iter10_reg;
reg   [15:0] tmp_105_i_i_reg_650_pp0_iter11_reg;
reg   [15:0] tmp_105_i_i_reg_650_pp0_iter12_reg;
reg   [15:0] tmp_105_i_i_reg_650_pp0_iter13_reg;
reg   [15:0] tmp_105_i_i_reg_650_pp0_iter14_reg;
reg   [15:0] tmp_105_i_i_reg_650_pp0_iter15_reg;
wire   [15:0] grp_fu_227_p2;
reg   [15:0] sub_i_i_i_reg_655;
wire   [15:0] grp_fu_231_p2;
reg   [15:0] normalized_reg_665;
wire   [15:0] grp_fu_223_p2;
reg   [15:0] biased_reg_675;
reg    ap_block_state1;
wire    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_exit_iter0_state2;
reg    ap_enable_reg_pp0_iter2;
reg    ap_enable_reg_pp0_iter3;
reg    ap_enable_reg_pp0_iter4;
reg    ap_enable_reg_pp0_iter5;
reg    ap_enable_reg_pp0_iter6;
reg    ap_enable_reg_pp0_iter7;
reg    ap_enable_reg_pp0_iter8;
reg    ap_enable_reg_pp0_iter9;
reg    ap_enable_reg_pp0_iter10;
reg    ap_enable_reg_pp0_iter11;
reg    ap_enable_reg_pp0_iter12;
reg    ap_enable_reg_pp0_iter13;
reg    ap_enable_reg_pp0_iter14;
reg    ap_enable_reg_pp0_iter15;
reg    ap_enable_reg_pp0_iter16;
reg    ap_enable_reg_pp0_iter17;
reg    ap_enable_reg_pp0_iter18;
reg    ap_enable_reg_pp0_iter19;
reg    ap_enable_reg_pp0_iter20;
reg    ap_enable_reg_pp0_iter21;
reg    ap_enable_reg_pp0_iter22;
wire    ap_block_pp0_stage0;
wire   [63:0] sext_ln109_fu_509_p1;
reg   [15:0] quad_3_39_fu_114;
wire   [15:0] quad_3_58_fu_475_p3;
reg   [15:0] quad_3_36_fu_118;
wire   [15:0] quad_3_57_fu_467_p3;
reg   [15:0] quad_3_40_fu_122;
wire   [15:0] quad_3_55_fu_451_p3;
reg   [15:0] quad_3_41_fu_126;
wire   [15:0] quad_3_52_fu_427_p3;
wire   [15:0] grp_fu_223_p1;
wire   [15:0] grp_fu_227_p1;
wire   [15:0] grp_fu_231_p1;
wire   [7:0] tmp_fu_235_p3;
wire   [4:0] tmp_s_fu_247_p3;
wire   [8:0] zext_ln109_fu_243_p1;
wire   [8:0] zext_ln109_7_fu_255_p1;
wire   [8:0] sub_ln109_fu_259_p2;
wire   [9:0] sub_ln109_cast_fu_265_p1;
wire   [9:0] zext_ln109_8_fu_269_p1;
wire   [0:0] icmp_ln103_fu_301_p2;
wire   [15:0] trunc_ln95_fu_329_p1;
wire   [15:0] data_V_fu_378_p1;
wire   [0:0] p_Result_s_fu_381_p3;
wire   [0:0] icmp_ln99_fu_396_p2;
wire   [15:0] quad_0_fu_389_p3;
wire   [0:0] icmp_ln99_7_fu_409_p2;
wire   [15:0] quad_3_fu_401_p3;
wire   [0:0] icmp_ln99_8_fu_422_p2;
wire   [15:0] quad_3_51_fu_414_p3;
wire   [15:0] quad_3_53_fu_435_p3;
wire   [15:0] quad_3_54_fu_443_p3;
wire   [15:0] quad_3_56_fu_459_p3;
wire   [13:0] tmp_74_fu_503_p3;
wire   [15:0] bitcast_ln109_12_fu_526_p1;
wire   [15:0] bitcast_ln109_11_fu_522_p1;
wire   [15:0] bitcast_ln109_10_fu_518_p1;
wire   [15:0] bitcast_ln109_fu_514_p1;
wire    ap_CS_fsm_state25;
reg   [2:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
#0 ap_enable_reg_pp0_iter4 = 1'b0;
#0 ap_enable_reg_pp0_iter5 = 1'b0;
#0 ap_enable_reg_pp0_iter6 = 1'b0;
#0 ap_enable_reg_pp0_iter7 = 1'b0;
#0 ap_enable_reg_pp0_iter8 = 1'b0;
#0 ap_enable_reg_pp0_iter9 = 1'b0;
#0 ap_enable_reg_pp0_iter10 = 1'b0;
#0 ap_enable_reg_pp0_iter11 = 1'b0;
#0 ap_enable_reg_pp0_iter12 = 1'b0;
#0 ap_enable_reg_pp0_iter13 = 1'b0;
#0 ap_enable_reg_pp0_iter14 = 1'b0;
#0 ap_enable_reg_pp0_iter15 = 1'b0;
#0 ap_enable_reg_pp0_iter16 = 1'b0;
#0 ap_enable_reg_pp0_iter17 = 1'b0;
#0 ap_enable_reg_pp0_iter18 = 1'b0;
#0 ap_enable_reg_pp0_iter19 = 1'b0;
#0 ap_enable_reg_pp0_iter20 = 1'b0;
#0 ap_enable_reg_pp0_iter21 = 1'b0;
#0 ap_enable_reg_pp0_iter22 = 1'b0;
end

td_fused_top_tdf10_l2_writeOutputs_165_running_sums_3 #(
    .DataWidth( 16 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
running_sums_3_U(
    .reset(ap_rst),
    .clk(ap_clk),
    .address0(running_sums_3_addr_reg_597_pp0_iter6_reg),
    .ce0(running_sums_3_ce0),
    .we0(running_sums_3_we0),
    .d0(running_sums_3_d0),
    .address1(running_sums_3_address1),
    .ce1(running_sums_3_ce1),
    .q1(running_sums_3_q1)
);

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U642(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(running_sums_3_load_reg_624),
    .din1(val_reg_619),
    .dout(grp_fu_219_p2)
);

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U643(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(normalized_reg_665),
    .din1(grp_fu_223_p1),
    .dout(grp_fu_223_p2)
);

td_fused_top_hsub_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hsub_16ns_16ns_16_5_full_dsp_1_U644(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(sum_reg_634),
    .din1(grp_fu_227_p1),
    .dout(grp_fu_227_p2)
);

td_fused_top_hmul_16ns_16ns_16_4_max_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hmul_16ns_16ns_16_4_max_dsp_1_U645(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(sub_i_i_i_reg_655),
    .din1(grp_fu_231_p1),
    .dout(grp_fu_231_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state25)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b1 == ap_condition_pp0_exit_iter0_state2) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((~((ap_start == 1'b0) | (write4_empty_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            if ((1'b1 == ap_condition_pp0_exit_iter0_state2)) begin
                ap_enable_reg_pp0_iter1 <= (1'b1 ^ ap_condition_pp0_exit_iter0_state2);
            end else if ((1'b1 == 1'b1)) begin
                ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
            end
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter10 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter10 <= ap_enable_reg_pp0_iter9;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter11 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter11 <= ap_enable_reg_pp0_iter10;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter12 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter12 <= ap_enable_reg_pp0_iter11;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter13 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter13 <= ap_enable_reg_pp0_iter12;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter14 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter14 <= ap_enable_reg_pp0_iter13;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter15 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter15 <= ap_enable_reg_pp0_iter14;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter16 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter16 <= ap_enable_reg_pp0_iter15;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter17 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter17 <= ap_enable_reg_pp0_iter16;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter18 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter18 <= ap_enable_reg_pp0_iter17;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter19 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter19 <= ap_enable_reg_pp0_iter18;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter20 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter20 <= ap_enable_reg_pp0_iter19;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter21 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter21 <= ap_enable_reg_pp0_iter20;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter22 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter22 <= ap_enable_reg_pp0_iter21;
        end else if ((~((ap_start == 1'b0) | (write4_empty_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter22 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter4 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter5 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter5 <= ap_enable_reg_pp0_iter4;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter6 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter6 <= ap_enable_reg_pp0_iter5;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter7 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter7 <= ap_enable_reg_pp0_iter6;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter8 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter8 <= ap_enable_reg_pp0_iter7;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter9 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter9 <= ap_enable_reg_pp0_iter8;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (icmp_ln86_fu_285_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        ochan_reg_208 <= add_ln86_fu_279_p2;
    end else if ((~((ap_start == 1'b0) | (write4_empty_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ochan_reg_208 <= 7'd0;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state1)) begin
        add_ln109_reg_573 <= add_ln109_fu_273_p2;
        write4_read_reg_567 <= write4_dout;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (icmp_ln86_fu_285_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        and_ln103_reg_610 <= and_ln103_fu_307_p2;
        running_sums_3_addr_reg_597 <= zext_ln86_fu_291_p1;
        trunc_ln99_reg_603 <= trunc_ln99_fu_297_p1;
        zext_ln86_reg_587[6 : 0] <= zext_ln86_fu_291_p1[6 : 0];
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        and_ln103_reg_610_pp0_iter10_reg <= and_ln103_reg_610_pp0_iter9_reg;
        and_ln103_reg_610_pp0_iter11_reg <= and_ln103_reg_610_pp0_iter10_reg;
        and_ln103_reg_610_pp0_iter12_reg <= and_ln103_reg_610_pp0_iter11_reg;
        and_ln103_reg_610_pp0_iter13_reg <= and_ln103_reg_610_pp0_iter12_reg;
        and_ln103_reg_610_pp0_iter14_reg <= and_ln103_reg_610_pp0_iter13_reg;
        and_ln103_reg_610_pp0_iter15_reg <= and_ln103_reg_610_pp0_iter14_reg;
        and_ln103_reg_610_pp0_iter16_reg <= and_ln103_reg_610_pp0_iter15_reg;
        and_ln103_reg_610_pp0_iter17_reg <= and_ln103_reg_610_pp0_iter16_reg;
        and_ln103_reg_610_pp0_iter18_reg <= and_ln103_reg_610_pp0_iter17_reg;
        and_ln103_reg_610_pp0_iter19_reg <= and_ln103_reg_610_pp0_iter18_reg;
        and_ln103_reg_610_pp0_iter20_reg <= and_ln103_reg_610_pp0_iter19_reg;
        and_ln103_reg_610_pp0_iter2_reg <= and_ln103_reg_610_pp0_iter1_reg;
        and_ln103_reg_610_pp0_iter3_reg <= and_ln103_reg_610_pp0_iter2_reg;
        and_ln103_reg_610_pp0_iter4_reg <= and_ln103_reg_610_pp0_iter3_reg;
        and_ln103_reg_610_pp0_iter5_reg <= and_ln103_reg_610_pp0_iter4_reg;
        and_ln103_reg_610_pp0_iter6_reg <= and_ln103_reg_610_pp0_iter5_reg;
        and_ln103_reg_610_pp0_iter7_reg <= and_ln103_reg_610_pp0_iter6_reg;
        and_ln103_reg_610_pp0_iter8_reg <= and_ln103_reg_610_pp0_iter7_reg;
        and_ln103_reg_610_pp0_iter9_reg <= and_ln103_reg_610_pp0_iter8_reg;
        biased_reg_675 <= grp_fu_223_p2;
        lshr_ln_reg_614_pp0_iter10_reg <= lshr_ln_reg_614_pp0_iter9_reg;
        lshr_ln_reg_614_pp0_iter11_reg <= lshr_ln_reg_614_pp0_iter10_reg;
        lshr_ln_reg_614_pp0_iter12_reg <= lshr_ln_reg_614_pp0_iter11_reg;
        lshr_ln_reg_614_pp0_iter13_reg <= lshr_ln_reg_614_pp0_iter12_reg;
        lshr_ln_reg_614_pp0_iter14_reg <= lshr_ln_reg_614_pp0_iter13_reg;
        lshr_ln_reg_614_pp0_iter15_reg <= lshr_ln_reg_614_pp0_iter14_reg;
        lshr_ln_reg_614_pp0_iter16_reg <= lshr_ln_reg_614_pp0_iter15_reg;
        lshr_ln_reg_614_pp0_iter17_reg <= lshr_ln_reg_614_pp0_iter16_reg;
        lshr_ln_reg_614_pp0_iter18_reg <= lshr_ln_reg_614_pp0_iter17_reg;
        lshr_ln_reg_614_pp0_iter19_reg <= lshr_ln_reg_614_pp0_iter18_reg;
        lshr_ln_reg_614_pp0_iter20_reg <= lshr_ln_reg_614_pp0_iter19_reg;
        lshr_ln_reg_614_pp0_iter2_reg <= lshr_ln_reg_614_pp0_iter1_reg;
        lshr_ln_reg_614_pp0_iter3_reg <= lshr_ln_reg_614_pp0_iter2_reg;
        lshr_ln_reg_614_pp0_iter4_reg <= lshr_ln_reg_614_pp0_iter3_reg;
        lshr_ln_reg_614_pp0_iter5_reg <= lshr_ln_reg_614_pp0_iter4_reg;
        lshr_ln_reg_614_pp0_iter6_reg <= lshr_ln_reg_614_pp0_iter5_reg;
        lshr_ln_reg_614_pp0_iter7_reg <= lshr_ln_reg_614_pp0_iter6_reg;
        lshr_ln_reg_614_pp0_iter8_reg <= lshr_ln_reg_614_pp0_iter7_reg;
        lshr_ln_reg_614_pp0_iter9_reg <= lshr_ln_reg_614_pp0_iter8_reg;
        normalized_reg_665 <= grp_fu_231_p2;
        running_sums_3_addr_reg_597_pp0_iter2_reg <= running_sums_3_addr_reg_597_pp0_iter1_reg;
        running_sums_3_addr_reg_597_pp0_iter3_reg <= running_sums_3_addr_reg_597_pp0_iter2_reg;
        running_sums_3_addr_reg_597_pp0_iter4_reg <= running_sums_3_addr_reg_597_pp0_iter3_reg;
        running_sums_3_addr_reg_597_pp0_iter5_reg <= running_sums_3_addr_reg_597_pp0_iter4_reg;
        running_sums_3_addr_reg_597_pp0_iter6_reg <= running_sums_3_addr_reg_597_pp0_iter5_reg;
        sub_i_i_i_reg_655 <= grp_fu_227_p2;
        sum_reg_634 <= grp_fu_219_p2;
        tmp_104_i_i_reg_645 <= {{l2_adjustments_q0[31:16]}};
        tmp_104_i_i_reg_645_pp0_iter10_reg <= tmp_104_i_i_reg_645_pp0_iter9_reg;
        tmp_104_i_i_reg_645_pp0_iter11_reg <= tmp_104_i_i_reg_645_pp0_iter10_reg;
        tmp_104_i_i_reg_645_pp0_iter8_reg <= tmp_104_i_i_reg_645;
        tmp_104_i_i_reg_645_pp0_iter9_reg <= tmp_104_i_i_reg_645_pp0_iter8_reg;
        tmp_105_i_i_reg_650 <= {{l2_adjustments_q0[47:32]}};
        tmp_105_i_i_reg_650_pp0_iter10_reg <= tmp_105_i_i_reg_650_pp0_iter9_reg;
        tmp_105_i_i_reg_650_pp0_iter11_reg <= tmp_105_i_i_reg_650_pp0_iter10_reg;
        tmp_105_i_i_reg_650_pp0_iter12_reg <= tmp_105_i_i_reg_650_pp0_iter11_reg;
        tmp_105_i_i_reg_650_pp0_iter13_reg <= tmp_105_i_i_reg_650_pp0_iter12_reg;
        tmp_105_i_i_reg_650_pp0_iter14_reg <= tmp_105_i_i_reg_650_pp0_iter13_reg;
        tmp_105_i_i_reg_650_pp0_iter15_reg <= tmp_105_i_i_reg_650_pp0_iter14_reg;
        tmp_105_i_i_reg_650_pp0_iter8_reg <= tmp_105_i_i_reg_650;
        tmp_105_i_i_reg_650_pp0_iter9_reg <= tmp_105_i_i_reg_650_pp0_iter8_reg;
        trunc_ln99_reg_603_pp0_iter10_reg <= trunc_ln99_reg_603_pp0_iter9_reg;
        trunc_ln99_reg_603_pp0_iter11_reg <= trunc_ln99_reg_603_pp0_iter10_reg;
        trunc_ln99_reg_603_pp0_iter12_reg <= trunc_ln99_reg_603_pp0_iter11_reg;
        trunc_ln99_reg_603_pp0_iter13_reg <= trunc_ln99_reg_603_pp0_iter12_reg;
        trunc_ln99_reg_603_pp0_iter14_reg <= trunc_ln99_reg_603_pp0_iter13_reg;
        trunc_ln99_reg_603_pp0_iter15_reg <= trunc_ln99_reg_603_pp0_iter14_reg;
        trunc_ln99_reg_603_pp0_iter16_reg <= trunc_ln99_reg_603_pp0_iter15_reg;
        trunc_ln99_reg_603_pp0_iter17_reg <= trunc_ln99_reg_603_pp0_iter16_reg;
        trunc_ln99_reg_603_pp0_iter18_reg <= trunc_ln99_reg_603_pp0_iter17_reg;
        trunc_ln99_reg_603_pp0_iter19_reg <= trunc_ln99_reg_603_pp0_iter18_reg;
        trunc_ln99_reg_603_pp0_iter20_reg <= trunc_ln99_reg_603_pp0_iter19_reg;
        trunc_ln99_reg_603_pp0_iter2_reg <= trunc_ln99_reg_603_pp0_iter1_reg;
        trunc_ln99_reg_603_pp0_iter3_reg <= trunc_ln99_reg_603_pp0_iter2_reg;
        trunc_ln99_reg_603_pp0_iter4_reg <= trunc_ln99_reg_603_pp0_iter3_reg;
        trunc_ln99_reg_603_pp0_iter5_reg <= trunc_ln99_reg_603_pp0_iter4_reg;
        trunc_ln99_reg_603_pp0_iter6_reg <= trunc_ln99_reg_603_pp0_iter5_reg;
        trunc_ln99_reg_603_pp0_iter7_reg <= trunc_ln99_reg_603_pp0_iter6_reg;
        trunc_ln99_reg_603_pp0_iter8_reg <= trunc_ln99_reg_603_pp0_iter7_reg;
        trunc_ln99_reg_603_pp0_iter9_reg <= trunc_ln99_reg_603_pp0_iter8_reg;
        zext_ln86_reg_587_pp0_iter2_reg[6 : 0] <= zext_ln86_reg_587_pp0_iter1_reg[6 : 0];
        zext_ln86_reg_587_pp0_iter3_reg[6 : 0] <= zext_ln86_reg_587_pp0_iter2_reg[6 : 0];
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        and_ln103_reg_610_pp0_iter1_reg <= and_ln103_reg_610;
        lshr_ln_reg_614_pp0_iter1_reg <= lshr_ln_reg_614;
        running_sums_3_addr_reg_597_pp0_iter1_reg <= running_sums_3_addr_reg_597;
        trunc_ln99_reg_603_pp0_iter1_reg <= trunc_ln99_reg_603;
        val_reg_619 <= l2_partial_sums_q0;
        zext_ln86_reg_587_pp0_iter1_reg[6 : 0] <= zext_ln86_reg_587[6 : 0];
    end
end

always @ (posedge ap_clk) begin
    if (((1'd1 == and_ln103_fu_307_p2) & (1'b1 == ap_CS_fsm_pp0_stage0) & (icmp_ln86_fu_285_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        lshr_ln_reg_614 <= {{ochan_reg_208[5:2]}};
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        quad_3_36_fu_118 <= quad_3_57_fu_467_p3;
        quad_3_39_fu_114 <= quad_3_58_fu_475_p3;
        quad_3_40_fu_122 <= quad_3_55_fu_451_p3;
        quad_3_41_fu_126 <= quad_3_52_fu_427_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        running_sums_3_load_reg_624 <= running_sums_3_q1;
    end
end

always @ (*) begin
    if ((icmp_ln86_fu_285_p2 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state2 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state2 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state25)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter22 == 1'b0) & (ap_enable_reg_pp0_iter21 == 1'b0) & (ap_enable_reg_pp0_iter20 == 1'b0) & (ap_enable_reg_pp0_iter19 == 1'b0) & (ap_enable_reg_pp0_iter18 == 1'b0) & (ap_enable_reg_pp0_iter17 == 1'b0) & (ap_enable_reg_pp0_iter16 == 1'b0) & (ap_enable_reg_pp0_iter15 == 1'b0) & (ap_enable_reg_pp0_iter14 == 1'b0) & (ap_enable_reg_pp0_iter13 == 1'b0) & (ap_enable_reg_pp0_iter12 == 1'b0) & (ap_enable_reg_pp0_iter11 == 1'b0) & (ap_enable_reg_pp0_iter10 == 1'b0) & (ap_enable_reg_pp0_iter9 == 1'b0) & (ap_enable_reg_pp0_iter8 == 1'b0) & (ap_enable_reg_pp0_iter7 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state25)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_01_blk_n = indices_01_empty_n;
    end else begin
        indices_01_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (write4_empty_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_01_read = 1'b1;
    end else begin
        indices_01_read = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_12_blk_n = indices_12_empty_n;
    end else begin
        indices_12_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (write4_empty_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_12_read = 1'b1;
    end else begin
        indices_12_read = 1'b0;
    end
end

always @ (*) begin
    if ((((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001)) | ((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001)) | ((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001)) | ((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
        l2_adjustments_ce0 = 1'b1;
    end else begin
        l2_adjustments_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        l2_partial_sums_ce0 = 1'b1;
    end else begin
        l2_partial_sums_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001)) | ((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
        out_data_ce1 = 1'b1;
    end else begin
        out_data_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'd1 == and_ln103_reg_610_pp0_iter20_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        out_data_we1 = 1'b1;
    end else begin
        out_data_we1 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        running_sums_3_ce0 = 1'b1;
    end else begin
        running_sums_3_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        running_sums_3_ce1 = 1'b1;
    end else begin
        running_sums_3_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        running_sums_3_we0 = 1'b1;
    end else begin
        running_sums_3_we0 = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        write4_blk_n = write4_empty_n;
    end else begin
        write4_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (write4_empty_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        write4_read = 1'b1;
    end else begin
        write4_read = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_start == 1'b0) | (write4_empty_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((~((ap_enable_reg_pp0_iter0 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0) & (icmp_ln86_fu_285_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone)) & ~((ap_enable_reg_pp0_iter22 == 1'b1) & (ap_enable_reg_pp0_iter21 == 1'b0) & (1'b0 == ap_block_pp0_stage0_subdone)))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0) & (icmp_ln86_fu_285_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone)) | ((ap_enable_reg_pp0_iter22 == 1'b1) & (ap_enable_reg_pp0_iter21 == 1'b0) & (1'b0 == ap_block_pp0_stage0_subdone)))) begin
                ap_NS_fsm = ap_ST_fsm_state25;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state25 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln109_fu_273_p2 = ((sub_ln109_cast_fu_265_p1) + (zext_ln109_8_fu_269_p1));

assign add_ln86_fu_279_p2 = (ochan_reg_208 + 7'd1);

assign and_ln103_fu_307_p2 = (write4_read_reg_567 & icmp_ln103_fu_301_p2);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state25 = ap_CS_fsm[32'd2];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (write4_empty_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1));
end

assign ap_block_state10_pp0_stage0_iter8 = ~(1'b1 == 1'b1);

assign ap_block_state11_pp0_stage0_iter9 = ~(1'b1 == 1'b1);

assign ap_block_state12_pp0_stage0_iter10 = ~(1'b1 == 1'b1);

assign ap_block_state13_pp0_stage0_iter11 = ~(1'b1 == 1'b1);

assign ap_block_state14_pp0_stage0_iter12 = ~(1'b1 == 1'b1);

assign ap_block_state15_pp0_stage0_iter13 = ~(1'b1 == 1'b1);

assign ap_block_state16_pp0_stage0_iter14 = ~(1'b1 == 1'b1);

assign ap_block_state17_pp0_stage0_iter15 = ~(1'b1 == 1'b1);

assign ap_block_state18_pp0_stage0_iter16 = ~(1'b1 == 1'b1);

assign ap_block_state19_pp0_stage0_iter17 = ~(1'b1 == 1'b1);

assign ap_block_state20_pp0_stage0_iter18 = ~(1'b1 == 1'b1);

assign ap_block_state21_pp0_stage0_iter19 = ~(1'b1 == 1'b1);

assign ap_block_state22_pp0_stage0_iter20 = ~(1'b1 == 1'b1);

assign ap_block_state23_pp0_stage0_iter21 = ~(1'b1 == 1'b1);

assign ap_block_state24_pp0_stage0_iter22 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter4 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage0_iter5 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage0_iter6 = ~(1'b1 == 1'b1);

assign ap_block_state9_pp0_stage0_iter7 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign bitcast_ln109_10_fu_518_p1 = quad_3_57_fu_467_p3;

assign bitcast_ln109_11_fu_522_p1 = quad_3_55_fu_451_p3;

assign bitcast_ln109_12_fu_526_p1 = quad_3_52_fu_427_p3;

assign bitcast_ln109_fu_514_p1 = quad_3_58_fu_475_p3;

assign data_V_fu_378_p1 = biased_reg_675;

assign grp_fu_223_p1 = tmp_105_i_i_reg_650_pp0_iter15_reg;

assign grp_fu_227_p1 = trunc_ln95_fu_329_p1;

assign grp_fu_231_p1 = tmp_104_i_i_reg_645_pp0_iter11_reg;

assign icmp_ln103_fu_301_p2 = ((trunc_ln99_fu_297_p1 == 2'd3) ? 1'b1 : 1'b0);

assign icmp_ln86_fu_285_p2 = ((ochan_reg_208 == 7'd64) ? 1'b1 : 1'b0);

assign icmp_ln99_7_fu_409_p2 = ((trunc_ln99_reg_603_pp0_iter20_reg == 2'd1) ? 1'b1 : 1'b0);

assign icmp_ln99_8_fu_422_p2 = ((trunc_ln99_reg_603_pp0_iter20_reg == 2'd0) ? 1'b1 : 1'b0);

assign icmp_ln99_fu_396_p2 = ((trunc_ln99_reg_603_pp0_iter20_reg == 2'd2) ? 1'b1 : 1'b0);

assign l2_adjustments_address0 = zext_ln86_reg_587_pp0_iter3_reg;

assign l2_partial_sums_address0 = zext_ln86_fu_291_p1;

assign out_data_address1 = sext_ln109_fu_509_p1;

assign out_data_d1 = {{{{bitcast_ln109_12_fu_526_p1}, {bitcast_ln109_11_fu_522_p1}}, {bitcast_ln109_10_fu_518_p1}}, {bitcast_ln109_fu_514_p1}};

assign p_Result_s_fu_381_p3 = data_V_fu_378_p1[32'd15];

assign quad_0_fu_389_p3 = ((p_Result_s_fu_381_p3[0:0] == 1'b1) ? 16'd0 : biased_reg_675);

assign quad_3_51_fu_414_p3 = ((icmp_ln99_7_fu_409_p2[0:0] == 1'b1) ? quad_3_41_fu_126 : quad_3_fu_401_p3);

assign quad_3_52_fu_427_p3 = ((icmp_ln99_8_fu_422_p2[0:0] == 1'b1) ? quad_3_41_fu_126 : quad_3_51_fu_414_p3);

assign quad_3_53_fu_435_p3 = ((icmp_ln99_fu_396_p2[0:0] == 1'b1) ? quad_0_fu_389_p3 : quad_3_40_fu_122);

assign quad_3_54_fu_443_p3 = ((icmp_ln99_7_fu_409_p2[0:0] == 1'b1) ? quad_3_40_fu_122 : quad_3_53_fu_435_p3);

assign quad_3_55_fu_451_p3 = ((icmp_ln99_8_fu_422_p2[0:0] == 1'b1) ? quad_3_40_fu_122 : quad_3_54_fu_443_p3);

assign quad_3_56_fu_459_p3 = ((icmp_ln99_7_fu_409_p2[0:0] == 1'b1) ? quad_0_fu_389_p3 : quad_3_36_fu_118);

assign quad_3_57_fu_467_p3 = ((icmp_ln99_8_fu_422_p2[0:0] == 1'b1) ? quad_3_36_fu_118 : quad_3_56_fu_459_p3);

assign quad_3_58_fu_475_p3 = ((icmp_ln99_8_fu_422_p2[0:0] == 1'b1) ? quad_0_fu_389_p3 : quad_3_39_fu_114);

assign quad_3_fu_401_p3 = ((icmp_ln99_fu_396_p2[0:0] == 1'b1) ? quad_3_41_fu_126 : quad_0_fu_389_p3);

assign running_sums_3_address1 = zext_ln86_fu_291_p1;

assign running_sums_3_d0 = ((write4_read_reg_567[0:0] == 1'b1) ? 16'd0 : sum_reg_634);

assign sext_ln109_fu_509_p1 = (tmp_74_fu_503_p3);

assign sub_ln109_cast_fu_265_p1 = (sub_ln109_fu_259_p2);

assign sub_ln109_fu_259_p2 = (zext_ln109_fu_243_p1 - zext_ln109_7_fu_255_p1);

assign tmp_74_fu_503_p3 = {{add_ln109_reg_573}, {lshr_ln_reg_614_pp0_iter20_reg}};

assign tmp_fu_235_p3 = {{indices_01_dout}, {4'd0}};

assign tmp_s_fu_247_p3 = {{indices_01_dout}, {1'd0}};

assign trunc_ln95_fu_329_p1 = l2_adjustments_q0[15:0];

assign trunc_ln99_fu_297_p1 = ochan_reg_208[1:0];

assign zext_ln109_7_fu_255_p1 = tmp_s_fu_247_p3;

assign zext_ln109_8_fu_269_p1 = indices_12_dout;

assign zext_ln109_fu_243_p1 = tmp_fu_235_p3;

assign zext_ln86_fu_291_p1 = ochan_reg_208;

always @ (posedge ap_clk) begin
    zext_ln86_reg_587[63:7] <= 57'b000000000000000000000000000000000000000000000000000000000;
    zext_ln86_reg_587_pp0_iter1_reg[63:7] <= 57'b000000000000000000000000000000000000000000000000000000000;
    zext_ln86_reg_587_pp0_iter2_reg[63:7] <= 57'b000000000000000000000000000000000000000000000000000000000;
    zext_ln86_reg_587_pp0_iter3_reg[63:7] <= 57'b000000000000000000000000000000000000000000000000000000000;
end

endmodule //td_fused_top_tdf10_l2_writeOutputs_165
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf10_readFilters68 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        filter_data_address0,
        filter_data_ce0,
        filter_data_q0,
        indices_23_dout,
        indices_23_empty_n,
        indices_23_read,
        weight_vecs_0_address0,
        weight_vecs_0_ce0,
        weight_vecs_0_we0,
        weight_vecs_0_d0,
        weight_vecs_0_address1,
        weight_vecs_0_ce1,
        weight_vecs_0_we1,
        weight_vecs_0_d1
);

parameter    ap_ST_fsm_state1 = 4'd1;
parameter    ap_ST_fsm_pp0_stage0 = 4'd2;
parameter    ap_ST_fsm_pp0_stage1 = 4'd4;
parameter    ap_ST_fsm_state7 = 4'd8;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [16:0] filter_data_address0;
output   filter_data_ce0;
input  [63:0] filter_data_q0;
input  [8:0] indices_23_dout;
input   indices_23_empty_n;
output   indices_23_read;
output  [9:0] weight_vecs_0_address0;
output   weight_vecs_0_ce0;
output   weight_vecs_0_we0;
output  [15:0] weight_vecs_0_d0;
output  [9:0] weight_vecs_0_address1;
output   weight_vecs_0_ce1;
output   weight_vecs_0_we1;
output  [15:0] weight_vecs_0_d1;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg filter_data_ce0;
reg indices_23_read;
reg[9:0] weight_vecs_0_address0;
reg weight_vecs_0_ce0;
reg weight_vecs_0_we0;
reg[15:0] weight_vecs_0_d0;
reg[9:0] weight_vecs_0_address1;
reg weight_vecs_0_ce1;
reg weight_vecs_0_we1;
reg[15:0] weight_vecs_0_d1;

reg    ap_done_reg;
  reg   [3:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    indices_23_blk_n;
reg   [7:0] indvar_flatten13_reg_174;
reg   [1:0] ii_reg_185;
reg   [6:0] indvar_flatten_reg_196;
reg   [1:0] jj_reg_207;
reg   [6:0] kk_0_i_i_reg_218;
wire   [12:0] sext_ln47_fu_251_p1;
reg   [12:0] sext_ln47_reg_583;
wire   [7:0] add_ln47_8_fu_255_p2;
reg   [7:0] add_ln47_8_reg_588;
wire    ap_CS_fsm_pp0_stage0;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state4_pp0_stage0_iter1;
wire    ap_block_state6_pp0_stage0_iter2;
wire    ap_block_pp0_stage0_11001;
wire   [0:0] icmp_ln47_fu_261_p2;
reg   [0:0] icmp_ln47_reg_593;
reg   [0:0] icmp_ln47_reg_593_pp0_iter1_reg;
wire   [0:0] icmp_ln48_fu_273_p2;
reg   [0:0] icmp_ln48_reg_597;
wire   [1:0] select_ln47_8_fu_287_p3;
reg   [1:0] select_ln47_8_reg_602;
wire   [6:0] select_ln48_fu_356_p3;
reg   [6:0] select_ln48_reg_609;
wire   [1:0] select_ln48_15_fu_364_p3;
reg   [1:0] select_ln48_15_reg_615;
wire   [5:0] empty_149_fu_382_p1;
reg   [5:0] empty_149_reg_621;
reg   [5:0] empty_149_reg_621_pp0_iter1_reg;
wire   [6:0] add_ln48_8_fu_405_p2;
reg   [6:0] add_ln48_8_reg_633;
wire   [6:0] add_ln49_fu_411_p2;
reg   [6:0] add_ln49_reg_638;
wire    ap_CS_fsm_pp0_stage1;
wire    ap_block_state3_pp0_stage1_iter0;
wire    ap_block_state5_pp0_stage1_iter1;
wire    ap_block_pp0_stage1_11001;
wire   [6:0] select_ln48_16_fu_416_p3;
reg   [6:0] select_ln48_16_reg_643;
wire   [5:0] add_ln55_29_fu_449_p2;
reg   [5:0] add_ln55_29_reg_648;
wire   [9:0] add_ln55_30_fu_470_p2;
reg   [9:0] add_ln55_30_reg_655;
reg   [15:0] tmp_102_i_i_reg_660;
reg   [15:0] tmp_103_i_i_reg_665;
reg    ap_block_state1;
wire    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_exit_iter0_state2;
reg    ap_enable_reg_pp0_iter1;
wire    ap_block_pp0_stage1_subdone;
reg    ap_enable_reg_pp0_iter2;
reg   [7:0] ap_phi_mux_indvar_flatten13_phi_fu_178_p4;
wire    ap_block_pp0_stage0;
reg   [1:0] ap_phi_mux_ii_phi_fu_189_p4;
reg   [6:0] ap_phi_mux_indvar_flatten_phi_fu_200_p4;
reg   [1:0] ap_phi_mux_jj_phi_fu_211_p4;
reg   [6:0] ap_phi_mux_kk_0_i_i_phi_fu_222_p4;
wire   [63:0] tmp_19_fu_396_p3;
wire   [63:0] zext_ln55_75_fu_476_p1;
wire    ap_block_pp0_stage1;
wire   [63:0] sext_ln55_7_fu_501_p1;
wire   [63:0] sext_ln55_8_fu_553_p1;
wire   [63:0] sext_ln55_9_fu_574_p1;
wire   [15:0] bitcast_ln55_fu_484_p1;
wire   [15:0] bitcast_ln55_4_fu_516_p1;
wire   [15:0] bitcast_ln55_5_fu_558_p1;
wire   [15:0] bitcast_ln55_6_fu_579_p1;
wire   [10:0] tmp_fu_233_p3;
wire   [11:0] zext_ln55_68_fu_241_p1;
wire   [11:0] zext_ln55_fu_229_p1;
wire   [11:0] sub_ln55_fu_245_p2;
wire   [1:0] add_ln47_fu_267_p2;
wire   [12:0] zext_ln55_70_fu_295_p1;
wire   [12:0] add_ln55_fu_299_p2;
wire   [14:0] tmp_69_fu_308_p3;
wire   [59:0] sext_ln55_6_fu_316_p1;
wire   [59:0] sext_ln55_fu_304_p1;
wire   [0:0] icmp_ln49_fu_332_p2;
wire   [0:0] xor_ln47_fu_326_p2;
wire   [1:0] select_ln47_fu_279_p3;
wire   [0:0] and_ln47_fu_338_p2;
wire   [0:0] or_ln48_fu_350_p2;
wire   [1:0] add_ln48_fu_344_p2;
wire   [59:0] sub_ln55_17_fu_320_p2;
wire   [59:0] zext_ln55_73_fu_372_p1;
wire   [59:0] add_ln55_28_fu_376_p2;
wire   [3:0] lshr_ln_fu_386_p4;
wire   [3:0] tmp_s_fu_425_p3;
wire   [4:0] zext_ln55_71_fu_432_p1;
wire   [4:0] zext_ln55_69_fu_422_p1;
wire   [4:0] sub_ln55_18_fu_436_p2;
wire   [5:0] sext_ln48_fu_442_p1;
wire   [5:0] zext_ln55_72_fu_446_p1;
wire   [3:0] trunc_ln55_fu_455_p1;
wire   [9:0] tmp_191_cast_fu_459_p3;
wire   [9:0] zext_ln55_74_fu_467_p1;
wire   [15:0] trunc_ln55_5_fu_480_p1;
wire   [5:0] or_ln49_fu_489_p2;
wire   [11:0] tmp_70_fu_494_p3;
wire   [15:0] tmp_101_i_i_fu_506_p4;
wire   [5:0] or_ln49_3_fu_541_p2;
wire   [11:0] tmp_71_fu_546_p3;
wire   [5:0] or_ln49_4_fu_562_p2;
wire   [11:0] tmp_72_fu_567_p3;
wire    ap_CS_fsm_state7;
reg   [3:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 4'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state7)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b1 == ap_condition_pp0_exit_iter0_state2))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1)) | ((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b0)))) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end else if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter2 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_reg_593 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ii_reg_185 <= select_ln47_8_reg_602;
    end else if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ii_reg_185 <= 2'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_reg_593 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        indvar_flatten13_reg_174 <= add_ln47_8_reg_588;
    end else if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indvar_flatten13_reg_174 <= 8'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_reg_593 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        indvar_flatten_reg_196 <= select_ln48_16_reg_643;
    end else if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indvar_flatten_reg_196 <= 7'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_reg_593 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        jj_reg_207 <= select_ln48_15_reg_615;
    end else if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        jj_reg_207 <= 2'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_reg_593 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        kk_0_i_i_reg_218 <= add_ln49_reg_638;
    end else if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        kk_0_i_i_reg_218 <= 7'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        add_ln47_8_reg_588 <= add_ln47_8_fu_255_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_fu_261_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        add_ln48_8_reg_633 <= add_ln48_8_fu_405_p2;
        empty_149_reg_621 <= empty_149_fu_382_p1;
        icmp_ln48_reg_597 <= icmp_ln48_fu_273_p2;
        select_ln48_reg_609 <= select_ln48_fu_356_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_reg_593 == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
        add_ln49_reg_638 <= add_ln49_fu_411_p2;
        select_ln48_16_reg_643 <= select_ln48_16_fu_416_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_reg_593 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        add_ln55_29_reg_648 <= add_ln55_29_fu_449_p2;
        add_ln55_30_reg_655 <= add_ln55_30_fu_470_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        empty_149_reg_621_pp0_iter1_reg <= empty_149_reg_621;
        icmp_ln47_reg_593 <= icmp_ln47_fu_261_p2;
        icmp_ln47_reg_593_pp0_iter1_reg <= icmp_ln47_reg_593;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_fu_261_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        select_ln47_8_reg_602 <= select_ln47_8_fu_287_p3;
        select_ln48_15_reg_615 <= select_ln48_15_fu_364_p3;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state1)) begin
        sext_ln47_reg_583 <= sext_ln47_fu_251_p1;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_reg_593_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
        tmp_102_i_i_reg_660 <= {{filter_data_q0[47:32]}};
        tmp_103_i_i_reg_665 <= {{filter_data_q0[63:48]}};
    end
end

always @ (*) begin
    if ((icmp_ln47_fu_261_p2 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state2 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state2 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state7)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln47_reg_593 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_ii_phi_fu_189_p4 = select_ln47_8_reg_602;
    end else begin
        ap_phi_mux_ii_phi_fu_189_p4 = ii_reg_185;
    end
end

always @ (*) begin
    if (((icmp_ln47_reg_593 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_indvar_flatten13_phi_fu_178_p4 = add_ln47_8_reg_588;
    end else begin
        ap_phi_mux_indvar_flatten13_phi_fu_178_p4 = indvar_flatten13_reg_174;
    end
end

always @ (*) begin
    if (((icmp_ln47_reg_593 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_indvar_flatten_phi_fu_200_p4 = select_ln48_16_reg_643;
    end else begin
        ap_phi_mux_indvar_flatten_phi_fu_200_p4 = indvar_flatten_reg_196;
    end
end

always @ (*) begin
    if (((icmp_ln47_reg_593 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_jj_phi_fu_211_p4 = select_ln48_15_reg_615;
    end else begin
        ap_phi_mux_jj_phi_fu_211_p4 = jj_reg_207;
    end
end

always @ (*) begin
    if (((icmp_ln47_reg_593 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_kk_0_i_i_phi_fu_222_p4 = add_ln49_reg_638;
    end else begin
        ap_phi_mux_kk_0_i_i_phi_fu_222_p4 = kk_0_i_i_reg_218;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state7)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1)) | ((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)) | ((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1)))) begin
        filter_data_ce0 = 1'b1;
    end else begin
        filter_data_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_23_blk_n = indices_23_empty_n;
    end else begin
        indices_23_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_23_read = 1'b1;
    end else begin
        indices_23_read = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        weight_vecs_0_address0 = sext_ln55_9_fu_574_p1;
    end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        weight_vecs_0_address0 = sext_ln55_7_fu_501_p1;
    end else begin
        weight_vecs_0_address0 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        weight_vecs_0_address1 = sext_ln55_8_fu_553_p1;
    end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        weight_vecs_0_address1 = zext_ln55_75_fu_476_p1;
    end else begin
        weight_vecs_0_address1 = 'bx;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1)) | ((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1)))) begin
        weight_vecs_0_ce0 = 1'b1;
    end else begin
        weight_vecs_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1)) | ((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1)))) begin
        weight_vecs_0_ce1 = 1'b1;
    end else begin
        weight_vecs_0_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        weight_vecs_0_d0 = bitcast_ln55_6_fu_579_p1;
    end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        weight_vecs_0_d0 = bitcast_ln55_4_fu_516_p1;
    end else begin
        weight_vecs_0_d0 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        weight_vecs_0_d1 = bitcast_ln55_5_fu_558_p1;
    end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        weight_vecs_0_d1 = bitcast_ln55_fu_484_p1;
    end else begin
        weight_vecs_0_d1 = 'bx;
    end
end

always @ (*) begin
    if ((((icmp_ln47_reg_593_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1)) | ((icmp_ln47_reg_593_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1)))) begin
        weight_vecs_0_we0 = 1'b1;
    end else begin
        weight_vecs_0_we0 = 1'b0;
    end
end

always @ (*) begin
    if ((((icmp_ln47_reg_593_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1)) | ((icmp_ln47_reg_593_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1)))) begin
        weight_vecs_0_we1 = 1'b1;
    end else begin
        weight_vecs_0_we1 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((~((icmp_ln47_fu_261_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0)) & ~((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0)) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end else if ((((icmp_ln47_fu_261_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0)) | ((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_state7;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_pp0_stage1 : begin
            if ((1'b0 == ap_block_pp0_stage1_subdone)) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end
        end
        ap_ST_fsm_state7 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln47_8_fu_255_p2 = (ap_phi_mux_indvar_flatten13_phi_fu_178_p4 + 8'd1);

assign add_ln47_fu_267_p2 = (ap_phi_mux_ii_phi_fu_189_p4 + 2'd1);

assign add_ln48_8_fu_405_p2 = (ap_phi_mux_indvar_flatten_phi_fu_200_p4 + 7'd1);

assign add_ln48_fu_344_p2 = (select_ln47_fu_279_p3 + 2'd1);

assign add_ln49_fu_411_p2 = (select_ln48_reg_609 + 7'd4);

assign add_ln55_28_fu_376_p2 = (sub_ln55_17_fu_320_p2 + zext_ln55_73_fu_372_p1);

assign add_ln55_29_fu_449_p2 = ((sext_ln48_fu_442_p1) + (zext_ln55_72_fu_446_p1));

assign add_ln55_30_fu_470_p2 = (tmp_191_cast_fu_459_p3 + zext_ln55_74_fu_467_p1);

assign add_ln55_fu_299_p2 = ((sext_ln47_reg_583) + (zext_ln55_70_fu_295_p1));

assign and_ln47_fu_338_p2 = (xor_ln47_fu_326_p2 & icmp_ln49_fu_332_p2);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_pp0_stage1 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state7 = ap_CS_fsm[32'd3];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1));
end

assign ap_block_state2_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage1_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage1_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign bitcast_ln55_4_fu_516_p1 = tmp_101_i_i_fu_506_p4;

assign bitcast_ln55_5_fu_558_p1 = tmp_102_i_i_reg_660;

assign bitcast_ln55_6_fu_579_p1 = tmp_103_i_i_reg_665;

assign bitcast_ln55_fu_484_p1 = trunc_ln55_5_fu_480_p1;

assign empty_149_fu_382_p1 = select_ln48_fu_356_p3[5:0];

assign filter_data_address0 = tmp_19_fu_396_p3;

assign icmp_ln47_fu_261_p2 = ((ap_phi_mux_indvar_flatten13_phi_fu_178_p4 == 8'd144) ? 1'b1 : 1'b0);

assign icmp_ln48_fu_273_p2 = ((ap_phi_mux_indvar_flatten_phi_fu_200_p4 == 7'd48) ? 1'b1 : 1'b0);

assign icmp_ln49_fu_332_p2 = ((ap_phi_mux_kk_0_i_i_phi_fu_222_p4 == 7'd64) ? 1'b1 : 1'b0);

assign lshr_ln_fu_386_p4 = {{select_ln48_fu_356_p3[5:2]}};

assign or_ln48_fu_350_p2 = (icmp_ln48_fu_273_p2 | and_ln47_fu_338_p2);

assign or_ln49_3_fu_541_p2 = (empty_149_reg_621_pp0_iter1_reg | 6'd2);

assign or_ln49_4_fu_562_p2 = (empty_149_reg_621_pp0_iter1_reg | 6'd3);

assign or_ln49_fu_489_p2 = (empty_149_reg_621_pp0_iter1_reg | 6'd1);

assign select_ln47_8_fu_287_p3 = ((icmp_ln48_fu_273_p2[0:0] == 1'b1) ? add_ln47_fu_267_p2 : ap_phi_mux_ii_phi_fu_189_p4);

assign select_ln47_fu_279_p3 = ((icmp_ln48_fu_273_p2[0:0] == 1'b1) ? 2'd0 : ap_phi_mux_jj_phi_fu_211_p4);

assign select_ln48_15_fu_364_p3 = ((and_ln47_fu_338_p2[0:0] == 1'b1) ? add_ln48_fu_344_p2 : select_ln47_fu_279_p3);

assign select_ln48_16_fu_416_p3 = ((icmp_ln48_reg_597[0:0] == 1'b1) ? 7'd1 : add_ln48_8_reg_633);

assign select_ln48_fu_356_p3 = ((or_ln48_fu_350_p2[0:0] == 1'b1) ? 7'd0 : ap_phi_mux_kk_0_i_i_phi_fu_222_p4);

assign sext_ln47_fu_251_p1 = (sub_ln55_fu_245_p2);

assign sext_ln48_fu_442_p1 = (sub_ln55_18_fu_436_p2);

assign sext_ln55_6_fu_316_p1 = (tmp_69_fu_308_p3);

assign sext_ln55_7_fu_501_p1 = (tmp_70_fu_494_p3);

assign sext_ln55_8_fu_553_p1 = (tmp_71_fu_546_p3);

assign sext_ln55_9_fu_574_p1 = (tmp_72_fu_567_p3);

assign sext_ln55_fu_304_p1 = add_ln55_fu_299_p2;

assign sub_ln55_17_fu_320_p2 = ((sext_ln55_6_fu_316_p1) - (sext_ln55_fu_304_p1));

assign sub_ln55_18_fu_436_p2 = (zext_ln55_71_fu_432_p1 - zext_ln55_69_fu_422_p1);

assign sub_ln55_fu_245_p2 = (zext_ln55_68_fu_241_p1 - zext_ln55_fu_229_p1);

assign tmp_101_i_i_fu_506_p4 = {{filter_data_q0[31:16]}};

assign tmp_191_cast_fu_459_p3 = {{trunc_ln55_fu_455_p1}, {6'd0}};

assign tmp_19_fu_396_p3 = {{add_ln55_28_fu_376_p2}, {lshr_ln_fu_386_p4}};

assign tmp_69_fu_308_p3 = {{add_ln55_fu_299_p2}, {2'd0}};

assign tmp_70_fu_494_p3 = {{add_ln55_29_reg_648}, {or_ln49_fu_489_p2}};

assign tmp_71_fu_546_p3 = {{add_ln55_29_reg_648}, {or_ln49_3_fu_541_p2}};

assign tmp_72_fu_567_p3 = {{add_ln55_29_reg_648}, {or_ln49_4_fu_562_p2}};

assign tmp_fu_233_p3 = {{indices_23_dout}, {2'd0}};

assign tmp_s_fu_425_p3 = {{select_ln47_8_reg_602}, {2'd0}};

assign trunc_ln55_5_fu_480_p1 = filter_data_q0[15:0];

assign trunc_ln55_fu_455_p1 = add_ln55_29_fu_449_p2[3:0];

assign xor_ln47_fu_326_p2 = (icmp_ln48_fu_273_p2 ^ 1'd1);

assign zext_ln55_68_fu_241_p1 = tmp_fu_233_p3;

assign zext_ln55_69_fu_422_p1 = select_ln47_8_reg_602;

assign zext_ln55_70_fu_295_p1 = select_ln47_8_fu_287_p3;

assign zext_ln55_71_fu_432_p1 = tmp_s_fu_425_p3;

assign zext_ln55_72_fu_446_p1 = select_ln48_15_reg_615;

assign zext_ln55_73_fu_372_p1 = select_ln48_15_fu_364_p3;

assign zext_ln55_74_fu_467_p1 = select_ln48_reg_609;

assign zext_ln55_75_fu_476_p1 = add_ln55_30_reg_655;

assign zext_ln55_fu_229_p1 = indices_23_dout;

endmodule //td_fused_top_tdf10_readFilters68
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf10_readInputs69 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        in_data_address0,
        in_data_ce0,
        in_data_q0,
        indices_01_dout,
        indices_01_empty_n,
        indices_01_read,
        indices_12_dout,
        indices_12_empty_n,
        indices_12_read,
        ifmap_vec_address0,
        ifmap_vec_ce0,
        ifmap_vec_we0,
        ifmap_vec_d0,
        ifmap_vec_address1,
        ifmap_vec_ce1,
        ifmap_vec_we1,
        ifmap_vec_d1,
        indices_01_out_din,
        indices_01_out_full_n,
        indices_01_out_write,
        indices_12_out_din,
        indices_12_out_full_n,
        indices_12_out_write
);

parameter    ap_ST_fsm_state1 = 5'd1;
parameter    ap_ST_fsm_state2 = 5'd2;
parameter    ap_ST_fsm_pp0_stage0 = 5'd4;
parameter    ap_ST_fsm_pp0_stage1 = 5'd8;
parameter    ap_ST_fsm_state9 = 5'd16;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [11:0] in_data_address0;
output   in_data_ce0;
input  [63:0] in_data_q0;
input  [15:0] indices_01_dout;
input   indices_01_empty_n;
output   indices_01_read;
input  [15:0] indices_12_dout;
input   indices_12_empty_n;
output   indices_12_read;
output  [9:0] ifmap_vec_address0;
output   ifmap_vec_ce0;
output   ifmap_vec_we0;
output  [15:0] ifmap_vec_d0;
output  [9:0] ifmap_vec_address1;
output   ifmap_vec_ce1;
output   ifmap_vec_we1;
output  [15:0] ifmap_vec_d1;
output  [3:0] indices_01_out_din;
input   indices_01_out_full_n;
output   indices_01_out_write;
output  [7:0] indices_12_out_din;
input   indices_12_out_full_n;
output   indices_12_out_write;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg in_data_ce0;
reg indices_01_read;
reg indices_12_read;
reg[9:0] ifmap_vec_address0;
reg ifmap_vec_ce0;
reg ifmap_vec_we0;
reg[15:0] ifmap_vec_d0;
reg[9:0] ifmap_vec_address1;
reg ifmap_vec_ce1;
reg ifmap_vec_we1;
reg[15:0] ifmap_vec_d1;
reg indices_01_out_write;
reg indices_12_out_write;

reg    ap_done_reg;
  reg   [4:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    indices_01_blk_n;
reg    indices_12_blk_n;
reg    indices_01_out_blk_n;
reg    indices_12_out_blk_n;
reg   [7:0] indvar_flatten47_reg_224;
reg   [1:0] ii_reg_236;
reg   [6:0] indvar_flatten_reg_248;
reg   [1:0] jj_reg_259;
reg   [6:0] kk_0_i_i_reg_271;
reg   [15:0] indices_01_read_reg_960;
wire   [3:0] trunc_ln250_fu_282_p1;
reg   [3:0] trunc_ln250_reg_965;
reg   [15:0] indices_12_read_reg_970;
wire   [7:0] empty_fu_287_p1;
reg   [7:0] empty_reg_975;
wire   [17:0] p_cast_i_i_fu_304_p1;
reg   [17:0] p_cast_i_i_reg_982;
wire    ap_CS_fsm_state2;
wire   [17:0] sext_ln22_fu_314_p1;
reg   [17:0] sext_ln22_reg_988;
wire   [3:0] p_cast_fu_318_p2;
reg   [3:0] p_cast_reg_994;
wire   [0:0] or_ln23_36_fu_337_p2;
reg   [0:0] or_ln23_36_reg_1000;
wire   [7:0] p_mid137_fu_343_p2;
reg   [7:0] p_mid137_reg_1005;
wire   [3:0] p_cast5_i_i_fu_361_p2;
reg   [3:0] p_cast5_i_i_reg_1010;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_block_state3_pp0_stage0_iter0;
wire    ap_block_state5_pp0_stage0_iter1;
wire    ap_block_state7_pp0_stage0_iter2;
wire    ap_block_pp0_stage0_11001;
wire   [0:0] is_padding_fu_401_p2;
reg   [0:0] is_padding_reg_1016;
wire   [0:0] icmp_ln19_fu_407_p2;
reg   [0:0] icmp_ln19_reg_1023;
reg   [0:0] icmp_ln19_reg_1023_pp0_iter1_reg;
reg   [0:0] icmp_ln19_reg_1023_pp0_iter2_reg;
wire   [1:0] add_ln19_fu_413_p2;
reg   [1:0] add_ln19_reg_1027;
wire   [0:0] icmp_ln20_fu_419_p2;
reg   [0:0] icmp_ln20_reg_1033;
wire   [1:0] select_ln19_fu_425_p3;
reg   [1:0] select_ln19_reg_1045;
wire   [0:0] or_ln23_38_fu_456_p2;
reg   [0:0] or_ln23_38_reg_1050;
wire   [1:0] add_ln20_fu_461_p2;
reg   [1:0] add_ln20_reg_1057;
wire   [0:0] or_ln23_40_fu_496_p2;
reg   [0:0] or_ln23_40_reg_1063;
wire   [6:0] add_ln20_8_fu_502_p2;
reg   [6:0] add_ln20_8_reg_1070;
wire   [7:0] add_ln19_8_fu_508_p2;
reg   [7:0] add_ln19_8_reg_1075;
wire    ap_CS_fsm_pp0_stage1;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_state4_pp0_stage1_iter0;
wire    ap_block_state6_pp0_stage1_iter1;
wire    ap_block_state8_pp0_stage1_iter2;
wire    ap_block_pp0_stage1_11001;
wire   [1:0] select_ln19_42_fu_546_p3;
reg   [1:0] select_ln19_42_reg_1080;
wire   [6:0] select_ln20_fu_620_p3;
reg   [6:0] select_ln20_reg_1087;
wire   [1:0] select_ln20_35_fu_628_p3;
reg   [1:0] select_ln20_35_reg_1093;
wire   [0:0] select_ln20_36_fu_637_p3;
reg   [0:0] select_ln20_36_reg_1099;
reg   [0:0] select_ln20_36_reg_1099_pp0_iter1_reg;
wire   [5:0] empty_148_fu_733_p1;
reg   [5:0] empty_148_reg_1107;
reg   [5:0] empty_148_reg_1107_pp0_iter1_reg;
wire   [6:0] select_ln20_39_fu_760_p3;
reg   [6:0] select_ln20_39_reg_1119;
wire   [6:0] add_ln25_fu_766_p2;
reg   [6:0] add_ln25_reg_1124;
reg    ap_enable_reg_pp0_iter1;
wire   [5:0] add_ln33_fu_798_p2;
reg   [5:0] add_ln33_reg_1129;
wire   [9:0] add_ln33_8_fu_819_p2;
reg   [9:0] add_ln33_8_reg_1136;
wire   [15:0] select_ln33_32_fu_898_p3;
reg   [15:0] select_ln33_32_reg_1141;
wire   [15:0] select_ln33_33_fu_919_p3;
reg   [15:0] select_ln33_33_reg_1146;
wire    ap_block_pp0_stage1_subdone;
reg    ap_condition_pp0_exit_iter0_state4;
reg    ap_enable_reg_pp0_iter2;
reg   [7:0] ap_phi_mux_indvar_flatten47_phi_fu_228_p4;
wire    ap_block_pp0_stage0;
reg   [1:0] ap_phi_mux_ii_phi_fu_240_p4;
reg   [6:0] ap_phi_mux_indvar_flatten_phi_fu_252_p4;
reg   [1:0] ap_phi_mux_jj_phi_fu_263_p4;
reg   [6:0] ap_phi_mux_kk_0_i_i_phi_fu_275_p4;
wire    ap_block_pp0_stage1;
wire   [63:0] sext_ln32_fu_755_p1;
wire   [63:0] zext_ln33_33_fu_825_p1;
wire   [63:0] sext_ln33_fu_857_p1;
wire   [63:0] sext_ln33_13_fu_938_p1;
wire   [63:0] sext_ln33_14_fu_955_p1;
reg    ap_block_state1;
wire   [15:0] select_ln33_fu_837_p3;
wire   [15:0] select_ln33_31_fu_876_p3;
wire   [16:0] zext_ln19_fu_295_p1;
wire   [16:0] empty_143_fu_298_p2;
wire   [16:0] j_cast_i_i_fu_292_p1;
wire   [16:0] add_ln22_fu_308_p2;
wire   [0:0] tmp_62_fu_323_p3;
wire   [0:0] icmp_ln24_fu_331_p2;
wire   [17:0] ii_cast_i_i_fu_348_p1;
wire   [3:0] ii_cast_fu_352_p1;
wire   [17:0] empty_144_fu_356_p2;
wire   [17:0] zext_ln20_fu_372_p1;
wire   [17:0] add_ln22_8_fu_376_p2;
wire   [0:0] tmp_63_fu_381_p3;
wire   [0:0] icmp_ln24_8_fu_389_p2;
wire   [0:0] or_ln23_fu_395_p2;
wire   [0:0] empty_145_fu_366_p2;
wire   [17:0] ii_cast_i_i_mid1_fu_433_p1;
wire   [17:0] p_mid111_fu_437_p2;
wire   [0:0] p_mid113_fu_442_p2;
wire   [17:0] zext_ln20_8_fu_467_p1;
wire   [17:0] add_ln22_9_fu_471_p2;
wire   [0:0] tmp_64_fu_476_p3;
wire   [0:0] icmp_ln24_9_fu_484_p2;
wire   [0:0] or_ln23_39_fu_490_p2;
wire   [0:0] select_ln19_44_fu_448_p3;
wire   [2:0] zext_ln22_fu_514_p1;
wire   [2:0] tmp1_fu_524_p2;
wire   [7:0] tmp1_cast_fu_530_p1;
wire   [7:0] empty_146_fu_534_p2;
wire   [3:0] ii_cast_mid1_fu_552_p1;
wire   [3:0] p_cast5_i_i_mid1_fu_555_p2;
wire   [3:0] row_coord_int_mid131_fu_571_p3;
wire   [3:0] row_coord_int_fu_518_p3;
wire   [7:0] col_coord_int_mid139_fu_578_p3;
wire   [7:0] col_coord_int_fu_539_p3;
wire   [0:0] icmp_ln25_fu_603_p2;
wire   [0:0] xor_ln19_fu_598_p2;
wire   [0:0] and_ln19_fu_609_p2;
wire   [0:0] or_ln20_fu_615_p2;
wire   [0:0] select_ln19_45_fu_566_p3;
wire   [3:0] select_ln19_43_fu_560_p3;
wire   [2:0] zext_ln22_8_fu_634_p1;
wire   [2:0] tmp1_mid1_fu_651_p2;
wire   [7:0] tmp1_cast_mid1_fu_657_p1;
wire   [7:0] p_mid1_fu_661_p2;
wire   [3:0] row_coord_int_mid1_fu_644_p3;
wire   [3:0] select_ln19_46_fu_584_p3;
wire   [3:0] select_ln20_37_fu_673_p3;
wire   [7:0] tmp_s_fu_681_p3;
wire   [4:0] tmp_18_fu_693_p3;
wire   [8:0] zext_ln32_fu_689_p1;
wire   [8:0] zext_ln32_36_fu_701_p1;
wire   [8:0] sub_ln32_fu_705_p2;
wire   [7:0] col_coord_int_mid1_fu_666_p3;
wire   [7:0] select_ln19_47_fu_591_p3;
wire   [7:0] select_ln20_38_fu_715_p3;
wire   [9:0] sext_ln20_fu_711_p1;
wire   [9:0] zext_ln32_37_fu_723_p1;
wire   [9:0] add_ln32_fu_727_p2;
wire   [3:0] lshr_ln_fu_737_p4;
wire   [13:0] tmp_65_fu_747_p3;
wire   [3:0] tmp_fu_774_p3;
wire   [4:0] zext_ln33_30_fu_781_p1;
wire   [4:0] zext_ln33_fu_771_p1;
wire   [4:0] sub_ln33_fu_785_p2;
wire   [5:0] sub_ln33_cast_fu_791_p1;
wire   [5:0] zext_ln33_31_fu_795_p1;
wire   [3:0] trunc_ln33_fu_804_p1;
wire   [9:0] tmp_180_cast_fu_808_p3;
wire   [9:0] zext_ln33_32_fu_816_p1;
wire   [15:0] trunc_ln32_fu_829_p1;
wire   [15:0] bitcast_ln32_fu_833_p1;
wire   [5:0] or_ln25_fu_845_p2;
wire   [11:0] tmp_66_fu_850_p3;
wire   [15:0] tmp_98_i_i_fu_862_p4;
wire   [15:0] bitcast_ln32_31_fu_872_p1;
wire   [15:0] tmp_99_i_i_fu_884_p4;
wire   [15:0] bitcast_ln32_32_fu_894_p1;
wire   [15:0] tmp_100_i_i_fu_905_p4;
wire   [15:0] bitcast_ln32_33_fu_915_p1;
wire   [5:0] or_ln25_21_fu_926_p2;
wire   [11:0] tmp_67_fu_931_p3;
wire   [5:0] or_ln25_22_fu_943_p2;
wire   [11:0] tmp_68_fu_948_p3;
wire    ap_CS_fsm_state9;
reg   [4:0] ap_NS_fsm;
wire    ap_block_pp0_stage0_subdone;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 5'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b1 == ap_condition_pp0_exit_iter0_state4) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_subdone))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_subdone))) begin
            if ((1'b1 == ap_condition_pp0_exit_iter0_state4)) begin
                ap_enable_reg_pp0_iter1 <= (1'b1 ^ ap_condition_pp0_exit_iter0_state4);
            end else if ((1'b1 == 1'b1)) begin
                ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
            end
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_subdone))) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            ap_enable_reg_pp0_iter2 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln19_reg_1023 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        ii_reg_236 <= select_ln19_42_reg_1080;
    end else if ((1'b1 == ap_CS_fsm_state2)) begin
        ii_reg_236 <= 2'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln19_reg_1023 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        indvar_flatten47_reg_224 <= add_ln19_8_reg_1075;
    end else if ((1'b1 == ap_CS_fsm_state2)) begin
        indvar_flatten47_reg_224 <= 8'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln19_reg_1023 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        indvar_flatten_reg_248 <= select_ln20_39_reg_1119;
    end else if ((1'b1 == ap_CS_fsm_state2)) begin
        indvar_flatten_reg_248 <= 7'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln19_reg_1023 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        jj_reg_259 <= select_ln20_35_reg_1093;
    end else if ((1'b1 == ap_CS_fsm_state2)) begin
        jj_reg_259 <= 2'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln19_reg_1023_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001))) begin
        kk_0_i_i_reg_271 <= add_ln25_reg_1124;
    end else if ((1'b1 == ap_CS_fsm_state2)) begin
        kk_0_i_i_reg_271 <= 7'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
        add_ln19_8_reg_1075 <= add_ln19_8_fu_508_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (icmp_ln19_fu_407_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        add_ln19_reg_1027 <= add_ln19_fu_413_p2;
        add_ln20_8_reg_1070 <= add_ln20_8_fu_502_p2;
        add_ln20_reg_1057 <= add_ln20_fu_461_p2;
        icmp_ln20_reg_1033 <= icmp_ln20_fu_419_p2;
        or_ln23_38_reg_1050 <= or_ln23_38_fu_456_p2;
        or_ln23_40_reg_1063 <= or_ln23_40_fu_496_p2;
        select_ln19_reg_1045 <= select_ln19_fu_425_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln19_reg_1023 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        add_ln25_reg_1124 <= add_ln25_fu_766_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln19_reg_1023_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001))) begin
        add_ln33_8_reg_1136 <= add_ln33_8_fu_819_p2;
        add_ln33_reg_1129 <= add_ln33_fu_798_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln19_reg_1023 == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001))) begin
        empty_148_reg_1107 <= empty_148_fu_733_p1;
        select_ln20_36_reg_1099 <= select_ln20_36_fu_637_p3;
        select_ln20_reg_1087 <= select_ln20_fu_620_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
        empty_148_reg_1107_pp0_iter1_reg <= empty_148_reg_1107;
        select_ln20_36_reg_1099_pp0_iter1_reg <= select_ln20_36_reg_1099;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state1)) begin
        empty_reg_975 <= empty_fu_287_p1;
        indices_01_read_reg_960 <= indices_01_dout;
        indices_12_read_reg_970 <= indices_12_dout;
        trunc_ln250_reg_965 <= trunc_ln250_fu_282_p1;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        icmp_ln19_reg_1023 <= icmp_ln19_fu_407_p2;
        icmp_ln19_reg_1023_pp0_iter1_reg <= icmp_ln19_reg_1023;
        icmp_ln19_reg_1023_pp0_iter2_reg <= icmp_ln19_reg_1023_pp0_iter1_reg;
        is_padding_reg_1016 <= is_padding_fu_401_p2;
        p_cast5_i_i_reg_1010 <= p_cast5_i_i_fu_361_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        or_ln23_36_reg_1000 <= or_ln23_36_fu_337_p2;
        p_cast_i_i_reg_982 <= p_cast_i_i_fu_304_p1;
        p_cast_reg_994 <= p_cast_fu_318_p2;
        p_mid137_reg_1005 <= p_mid137_fu_343_p2;
        sext_ln22_reg_988 <= sext_ln22_fu_314_p1;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln19_reg_1023 == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001))) begin
        select_ln19_42_reg_1080 <= select_ln19_42_fu_546_p3;
        select_ln20_35_reg_1093 <= select_ln20_35_fu_628_p3;
        select_ln20_39_reg_1119 <= select_ln20_39_fu_760_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (icmp_ln19_reg_1023_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        select_ln33_32_reg_1141 <= select_ln33_32_fu_898_p3;
        select_ln33_33_reg_1146 <= select_ln33_33_fu_919_p3;
    end
end

always @ (*) begin
    if ((icmp_ln19_reg_1023 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state4 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state4 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state9)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln19_reg_1023 == 1'd0) & (1'b0 == ap_block_pp0_stage0))) begin
        ap_phi_mux_ii_phi_fu_240_p4 = select_ln19_42_reg_1080;
    end else begin
        ap_phi_mux_ii_phi_fu_240_p4 = ii_reg_236;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln19_reg_1023 == 1'd0) & (1'b0 == ap_block_pp0_stage0))) begin
        ap_phi_mux_indvar_flatten47_phi_fu_228_p4 = add_ln19_8_reg_1075;
    end else begin
        ap_phi_mux_indvar_flatten47_phi_fu_228_p4 = indvar_flatten47_reg_224;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln19_reg_1023 == 1'd0) & (1'b0 == ap_block_pp0_stage0))) begin
        ap_phi_mux_indvar_flatten_phi_fu_252_p4 = select_ln20_39_reg_1119;
    end else begin
        ap_phi_mux_indvar_flatten_phi_fu_252_p4 = indvar_flatten_reg_248;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln19_reg_1023 == 1'd0) & (1'b0 == ap_block_pp0_stage0))) begin
        ap_phi_mux_jj_phi_fu_263_p4 = select_ln20_35_reg_1093;
    end else begin
        ap_phi_mux_jj_phi_fu_263_p4 = jj_reg_259;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln19_reg_1023_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage1))) begin
        ap_phi_mux_kk_0_i_i_phi_fu_275_p4 = add_ln25_reg_1124;
    end else begin
        ap_phi_mux_kk_0_i_i_phi_fu_275_p4 = kk_0_i_i_reg_271;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state9)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((ap_enable_reg_pp0_iter2 == 1'b1)) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ifmap_vec_address0 = sext_ln33_14_fu_955_p1;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0))) begin
            ifmap_vec_address0 = sext_ln33_fu_857_p1;
        end else begin
            ifmap_vec_address0 = 'bx;
        end
    end else begin
        ifmap_vec_address0 = 'bx;
    end
end

always @ (*) begin
    if ((ap_enable_reg_pp0_iter2 == 1'b1)) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ifmap_vec_address1 = sext_ln33_13_fu_938_p1;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0))) begin
            ifmap_vec_address1 = zext_ln33_33_fu_825_p1;
        end else begin
            ifmap_vec_address1 = 'bx;
        end
    end else begin
        ifmap_vec_address1 = 'bx;
    end
end

always @ (*) begin
    if ((((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_11001)) | ((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
        ifmap_vec_ce0 = 1'b1;
    end else begin
        ifmap_vec_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_11001)) | ((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
        ifmap_vec_ce1 = 1'b1;
    end else begin
        ifmap_vec_ce1 = 1'b0;
    end
end

always @ (*) begin
    if ((ap_enable_reg_pp0_iter2 == 1'b1)) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ifmap_vec_d0 = select_ln33_33_reg_1146;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0))) begin
            ifmap_vec_d0 = select_ln33_31_fu_876_p3;
        end else begin
            ifmap_vec_d0 = 'bx;
        end
    end else begin
        ifmap_vec_d0 = 'bx;
    end
end

always @ (*) begin
    if ((ap_enable_reg_pp0_iter2 == 1'b1)) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ifmap_vec_d1 = select_ln33_32_reg_1141;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0))) begin
            ifmap_vec_d1 = select_ln33_fu_837_p3;
        end else begin
            ifmap_vec_d1 = 'bx;
        end
    end else begin
        ifmap_vec_d1 = 'bx;
    end
end

always @ (*) begin
    if ((((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln19_reg_1023_pp0_iter2_reg == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001)) | ((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (icmp_ln19_reg_1023_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
        ifmap_vec_we0 = 1'b1;
    end else begin
        ifmap_vec_we0 = 1'b0;
    end
end

always @ (*) begin
    if ((((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln19_reg_1023_pp0_iter2_reg == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001)) | ((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (icmp_ln19_reg_1023_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
        ifmap_vec_we1 = 1'b1;
    end else begin
        ifmap_vec_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001)) | ((1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b0 == ap_block_pp0_stage1_11001)) | ((1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage1_11001)) | ((1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
        in_data_ce0 = 1'b1;
    end else begin
        in_data_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_01_blk_n = indices_01_empty_n;
    end else begin
        indices_01_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_01_out_blk_n = indices_01_out_full_n;
    end else begin
        indices_01_out_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((indices_12_out_full_n == 1'b0) | (indices_01_out_full_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_01_out_write = 1'b1;
    end else begin
        indices_01_out_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((indices_12_out_full_n == 1'b0) | (indices_01_out_full_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_01_read = 1'b1;
    end else begin
        indices_01_read = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_12_blk_n = indices_12_empty_n;
    end else begin
        indices_12_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_12_out_blk_n = indices_12_out_full_n;
    end else begin
        indices_12_out_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((indices_12_out_full_n == 1'b0) | (indices_01_out_full_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_12_out_write = 1'b1;
    end else begin
        indices_12_out_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((indices_12_out_full_n == 1'b0) | (indices_01_out_full_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_12_read = 1'b1;
    end else begin
        indices_12_read = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((indices_12_out_full_n == 1'b0) | (indices_01_out_full_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_state2 : begin
            ap_NS_fsm = ap_ST_fsm_pp0_stage0;
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_pp0_stage1 : begin
            if ((~((ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln19_reg_1023 == 1'd1) & (1'b0 == ap_block_pp0_stage1_subdone)) & ~((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b0) & (1'b0 == ap_block_pp0_stage1_subdone)) & (1'b0 == ap_block_pp0_stage1_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if ((((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b0) & (1'b0 == ap_block_pp0_stage1_subdone)) | ((ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln19_reg_1023 == 1'd1) & (1'b0 == ap_block_pp0_stage1_subdone)))) begin
                ap_NS_fsm = ap_ST_fsm_state9;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end
        end
        ap_ST_fsm_state9 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln19_8_fu_508_p2 = (indvar_flatten47_reg_224 + 8'd1);

assign add_ln19_fu_413_p2 = (ap_phi_mux_ii_phi_fu_240_p4 + 2'd1);

assign add_ln20_8_fu_502_p2 = (ap_phi_mux_indvar_flatten_phi_fu_252_p4 + 7'd1);

assign add_ln20_fu_461_p2 = (select_ln19_fu_425_p3 + 2'd1);

assign add_ln22_8_fu_376_p2 = ((sext_ln22_reg_988) + (zext_ln20_fu_372_p1));

assign add_ln22_9_fu_471_p2 = ((sext_ln22_reg_988) + (zext_ln20_8_fu_467_p1));

assign add_ln22_fu_308_p2 = ((j_cast_i_i_fu_292_p1) + (17'd131071));

assign add_ln25_fu_766_p2 = (select_ln20_reg_1087 + 7'd4);

assign add_ln32_fu_727_p2 = ((sext_ln20_fu_711_p1) + (zext_ln32_37_fu_723_p1));

assign add_ln33_8_fu_819_p2 = (tmp_180_cast_fu_808_p3 + zext_ln33_32_fu_816_p1);

assign add_ln33_fu_798_p2 = ((sub_ln33_cast_fu_791_p1) + (zext_ln33_31_fu_795_p1));

assign and_ln19_fu_609_p2 = (xor_ln19_fu_598_p2 & icmp_ln25_fu_603_p2);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_pp0_stage1 = ap_CS_fsm[32'd3];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state9 = ap_CS_fsm[32'd4];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((indices_12_out_full_n == 1'b0) | (indices_01_out_full_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0));
end

assign ap_block_state3_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage1_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage1_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage1_iter2 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign bitcast_ln32_31_fu_872_p1 = tmp_98_i_i_fu_862_p4;

assign bitcast_ln32_32_fu_894_p1 = tmp_99_i_i_fu_884_p4;

assign bitcast_ln32_33_fu_915_p1 = tmp_100_i_i_fu_905_p4;

assign bitcast_ln32_fu_833_p1 = trunc_ln32_fu_829_p1;

assign col_coord_int_fu_539_p3 = ((is_padding_reg_1016[0:0] == 1'b1) ? 8'd0 : empty_146_fu_534_p2);

assign col_coord_int_mid139_fu_578_p3 = ((or_ln23_38_reg_1050[0:0] == 1'b1) ? 8'd0 : p_mid137_reg_1005);

assign col_coord_int_mid1_fu_666_p3 = ((or_ln23_40_reg_1063[0:0] == 1'b1) ? 8'd0 : p_mid1_fu_661_p2);

assign empty_143_fu_298_p2 = ((zext_ln19_fu_295_p1) + (17'd131071));

assign empty_144_fu_356_p2 = ((p_cast_i_i_reg_982) + (ii_cast_i_i_fu_348_p1));

assign empty_145_fu_366_p2 = ((empty_144_fu_356_p2 > 18'd13) ? 1'b1 : 1'b0);

assign empty_146_fu_534_p2 = ((tmp1_cast_fu_530_p1) + (empty_reg_975));

assign empty_148_fu_733_p1 = select_ln20_fu_620_p3[5:0];

assign empty_fu_287_p1 = indices_12_dout[7:0];

assign icmp_ln19_fu_407_p2 = ((ap_phi_mux_indvar_flatten47_phi_fu_228_p4 == 8'd144) ? 1'b1 : 1'b0);

assign icmp_ln20_fu_419_p2 = ((ap_phi_mux_indvar_flatten_phi_fu_252_p4 == 7'd48) ? 1'b1 : 1'b0);

assign icmp_ln24_8_fu_389_p2 = (((add_ln22_8_fu_376_p2) > (18'd13)) ? 1'b1 : 1'b0);

assign icmp_ln24_9_fu_484_p2 = (((add_ln22_9_fu_471_p2) > (18'd13)) ? 1'b1 : 1'b0);

assign icmp_ln24_fu_331_p2 = (((add_ln22_fu_308_p2) > (17'd13)) ? 1'b1 : 1'b0);

assign icmp_ln25_fu_603_p2 = ((ap_phi_mux_kk_0_i_i_phi_fu_275_p4 == 7'd64) ? 1'b1 : 1'b0);

assign ii_cast_fu_352_p1 = ap_phi_mux_ii_phi_fu_240_p4;

assign ii_cast_i_i_fu_348_p1 = ap_phi_mux_ii_phi_fu_240_p4;

assign ii_cast_i_i_mid1_fu_433_p1 = add_ln19_fu_413_p2;

assign ii_cast_mid1_fu_552_p1 = add_ln19_reg_1027;

assign in_data_address0 = sext_ln32_fu_755_p1;

assign indices_01_out_din = indices_01_dout[3:0];

assign indices_12_out_din = indices_12_dout[7:0];

assign is_padding_fu_401_p2 = (or_ln23_fu_395_p2 | empty_145_fu_366_p2);

assign j_cast_i_i_fu_292_p1 = indices_12_read_reg_970;

assign lshr_ln_fu_737_p4 = {{select_ln20_fu_620_p3[5:2]}};

assign or_ln20_fu_615_p2 = (icmp_ln20_reg_1033 | and_ln19_fu_609_p2);

assign or_ln23_36_fu_337_p2 = (tmp_62_fu_323_p3 | icmp_ln24_fu_331_p2);

assign or_ln23_38_fu_456_p2 = (p_mid113_fu_442_p2 | or_ln23_36_reg_1000);

assign or_ln23_39_fu_490_p2 = (tmp_64_fu_476_p3 | icmp_ln24_9_fu_484_p2);

assign or_ln23_40_fu_496_p2 = (select_ln19_44_fu_448_p3 | or_ln23_39_fu_490_p2);

assign or_ln23_fu_395_p2 = (tmp_63_fu_381_p3 | icmp_ln24_8_fu_389_p2);

assign or_ln25_21_fu_926_p2 = (empty_148_reg_1107_pp0_iter1_reg | 6'd2);

assign or_ln25_22_fu_943_p2 = (empty_148_reg_1107_pp0_iter1_reg | 6'd3);

assign or_ln25_fu_845_p2 = (empty_148_reg_1107_pp0_iter1_reg | 6'd1);

assign p_cast5_i_i_fu_361_p2 = (p_cast_reg_994 + ii_cast_fu_352_p1);

assign p_cast5_i_i_mid1_fu_555_p2 = (p_cast_reg_994 + ii_cast_mid1_fu_552_p1);

assign p_cast_fu_318_p2 = ((trunc_ln250_reg_965) + (4'd15));

assign p_cast_i_i_fu_304_p1 = (empty_143_fu_298_p2);

assign p_mid111_fu_437_p2 = ((p_cast_i_i_reg_982) + (ii_cast_i_i_mid1_fu_433_p1));

assign p_mid113_fu_442_p2 = ((p_mid111_fu_437_p2 > 18'd13) ? 1'b1 : 1'b0);

assign p_mid137_fu_343_p2 = ((empty_reg_975) + (8'd255));

assign p_mid1_fu_661_p2 = ((tmp1_cast_mid1_fu_657_p1) + (empty_reg_975));

assign row_coord_int_fu_518_p3 = ((is_padding_reg_1016[0:0] == 1'b1) ? 4'd0 : p_cast5_i_i_reg_1010);

assign row_coord_int_mid131_fu_571_p3 = ((or_ln23_38_reg_1050[0:0] == 1'b1) ? 4'd0 : p_cast5_i_i_mid1_fu_555_p2);

assign row_coord_int_mid1_fu_644_p3 = ((or_ln23_40_reg_1063[0:0] == 1'b1) ? 4'd0 : select_ln19_43_fu_560_p3);

assign select_ln19_42_fu_546_p3 = ((icmp_ln20_reg_1033[0:0] == 1'b1) ? add_ln19_reg_1027 : ii_reg_236);

assign select_ln19_43_fu_560_p3 = ((icmp_ln20_reg_1033[0:0] == 1'b1) ? p_cast5_i_i_mid1_fu_555_p2 : p_cast5_i_i_reg_1010);

assign select_ln19_44_fu_448_p3 = ((icmp_ln20_fu_419_p2[0:0] == 1'b1) ? p_mid113_fu_442_p2 : empty_145_fu_366_p2);

assign select_ln19_45_fu_566_p3 = ((icmp_ln20_reg_1033[0:0] == 1'b1) ? or_ln23_38_reg_1050 : is_padding_reg_1016);

assign select_ln19_46_fu_584_p3 = ((icmp_ln20_reg_1033[0:0] == 1'b1) ? row_coord_int_mid131_fu_571_p3 : row_coord_int_fu_518_p3);

assign select_ln19_47_fu_591_p3 = ((icmp_ln20_reg_1033[0:0] == 1'b1) ? col_coord_int_mid139_fu_578_p3 : col_coord_int_fu_539_p3);

assign select_ln19_fu_425_p3 = ((icmp_ln20_fu_419_p2[0:0] == 1'b1) ? 2'd0 : ap_phi_mux_jj_phi_fu_263_p4);

assign select_ln20_35_fu_628_p3 = ((and_ln19_fu_609_p2[0:0] == 1'b1) ? add_ln20_reg_1057 : select_ln19_reg_1045);

assign select_ln20_36_fu_637_p3 = ((and_ln19_fu_609_p2[0:0] == 1'b1) ? or_ln23_40_reg_1063 : select_ln19_45_fu_566_p3);

assign select_ln20_37_fu_673_p3 = ((and_ln19_fu_609_p2[0:0] == 1'b1) ? row_coord_int_mid1_fu_644_p3 : select_ln19_46_fu_584_p3);

assign select_ln20_38_fu_715_p3 = ((and_ln19_fu_609_p2[0:0] == 1'b1) ? col_coord_int_mid1_fu_666_p3 : select_ln19_47_fu_591_p3);

assign select_ln20_39_fu_760_p3 = ((icmp_ln20_reg_1033[0:0] == 1'b1) ? 7'd1 : add_ln20_8_reg_1070);

assign select_ln20_fu_620_p3 = ((or_ln20_fu_615_p2[0:0] == 1'b1) ? 7'd0 : ap_phi_mux_kk_0_i_i_phi_fu_275_p4);

assign select_ln33_31_fu_876_p3 = ((select_ln20_36_reg_1099_pp0_iter1_reg[0:0] == 1'b1) ? 16'd0 : bitcast_ln32_31_fu_872_p1);

assign select_ln33_32_fu_898_p3 = ((select_ln20_36_reg_1099_pp0_iter1_reg[0:0] == 1'b1) ? 16'd0 : bitcast_ln32_32_fu_894_p1);

assign select_ln33_33_fu_919_p3 = ((select_ln20_36_reg_1099_pp0_iter1_reg[0:0] == 1'b1) ? 16'd0 : bitcast_ln32_33_fu_915_p1);

assign select_ln33_fu_837_p3 = ((select_ln20_36_reg_1099_pp0_iter1_reg[0:0] == 1'b1) ? 16'd0 : bitcast_ln32_fu_833_p1);

assign sext_ln20_fu_711_p1 = (sub_ln32_fu_705_p2);

assign sext_ln22_fu_314_p1 = add_ln22_fu_308_p2;

assign sext_ln32_fu_755_p1 = (tmp_65_fu_747_p3);

assign sext_ln33_13_fu_938_p1 = (tmp_67_fu_931_p3);

assign sext_ln33_14_fu_955_p1 = (tmp_68_fu_948_p3);

assign sext_ln33_fu_857_p1 = (tmp_66_fu_850_p3);

assign sub_ln32_fu_705_p2 = (zext_ln32_fu_689_p1 - zext_ln32_36_fu_701_p1);

assign sub_ln33_cast_fu_791_p1 = (sub_ln33_fu_785_p2);

assign sub_ln33_fu_785_p2 = (zext_ln33_30_fu_781_p1 - zext_ln33_fu_771_p1);

assign tmp1_cast_fu_530_p1 = (tmp1_fu_524_p2);

assign tmp1_cast_mid1_fu_657_p1 = (tmp1_mid1_fu_651_p2);

assign tmp1_fu_524_p2 = ((zext_ln22_fu_514_p1) + (3'd7));

assign tmp1_mid1_fu_651_p2 = ((zext_ln22_8_fu_634_p1) + (3'd7));

assign tmp_100_i_i_fu_905_p4 = {{in_data_q0[63:48]}};

assign tmp_180_cast_fu_808_p3 = {{trunc_ln33_fu_804_p1}, {6'd0}};

assign tmp_18_fu_693_p3 = {{select_ln20_37_fu_673_p3}, {1'd0}};

assign tmp_62_fu_323_p3 = add_ln22_fu_308_p2[32'd16];

assign tmp_63_fu_381_p3 = add_ln22_8_fu_376_p2[32'd17];

assign tmp_64_fu_476_p3 = add_ln22_9_fu_471_p2[32'd17];

assign tmp_65_fu_747_p3 = {{add_ln32_fu_727_p2}, {lshr_ln_fu_737_p4}};

assign tmp_66_fu_850_p3 = {{add_ln33_reg_1129}, {or_ln25_fu_845_p2}};

assign tmp_67_fu_931_p3 = {{add_ln33_reg_1129}, {or_ln25_21_fu_926_p2}};

assign tmp_68_fu_948_p3 = {{add_ln33_reg_1129}, {or_ln25_22_fu_943_p2}};

assign tmp_98_i_i_fu_862_p4 = {{in_data_q0[31:16]}};

assign tmp_99_i_i_fu_884_p4 = {{in_data_q0[47:32]}};

assign tmp_fu_774_p3 = {{select_ln19_42_reg_1080}, {2'd0}};

assign tmp_s_fu_681_p3 = {{select_ln20_37_fu_673_p3}, {4'd0}};

assign trunc_ln250_fu_282_p1 = indices_01_dout[3:0];

assign trunc_ln32_fu_829_p1 = in_data_q0[15:0];

assign trunc_ln33_fu_804_p1 = add_ln33_fu_798_p2[3:0];

assign xor_ln19_fu_598_p2 = (icmp_ln20_reg_1033 ^ 1'd1);

assign zext_ln19_fu_295_p1 = indices_01_read_reg_960;

assign zext_ln20_8_fu_467_p1 = add_ln20_fu_461_p2;

assign zext_ln20_fu_372_p1 = ap_phi_mux_jj_phi_fu_263_p4;

assign zext_ln22_8_fu_634_p1 = add_ln20_reg_1057;

assign zext_ln22_fu_514_p1 = jj_reg_259;

assign zext_ln32_36_fu_701_p1 = tmp_18_fu_693_p3;

assign zext_ln32_37_fu_723_p1 = select_ln20_38_fu_715_p3;

assign zext_ln32_fu_689_p1 = tmp_s_fu_681_p3;

assign zext_ln33_30_fu_781_p1 = tmp_fu_774_p3;

assign zext_ln33_31_fu_795_p1 = select_ln20_35_reg_1093;

assign zext_ln33_32_fu_816_p1 = select_ln20_reg_1087;

assign zext_ln33_33_fu_825_p1 = add_ln33_8_reg_1136;

assign zext_ln33_fu_771_p1 = select_ln19_42_reg_1080;

endmodule //td_fused_top_tdf10_readInputs69
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf1_114 (
        in_data_address0,
        in_data_ce0,
        in_data_d0,
        in_data_q0,
        in_data_we0,
        in_data_address1,
        in_data_ce1,
        in_data_d1,
        in_data_q1,
        in_data_we1,
        out_data_address0,
        out_data_ce0,
        out_data_d0,
        out_data_q0,
        out_data_we0,
        out_data_address1,
        out_data_ce1,
        out_data_d1,
        out_data_q1,
        out_data_we1,
        filter_data_address0,
        filter_data_ce0,
        filter_data_d0,
        filter_data_q0,
        filter_data_we0,
        filter_data_address1,
        filter_data_ce1,
        filter_data_d1,
        filter_data_q1,
        filter_data_we1,
        adjustments_address0,
        adjustments_ce0,
        adjustments_d0,
        adjustments_q0,
        adjustments_we0,
        adjustments_address1,
        adjustments_ce1,
        adjustments_d1,
        adjustments_q1,
        adjustments_we1,
        ap_clk,
        ap_rst,
        in_data_empty_n,
        in_data_read,
        out_data_full_n,
        out_data_write,
        ap_start,
        ap_done,
        ap_ready,
        ap_idle,
        ap_continue
);


output  [15:0] in_data_address0;
output   in_data_ce0;
output  [63:0] in_data_d0;
input  [63:0] in_data_q0;
output   in_data_we0;
output  [15:0] in_data_address1;
output   in_data_ce1;
output  [63:0] in_data_d1;
input  [63:0] in_data_q1;
output   in_data_we1;
output  [15:0] out_data_address0;
output   out_data_ce0;
output  [63:0] out_data_d0;
input  [63:0] out_data_q0;
output   out_data_we0;
output  [15:0] out_data_address1;
output   out_data_ce1;
output  [63:0] out_data_d1;
input  [63:0] out_data_q1;
output   out_data_we1;
output  [8:0] filter_data_address0;
output   filter_data_ce0;
output  [15:0] filter_data_d0;
input  [15:0] filter_data_q0;
output   filter_data_we0;
output  [8:0] filter_data_address1;
output   filter_data_ce1;
output  [15:0] filter_data_d1;
input  [15:0] filter_data_q1;
output   filter_data_we1;
output  [3:0] adjustments_address0;
output   adjustments_ce0;
output  [47:0] adjustments_d0;
input  [47:0] adjustments_q0;
output   adjustments_we0;
output  [3:0] adjustments_address1;
output   adjustments_ce1;
output  [47:0] adjustments_d1;
input  [47:0] adjustments_q1;
output   adjustments_we1;
input   ap_clk;
input   ap_rst;
input   in_data_empty_n;
output   in_data_read;
input   out_data_full_n;
output   out_data_write;
input   ap_start;
output   ap_done;
output   ap_ready;
output   ap_idle;
input   ap_continue;

reg ap_done;
reg ap_ready;
reg ap_idle;

wire   [15:0] dataflow_in_loop_TOP_LOOP38116_U0_in_data_address0;
wire    dataflow_in_loop_TOP_LOOP38116_U0_in_data_ce0;
wire   [63:0] dataflow_in_loop_TOP_LOOP38116_U0_in_data_d0;
wire    dataflow_in_loop_TOP_LOOP38116_U0_in_data_we0;
wire   [15:0] dataflow_in_loop_TOP_LOOP38116_U0_in_data_address1;
wire    dataflow_in_loop_TOP_LOOP38116_U0_in_data_ce1;
wire   [63:0] dataflow_in_loop_TOP_LOOP38116_U0_in_data_d1;
wire    dataflow_in_loop_TOP_LOOP38116_U0_in_data_we1;
wire   [8:0] dataflow_in_loop_TOP_LOOP38116_U0_filter_data_address0;
wire    dataflow_in_loop_TOP_LOOP38116_U0_filter_data_ce0;
wire   [15:0] dataflow_in_loop_TOP_LOOP38116_U0_filter_data_d0;
wire    dataflow_in_loop_TOP_LOOP38116_U0_filter_data_we0;
wire   [8:0] dataflow_in_loop_TOP_LOOP38116_U0_filter_data_address1;
wire    dataflow_in_loop_TOP_LOOP38116_U0_filter_data_ce1;
wire   [15:0] dataflow_in_loop_TOP_LOOP38116_U0_filter_data_d1;
wire    dataflow_in_loop_TOP_LOOP38116_U0_filter_data_we1;
wire   [3:0] dataflow_in_loop_TOP_LOOP38116_U0_adjustments_address0;
wire    dataflow_in_loop_TOP_LOOP38116_U0_adjustments_ce0;
wire   [47:0] dataflow_in_loop_TOP_LOOP38116_U0_adjustments_d0;
wire    dataflow_in_loop_TOP_LOOP38116_U0_adjustments_we0;
wire   [3:0] dataflow_in_loop_TOP_LOOP38116_U0_adjustments_address1;
wire    dataflow_in_loop_TOP_LOOP38116_U0_adjustments_ce1;
wire   [47:0] dataflow_in_loop_TOP_LOOP38116_U0_adjustments_d1;
wire    dataflow_in_loop_TOP_LOOP38116_U0_adjustments_we1;
wire   [15:0] dataflow_in_loop_TOP_LOOP38116_U0_out_data_address0;
wire    dataflow_in_loop_TOP_LOOP38116_U0_out_data_ce0;
wire   [63:0] dataflow_in_loop_TOP_LOOP38116_U0_out_data_d0;
wire    dataflow_in_loop_TOP_LOOP38116_U0_out_data_we0;
wire   [15:0] dataflow_in_loop_TOP_LOOP38116_U0_out_data_address1;
wire    dataflow_in_loop_TOP_LOOP38116_U0_out_data_ce1;
wire   [63:0] dataflow_in_loop_TOP_LOOP38116_U0_out_data_d1;
wire    dataflow_in_loop_TOP_LOOP38116_U0_out_data_we1;
wire    dataflow_in_loop_TOP_LOOP38116_U0_ap_start;
wire    dataflow_in_loop_TOP_LOOP38116_U0_in_data_read;
wire    dataflow_in_loop_TOP_LOOP38116_U0_out_data_write;
wire    dataflow_in_loop_TOP_LOOP38116_U0_ap_done;
wire    dataflow_in_loop_TOP_LOOP38116_U0_ap_ready;
wire    dataflow_in_loop_TOP_LOOP38116_U0_ap_idle;
reg    dataflow_in_loop_TOP_LOOP38116_U0_ap_continue;
wire    dataflow_in_loop_TOP_LOOP38116_U0_in_data_full_n;
wire    dataflow_in_loop_TOP_LOOP38116_U0_in_data_write;
wire    ap_sync_continue;
wire    ap_sync_done;
wire    ap_sync_ready;
reg   [19:0] loop_dataflow_input_count;
reg   [19:0] loop_dataflow_output_count;
wire   [19:0] bound_minus_1;
wire    dataflow_in_loop_TOP_LOOP38116_U0_start_full_n;
wire    dataflow_in_loop_TOP_LOOP38116_U0_start_write;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 loop_dataflow_input_count = 20'd0;
#0 loop_dataflow_output_count = 20'd0;
end

td_fused_top_dataflow_in_loop_TOP_LOOP38116 dataflow_in_loop_TOP_LOOP38116_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .in_data_address0(dataflow_in_loop_TOP_LOOP38116_U0_in_data_address0),
    .in_data_ce0(dataflow_in_loop_TOP_LOOP38116_U0_in_data_ce0),
    .in_data_d0(dataflow_in_loop_TOP_LOOP38116_U0_in_data_d0),
    .in_data_q0(in_data_q0),
    .in_data_we0(dataflow_in_loop_TOP_LOOP38116_U0_in_data_we0),
    .in_data_address1(dataflow_in_loop_TOP_LOOP38116_U0_in_data_address1),
    .in_data_ce1(dataflow_in_loop_TOP_LOOP38116_U0_in_data_ce1),
    .in_data_d1(dataflow_in_loop_TOP_LOOP38116_U0_in_data_d1),
    .in_data_q1(64'd0),
    .in_data_we1(dataflow_in_loop_TOP_LOOP38116_U0_in_data_we1),
    .filter_data_address0(dataflow_in_loop_TOP_LOOP38116_U0_filter_data_address0),
    .filter_data_ce0(dataflow_in_loop_TOP_LOOP38116_U0_filter_data_ce0),
    .filter_data_d0(dataflow_in_loop_TOP_LOOP38116_U0_filter_data_d0),
    .filter_data_q0(filter_data_q0),
    .filter_data_we0(dataflow_in_loop_TOP_LOOP38116_U0_filter_data_we0),
    .filter_data_address1(dataflow_in_loop_TOP_LOOP38116_U0_filter_data_address1),
    .filter_data_ce1(dataflow_in_loop_TOP_LOOP38116_U0_filter_data_ce1),
    .filter_data_d1(dataflow_in_loop_TOP_LOOP38116_U0_filter_data_d1),
    .filter_data_q1(16'd0),
    .filter_data_we1(dataflow_in_loop_TOP_LOOP38116_U0_filter_data_we1),
    .adjustments_address0(dataflow_in_loop_TOP_LOOP38116_U0_adjustments_address0),
    .adjustments_ce0(dataflow_in_loop_TOP_LOOP38116_U0_adjustments_ce0),
    .adjustments_d0(dataflow_in_loop_TOP_LOOP38116_U0_adjustments_d0),
    .adjustments_q0(adjustments_q0),
    .adjustments_we0(dataflow_in_loop_TOP_LOOP38116_U0_adjustments_we0),
    .adjustments_address1(dataflow_in_loop_TOP_LOOP38116_U0_adjustments_address1),
    .adjustments_ce1(dataflow_in_loop_TOP_LOOP38116_U0_adjustments_ce1),
    .adjustments_d1(dataflow_in_loop_TOP_LOOP38116_U0_adjustments_d1),
    .adjustments_q1(48'd0),
    .adjustments_we1(dataflow_in_loop_TOP_LOOP38116_U0_adjustments_we1),
    .out_data_address0(dataflow_in_loop_TOP_LOOP38116_U0_out_data_address0),
    .out_data_ce0(dataflow_in_loop_TOP_LOOP38116_U0_out_data_ce0),
    .out_data_d0(dataflow_in_loop_TOP_LOOP38116_U0_out_data_d0),
    .out_data_q0(64'd0),
    .out_data_we0(dataflow_in_loop_TOP_LOOP38116_U0_out_data_we0),
    .out_data_address1(dataflow_in_loop_TOP_LOOP38116_U0_out_data_address1),
    .out_data_ce1(dataflow_in_loop_TOP_LOOP38116_U0_out_data_ce1),
    .out_data_d1(dataflow_in_loop_TOP_LOOP38116_U0_out_data_d1),
    .out_data_q1(64'd0),
    .out_data_we1(dataflow_in_loop_TOP_LOOP38116_U0_out_data_we1),
    .ap_start(dataflow_in_loop_TOP_LOOP38116_U0_ap_start),
    .in_data_empty_n(1'b0),
    .in_data_read(dataflow_in_loop_TOP_LOOP38116_U0_in_data_read),
    .out_data_full_n(out_data_full_n),
    .out_data_write(dataflow_in_loop_TOP_LOOP38116_U0_out_data_write),
    .ap_done(dataflow_in_loop_TOP_LOOP38116_U0_ap_done),
    .ap_ready(dataflow_in_loop_TOP_LOOP38116_U0_ap_ready),
    .ap_idle(dataflow_in_loop_TOP_LOOP38116_U0_ap_idle),
    .ap_continue(dataflow_in_loop_TOP_LOOP38116_U0_ap_continue)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        loop_dataflow_input_count <= 20'd0;
    end else begin
        if ((~(loop_dataflow_input_count == bound_minus_1) & (dataflow_in_loop_TOP_LOOP38116_U0_ap_ready == 1'b1) & (ap_start == 1'b1))) begin
            loop_dataflow_input_count <= (loop_dataflow_input_count + 20'd1);
        end else if (((dataflow_in_loop_TOP_LOOP38116_U0_ap_ready == 1'b1) & (loop_dataflow_input_count == bound_minus_1) & (ap_start == 1'b1))) begin
            loop_dataflow_input_count <= 20'd0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        loop_dataflow_output_count <= 20'd0;
    end else begin
        if ((~(loop_dataflow_output_count == bound_minus_1) & (dataflow_in_loop_TOP_LOOP38116_U0_ap_continue == 1'b1) & (dataflow_in_loop_TOP_LOOP38116_U0_ap_done == 1'b1))) begin
            loop_dataflow_output_count <= (loop_dataflow_output_count + 20'd1);
        end else if (((dataflow_in_loop_TOP_LOOP38116_U0_ap_continue == 1'b1) & (dataflow_in_loop_TOP_LOOP38116_U0_ap_done == 1'b1) & (loop_dataflow_output_count == bound_minus_1))) begin
            loop_dataflow_output_count <= 20'd0;
        end
    end
end

always @ (*) begin
    if (((dataflow_in_loop_TOP_LOOP38116_U0_ap_done == 1'b1) & (loop_dataflow_output_count == bound_minus_1))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = 1'b0;
    end
end

always @ (*) begin
    if (((dataflow_in_loop_TOP_LOOP38116_U0_ap_idle == 1'b1) & (loop_dataflow_output_count == 20'd0) & (ap_start == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((dataflow_in_loop_TOP_LOOP38116_U0_ap_ready == 1'b1) & (loop_dataflow_input_count == bound_minus_1) & (ap_start == 1'b1))) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((~(loop_dataflow_output_count == bound_minus_1) | (ap_continue == 1'b1))) begin
        dataflow_in_loop_TOP_LOOP38116_U0_ap_continue = 1'b1;
    end else begin
        dataflow_in_loop_TOP_LOOP38116_U0_ap_continue = 1'b0;
    end
end

assign adjustments_address0 = dataflow_in_loop_TOP_LOOP38116_U0_adjustments_address0;

assign adjustments_address1 = 4'd0;

assign adjustments_ce0 = dataflow_in_loop_TOP_LOOP38116_U0_adjustments_ce0;

assign adjustments_ce1 = 1'b0;

assign adjustments_d0 = 48'd0;

assign adjustments_d1 = 48'd0;

assign adjustments_we0 = 1'b0;

assign adjustments_we1 = 1'b0;

assign ap_sync_continue = ap_continue;

assign ap_sync_done = dataflow_in_loop_TOP_LOOP38116_U0_ap_done;

assign ap_sync_ready = dataflow_in_loop_TOP_LOOP38116_U0_ap_ready;

assign bound_minus_1 = (20'd802816 - 20'd1);

assign dataflow_in_loop_TOP_LOOP38116_U0_ap_start = ap_start;

assign dataflow_in_loop_TOP_LOOP38116_U0_in_data_full_n = in_data_empty_n;

assign dataflow_in_loop_TOP_LOOP38116_U0_in_data_write = 1'b0;

assign dataflow_in_loop_TOP_LOOP38116_U0_start_full_n = 1'b1;

assign dataflow_in_loop_TOP_LOOP38116_U0_start_write = 1'b0;

assign filter_data_address0 = dataflow_in_loop_TOP_LOOP38116_U0_filter_data_address0;

assign filter_data_address1 = 9'd0;

assign filter_data_ce0 = dataflow_in_loop_TOP_LOOP38116_U0_filter_data_ce0;

assign filter_data_ce1 = 1'b0;

assign filter_data_d0 = 16'd0;

assign filter_data_d1 = 16'd0;

assign filter_data_we0 = 1'b0;

assign filter_data_we1 = 1'b0;

assign in_data_address0 = dataflow_in_loop_TOP_LOOP38116_U0_in_data_address0;

assign in_data_address1 = 16'd0;

assign in_data_ce0 = dataflow_in_loop_TOP_LOOP38116_U0_in_data_ce0;

assign in_data_ce1 = 1'b0;

assign in_data_d0 = 64'd0;

assign in_data_d1 = 64'd0;

assign in_data_read = dataflow_in_loop_TOP_LOOP38116_U0_in_data_write;

assign in_data_we0 = 1'b0;

assign in_data_we1 = 1'b0;

assign out_data_address0 = 16'd0;

assign out_data_address1 = dataflow_in_loop_TOP_LOOP38116_U0_out_data_address1;

assign out_data_ce0 = 1'b0;

assign out_data_ce1 = dataflow_in_loop_TOP_LOOP38116_U0_out_data_ce1;

assign out_data_d0 = 64'd0;

assign out_data_d1 = dataflow_in_loop_TOP_LOOP38116_U0_out_data_d1;

assign out_data_we0 = 1'b0;

assign out_data_we1 = dataflow_in_loop_TOP_LOOP38116_U0_out_data_we1;

assign out_data_write = dataflow_in_loop_TOP_LOOP38116_U0_out_data_write;

endmodule //td_fused_top_tdf1_114
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf11_14 (
        in_data_address0,
        in_data_ce0,
        in_data_d0,
        in_data_q0,
        in_data_we0,
        in_data_address1,
        in_data_ce1,
        in_data_d1,
        in_data_q1,
        in_data_we1,
        out_data_address0,
        out_data_ce0,
        out_data_d0,
        out_data_q0,
        out_data_we0,
        out_data_address1,
        out_data_ce1,
        out_data_d1,
        out_data_q1,
        out_data_we1,
        l1_filter_data_address0,
        l1_filter_data_ce0,
        l1_filter_data_d0,
        l1_filter_data_q0,
        l1_filter_data_we0,
        l1_filter_data_address1,
        l1_filter_data_ce1,
        l1_filter_data_d1,
        l1_filter_data_q1,
        l1_filter_data_we1,
        l2_filter_data_address0,
        l2_filter_data_ce0,
        l2_filter_data_d0,
        l2_filter_data_q0,
        l2_filter_data_we0,
        l2_filter_data_address1,
        l2_filter_data_ce1,
        l2_filter_data_d1,
        l2_filter_data_q1,
        l2_filter_data_we1,
        l1_adjustments_address0,
        l1_adjustments_ce0,
        l1_adjustments_d0,
        l1_adjustments_q0,
        l1_adjustments_we0,
        l1_adjustments_address1,
        l1_adjustments_ce1,
        l1_adjustments_d1,
        l1_adjustments_q1,
        l1_adjustments_we1,
        l2_adjustments_address0,
        l2_adjustments_ce0,
        l2_adjustments_d0,
        l2_adjustments_q0,
        l2_adjustments_we0,
        l2_adjustments_address1,
        l2_adjustments_ce1,
        l2_adjustments_d1,
        l2_adjustments_q1,
        l2_adjustments_we1,
        ap_clk,
        ap_rst,
        in_data_empty_n,
        in_data_read,
        out_data_full_n,
        out_data_write,
        ap_start,
        ap_done,
        ap_ready,
        ap_idle,
        ap_continue
);


output  [11:0] in_data_address0;
output   in_data_ce0;
output  [63:0] in_data_d0;
input  [63:0] in_data_q0;
output   in_data_we0;
output  [11:0] in_data_address1;
output   in_data_ce1;
output  [63:0] in_data_d1;
input  [63:0] in_data_q1;
output   in_data_we1;
output  [12:0] out_data_address0;
output   out_data_ce0;
output  [63:0] out_data_d0;
input  [63:0] out_data_q0;
output   out_data_we0;
output  [12:0] out_data_address1;
output   out_data_ce1;
output  [63:0] out_data_d1;
input  [63:0] out_data_q1;
output   out_data_we1;
output  [16:0] l1_filter_data_address0;
output   l1_filter_data_ce0;
output  [63:0] l1_filter_data_d0;
input  [63:0] l1_filter_data_q0;
output   l1_filter_data_we0;
output  [16:0] l1_filter_data_address1;
output   l1_filter_data_ce1;
output  [63:0] l1_filter_data_d1;
input  [63:0] l1_filter_data_q1;
output   l1_filter_data_we1;
output  [15:0] l2_filter_data_address0;
output   l2_filter_data_ce0;
output  [15:0] l2_filter_data_d0;
input  [15:0] l2_filter_data_q0;
output   l2_filter_data_we0;
output  [15:0] l2_filter_data_address1;
output   l2_filter_data_ce1;
output  [15:0] l2_filter_data_d1;
input  [15:0] l2_filter_data_q1;
output   l2_filter_data_we1;
output  [8:0] l1_adjustments_address0;
output   l1_adjustments_ce0;
output  [47:0] l1_adjustments_d0;
input  [47:0] l1_adjustments_q0;
output   l1_adjustments_we0;
output  [8:0] l1_adjustments_address1;
output   l1_adjustments_ce1;
output  [47:0] l1_adjustments_d1;
input  [47:0] l1_adjustments_q1;
output   l1_adjustments_we1;
output  [6:0] l2_adjustments_address0;
output   l2_adjustments_ce0;
output  [47:0] l2_adjustments_d0;
input  [47:0] l2_adjustments_q0;
output   l2_adjustments_we0;
output  [6:0] l2_adjustments_address1;
output   l2_adjustments_ce1;
output  [47:0] l2_adjustments_d1;
input  [47:0] l2_adjustments_q1;
output   l2_adjustments_we1;
input   ap_clk;
input   ap_rst;
input   in_data_empty_n;
output   in_data_read;
input   out_data_full_n;
output   out_data_write;
input   ap_start;
output   ap_done;
output   ap_ready;
output   ap_idle;
input   ap_continue;

reg ap_done;
reg ap_ready;
reg ap_idle;

wire   [11:0] dataflow_in_loop_TOP_LOOP38270_U0_in_data_address0;
wire    dataflow_in_loop_TOP_LOOP38270_U0_in_data_ce0;
wire   [63:0] dataflow_in_loop_TOP_LOOP38270_U0_in_data_d0;
wire    dataflow_in_loop_TOP_LOOP38270_U0_in_data_we0;
wire   [11:0] dataflow_in_loop_TOP_LOOP38270_U0_in_data_address1;
wire    dataflow_in_loop_TOP_LOOP38270_U0_in_data_ce1;
wire   [63:0] dataflow_in_loop_TOP_LOOP38270_U0_in_data_d1;
wire    dataflow_in_loop_TOP_LOOP38270_U0_in_data_we1;
wire   [16:0] dataflow_in_loop_TOP_LOOP38270_U0_l1_filter_data_address0;
wire    dataflow_in_loop_TOP_LOOP38270_U0_l1_filter_data_ce0;
wire   [63:0] dataflow_in_loop_TOP_LOOP38270_U0_l1_filter_data_d0;
wire    dataflow_in_loop_TOP_LOOP38270_U0_l1_filter_data_we0;
wire   [16:0] dataflow_in_loop_TOP_LOOP38270_U0_l1_filter_data_address1;
wire    dataflow_in_loop_TOP_LOOP38270_U0_l1_filter_data_ce1;
wire   [63:0] dataflow_in_loop_TOP_LOOP38270_U0_l1_filter_data_d1;
wire    dataflow_in_loop_TOP_LOOP38270_U0_l1_filter_data_we1;
wire   [8:0] dataflow_in_loop_TOP_LOOP38270_U0_l1_adjustments_address0;
wire    dataflow_in_loop_TOP_LOOP38270_U0_l1_adjustments_ce0;
wire   [47:0] dataflow_in_loop_TOP_LOOP38270_U0_l1_adjustments_d0;
wire    dataflow_in_loop_TOP_LOOP38270_U0_l1_adjustments_we0;
wire   [8:0] dataflow_in_loop_TOP_LOOP38270_U0_l1_adjustments_address1;
wire    dataflow_in_loop_TOP_LOOP38270_U0_l1_adjustments_ce1;
wire   [47:0] dataflow_in_loop_TOP_LOOP38270_U0_l1_adjustments_d1;
wire    dataflow_in_loop_TOP_LOOP38270_U0_l1_adjustments_we1;
wire   [15:0] dataflow_in_loop_TOP_LOOP38270_U0_l2_filter_data_address0;
wire    dataflow_in_loop_TOP_LOOP38270_U0_l2_filter_data_ce0;
wire   [15:0] dataflow_in_loop_TOP_LOOP38270_U0_l2_filter_data_d0;
wire    dataflow_in_loop_TOP_LOOP38270_U0_l2_filter_data_we0;
wire   [15:0] dataflow_in_loop_TOP_LOOP38270_U0_l2_filter_data_address1;
wire    dataflow_in_loop_TOP_LOOP38270_U0_l2_filter_data_ce1;
wire   [15:0] dataflow_in_loop_TOP_LOOP38270_U0_l2_filter_data_d1;
wire    dataflow_in_loop_TOP_LOOP38270_U0_l2_filter_data_we1;
wire   [12:0] dataflow_in_loop_TOP_LOOP38270_U0_out_data_address0;
wire    dataflow_in_loop_TOP_LOOP38270_U0_out_data_ce0;
wire   [63:0] dataflow_in_loop_TOP_LOOP38270_U0_out_data_d0;
wire    dataflow_in_loop_TOP_LOOP38270_U0_out_data_we0;
wire   [12:0] dataflow_in_loop_TOP_LOOP38270_U0_out_data_address1;
wire    dataflow_in_loop_TOP_LOOP38270_U0_out_data_ce1;
wire   [63:0] dataflow_in_loop_TOP_LOOP38270_U0_out_data_d1;
wire    dataflow_in_loop_TOP_LOOP38270_U0_out_data_we1;
wire   [6:0] dataflow_in_loop_TOP_LOOP38270_U0_l2_adjustments_address0;
wire    dataflow_in_loop_TOP_LOOP38270_U0_l2_adjustments_ce0;
wire   [47:0] dataflow_in_loop_TOP_LOOP38270_U0_l2_adjustments_d0;
wire    dataflow_in_loop_TOP_LOOP38270_U0_l2_adjustments_we0;
wire   [6:0] dataflow_in_loop_TOP_LOOP38270_U0_l2_adjustments_address1;
wire    dataflow_in_loop_TOP_LOOP38270_U0_l2_adjustments_ce1;
wire   [47:0] dataflow_in_loop_TOP_LOOP38270_U0_l2_adjustments_d1;
wire    dataflow_in_loop_TOP_LOOP38270_U0_l2_adjustments_we1;
wire    dataflow_in_loop_TOP_LOOP38270_U0_ap_start;
wire    dataflow_in_loop_TOP_LOOP38270_U0_in_data_read;
wire    dataflow_in_loop_TOP_LOOP38270_U0_out_data_write;
wire    dataflow_in_loop_TOP_LOOP38270_U0_ap_done;
wire    dataflow_in_loop_TOP_LOOP38270_U0_ap_ready;
wire    dataflow_in_loop_TOP_LOOP38270_U0_ap_idle;
reg    dataflow_in_loop_TOP_LOOP38270_U0_ap_continue;
wire    dataflow_in_loop_TOP_LOOP38270_U0_in_data_full_n;
wire    dataflow_in_loop_TOP_LOOP38270_U0_in_data_write;
wire    ap_sync_continue;
wire    ap_sync_done;
wire    ap_sync_ready;
reg   [16:0] loop_dataflow_input_count;
reg   [16:0] loop_dataflow_output_count;
wire   [16:0] bound_minus_1;
wire    dataflow_in_loop_TOP_LOOP38270_U0_start_full_n;
wire    dataflow_in_loop_TOP_LOOP38270_U0_start_write;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 loop_dataflow_input_count = 17'd0;
#0 loop_dataflow_output_count = 17'd0;
end

td_fused_top_dataflow_in_loop_TOP_LOOP38270 dataflow_in_loop_TOP_LOOP38270_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .in_data_address0(dataflow_in_loop_TOP_LOOP38270_U0_in_data_address0),
    .in_data_ce0(dataflow_in_loop_TOP_LOOP38270_U0_in_data_ce0),
    .in_data_d0(dataflow_in_loop_TOP_LOOP38270_U0_in_data_d0),
    .in_data_q0(in_data_q0),
    .in_data_we0(dataflow_in_loop_TOP_LOOP38270_U0_in_data_we0),
    .in_data_address1(dataflow_in_loop_TOP_LOOP38270_U0_in_data_address1),
    .in_data_ce1(dataflow_in_loop_TOP_LOOP38270_U0_in_data_ce1),
    .in_data_d1(dataflow_in_loop_TOP_LOOP38270_U0_in_data_d1),
    .in_data_q1(64'd0),
    .in_data_we1(dataflow_in_loop_TOP_LOOP38270_U0_in_data_we1),
    .l1_filter_data_address0(dataflow_in_loop_TOP_LOOP38270_U0_l1_filter_data_address0),
    .l1_filter_data_ce0(dataflow_in_loop_TOP_LOOP38270_U0_l1_filter_data_ce0),
    .l1_filter_data_d0(dataflow_in_loop_TOP_LOOP38270_U0_l1_filter_data_d0),
    .l1_filter_data_q0(l1_filter_data_q0),
    .l1_filter_data_we0(dataflow_in_loop_TOP_LOOP38270_U0_l1_filter_data_we0),
    .l1_filter_data_address1(dataflow_in_loop_TOP_LOOP38270_U0_l1_filter_data_address1),
    .l1_filter_data_ce1(dataflow_in_loop_TOP_LOOP38270_U0_l1_filter_data_ce1),
    .l1_filter_data_d1(dataflow_in_loop_TOP_LOOP38270_U0_l1_filter_data_d1),
    .l1_filter_data_q1(64'd0),
    .l1_filter_data_we1(dataflow_in_loop_TOP_LOOP38270_U0_l1_filter_data_we1),
    .l1_adjustments_address0(dataflow_in_loop_TOP_LOOP38270_U0_l1_adjustments_address0),
    .l1_adjustments_ce0(dataflow_in_loop_TOP_LOOP38270_U0_l1_adjustments_ce0),
    .l1_adjustments_d0(dataflow_in_loop_TOP_LOOP38270_U0_l1_adjustments_d0),
    .l1_adjustments_q0(l1_adjustments_q0),
    .l1_adjustments_we0(dataflow_in_loop_TOP_LOOP38270_U0_l1_adjustments_we0),
    .l1_adjustments_address1(dataflow_in_loop_TOP_LOOP38270_U0_l1_adjustments_address1),
    .l1_adjustments_ce1(dataflow_in_loop_TOP_LOOP38270_U0_l1_adjustments_ce1),
    .l1_adjustments_d1(dataflow_in_loop_TOP_LOOP38270_U0_l1_adjustments_d1),
    .l1_adjustments_q1(48'd0),
    .l1_adjustments_we1(dataflow_in_loop_TOP_LOOP38270_U0_l1_adjustments_we1),
    .l2_filter_data_address0(dataflow_in_loop_TOP_LOOP38270_U0_l2_filter_data_address0),
    .l2_filter_data_ce0(dataflow_in_loop_TOP_LOOP38270_U0_l2_filter_data_ce0),
    .l2_filter_data_d0(dataflow_in_loop_TOP_LOOP38270_U0_l2_filter_data_d0),
    .l2_filter_data_q0(l2_filter_data_q0),
    .l2_filter_data_we0(dataflow_in_loop_TOP_LOOP38270_U0_l2_filter_data_we0),
    .l2_filter_data_address1(dataflow_in_loop_TOP_LOOP38270_U0_l2_filter_data_address1),
    .l2_filter_data_ce1(dataflow_in_loop_TOP_LOOP38270_U0_l2_filter_data_ce1),
    .l2_filter_data_d1(dataflow_in_loop_TOP_LOOP38270_U0_l2_filter_data_d1),
    .l2_filter_data_q1(16'd0),
    .l2_filter_data_we1(dataflow_in_loop_TOP_LOOP38270_U0_l2_filter_data_we1),
    .out_data_address0(dataflow_in_loop_TOP_LOOP38270_U0_out_data_address0),
    .out_data_ce0(dataflow_in_loop_TOP_LOOP38270_U0_out_data_ce0),
    .out_data_d0(dataflow_in_loop_TOP_LOOP38270_U0_out_data_d0),
    .out_data_q0(64'd0),
    .out_data_we0(dataflow_in_loop_TOP_LOOP38270_U0_out_data_we0),
    .out_data_address1(dataflow_in_loop_TOP_LOOP38270_U0_out_data_address1),
    .out_data_ce1(dataflow_in_loop_TOP_LOOP38270_U0_out_data_ce1),
    .out_data_d1(dataflow_in_loop_TOP_LOOP38270_U0_out_data_d1),
    .out_data_q1(64'd0),
    .out_data_we1(dataflow_in_loop_TOP_LOOP38270_U0_out_data_we1),
    .l2_adjustments_address0(dataflow_in_loop_TOP_LOOP38270_U0_l2_adjustments_address0),
    .l2_adjustments_ce0(dataflow_in_loop_TOP_LOOP38270_U0_l2_adjustments_ce0),
    .l2_adjustments_d0(dataflow_in_loop_TOP_LOOP38270_U0_l2_adjustments_d0),
    .l2_adjustments_q0(l2_adjustments_q0),
    .l2_adjustments_we0(dataflow_in_loop_TOP_LOOP38270_U0_l2_adjustments_we0),
    .l2_adjustments_address1(dataflow_in_loop_TOP_LOOP38270_U0_l2_adjustments_address1),
    .l2_adjustments_ce1(dataflow_in_loop_TOP_LOOP38270_U0_l2_adjustments_ce1),
    .l2_adjustments_d1(dataflow_in_loop_TOP_LOOP38270_U0_l2_adjustments_d1),
    .l2_adjustments_q1(48'd0),
    .l2_adjustments_we1(dataflow_in_loop_TOP_LOOP38270_U0_l2_adjustments_we1),
    .ap_start(dataflow_in_loop_TOP_LOOP38270_U0_ap_start),
    .in_data_empty_n(1'b0),
    .in_data_read(dataflow_in_loop_TOP_LOOP38270_U0_in_data_read),
    .out_data_full_n(out_data_full_n),
    .out_data_write(dataflow_in_loop_TOP_LOOP38270_U0_out_data_write),
    .ap_done(dataflow_in_loop_TOP_LOOP38270_U0_ap_done),
    .ap_ready(dataflow_in_loop_TOP_LOOP38270_U0_ap_ready),
    .ap_idle(dataflow_in_loop_TOP_LOOP38270_U0_ap_idle),
    .ap_continue(dataflow_in_loop_TOP_LOOP38270_U0_ap_continue)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        loop_dataflow_input_count <= 17'd0;
    end else begin
        if ((~(loop_dataflow_input_count == bound_minus_1) & (ap_start == 1'b1) & (dataflow_in_loop_TOP_LOOP38270_U0_ap_ready == 1'b1))) begin
            loop_dataflow_input_count <= (loop_dataflow_input_count + 17'd1);
        end else if (((loop_dataflow_input_count == bound_minus_1) & (ap_start == 1'b1) & (dataflow_in_loop_TOP_LOOP38270_U0_ap_ready == 1'b1))) begin
            loop_dataflow_input_count <= 17'd0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        loop_dataflow_output_count <= 17'd0;
    end else begin
        if ((~(loop_dataflow_output_count == bound_minus_1) & (dataflow_in_loop_TOP_LOOP38270_U0_ap_continue == 1'b1) & (dataflow_in_loop_TOP_LOOP38270_U0_ap_done == 1'b1))) begin
            loop_dataflow_output_count <= (loop_dataflow_output_count + 17'd1);
        end else if (((loop_dataflow_output_count == bound_minus_1) & (dataflow_in_loop_TOP_LOOP38270_U0_ap_continue == 1'b1) & (dataflow_in_loop_TOP_LOOP38270_U0_ap_done == 1'b1))) begin
            loop_dataflow_output_count <= 17'd0;
        end
    end
end

always @ (*) begin
    if (((loop_dataflow_output_count == bound_minus_1) & (dataflow_in_loop_TOP_LOOP38270_U0_ap_done == 1'b1))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = 1'b0;
    end
end

always @ (*) begin
    if (((loop_dataflow_output_count == 17'd0) & (ap_start == 1'b0) & (dataflow_in_loop_TOP_LOOP38270_U0_ap_idle == 1'b1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((loop_dataflow_input_count == bound_minus_1) & (ap_start == 1'b1) & (dataflow_in_loop_TOP_LOOP38270_U0_ap_ready == 1'b1))) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((~(loop_dataflow_output_count == bound_minus_1) | (ap_continue == 1'b1))) begin
        dataflow_in_loop_TOP_LOOP38270_U0_ap_continue = 1'b1;
    end else begin
        dataflow_in_loop_TOP_LOOP38270_U0_ap_continue = 1'b0;
    end
end

assign ap_sync_continue = ap_continue;

assign ap_sync_done = dataflow_in_loop_TOP_LOOP38270_U0_ap_done;

assign ap_sync_ready = dataflow_in_loop_TOP_LOOP38270_U0_ap_ready;

assign bound_minus_1 = (17'd100352 - 17'd1);

assign dataflow_in_loop_TOP_LOOP38270_U0_ap_start = ap_start;

assign dataflow_in_loop_TOP_LOOP38270_U0_in_data_full_n = in_data_empty_n;

assign dataflow_in_loop_TOP_LOOP38270_U0_in_data_write = 1'b0;

assign dataflow_in_loop_TOP_LOOP38270_U0_start_full_n = 1'b1;

assign dataflow_in_loop_TOP_LOOP38270_U0_start_write = 1'b0;

assign in_data_address0 = dataflow_in_loop_TOP_LOOP38270_U0_in_data_address0;

assign in_data_address1 = 12'd0;

assign in_data_ce0 = dataflow_in_loop_TOP_LOOP38270_U0_in_data_ce0;

assign in_data_ce1 = 1'b0;

assign in_data_d0 = 64'd0;

assign in_data_d1 = 64'd0;

assign in_data_read = dataflow_in_loop_TOP_LOOP38270_U0_in_data_write;

assign in_data_we0 = 1'b0;

assign in_data_we1 = 1'b0;

assign l1_adjustments_address0 = dataflow_in_loop_TOP_LOOP38270_U0_l1_adjustments_address0;

assign l1_adjustments_address1 = 9'd0;

assign l1_adjustments_ce0 = dataflow_in_loop_TOP_LOOP38270_U0_l1_adjustments_ce0;

assign l1_adjustments_ce1 = 1'b0;

assign l1_adjustments_d0 = 48'd0;

assign l1_adjustments_d1 = 48'd0;

assign l1_adjustments_we0 = 1'b0;

assign l1_adjustments_we1 = 1'b0;

assign l1_filter_data_address0 = dataflow_in_loop_TOP_LOOP38270_U0_l1_filter_data_address0;

assign l1_filter_data_address1 = 17'd0;

assign l1_filter_data_ce0 = dataflow_in_loop_TOP_LOOP38270_U0_l1_filter_data_ce0;

assign l1_filter_data_ce1 = 1'b0;

assign l1_filter_data_d0 = 64'd0;

assign l1_filter_data_d1 = 64'd0;

assign l1_filter_data_we0 = 1'b0;

assign l1_filter_data_we1 = 1'b0;

assign l2_adjustments_address0 = dataflow_in_loop_TOP_LOOP38270_U0_l2_adjustments_address0;

assign l2_adjustments_address1 = 7'd0;

assign l2_adjustments_ce0 = dataflow_in_loop_TOP_LOOP38270_U0_l2_adjustments_ce0;

assign l2_adjustments_ce1 = 1'b0;

assign l2_adjustments_d0 = 48'd0;

assign l2_adjustments_d1 = 48'd0;

assign l2_adjustments_we0 = 1'b0;

assign l2_adjustments_we1 = 1'b0;

assign l2_filter_data_address0 = dataflow_in_loop_TOP_LOOP38270_U0_l2_filter_data_address0;

assign l2_filter_data_address1 = 16'd0;

assign l2_filter_data_ce0 = dataflow_in_loop_TOP_LOOP38270_U0_l2_filter_data_ce0;

assign l2_filter_data_ce1 = 1'b0;

assign l2_filter_data_d0 = 16'd0;

assign l2_filter_data_d1 = 16'd0;

assign l2_filter_data_we0 = 1'b0;

assign l2_filter_data_we1 = 1'b0;

assign out_data_address0 = 13'd0;

assign out_data_address1 = dataflow_in_loop_TOP_LOOP38270_U0_out_data_address1;

assign out_data_ce0 = 1'b0;

assign out_data_ce1 = dataflow_in_loop_TOP_LOOP38270_U0_out_data_ce1;

assign out_data_d0 = 64'd0;

assign out_data_d1 = dataflow_in_loop_TOP_LOOP38270_U0_out_data_d1;

assign out_data_we0 = 1'b0;

assign out_data_we1 = dataflow_in_loop_TOP_LOOP38270_U0_out_data_we1;

assign out_data_write = dataflow_in_loop_TOP_LOOP38270_U0_out_data_write;

endmodule //td_fused_top_tdf11_14
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf11_accum_1 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        accum_in_0_address0,
        accum_in_0_ce0,
        accum_in_0_q0,
        accum_in_0_address1,
        accum_in_0_ce1,
        accum_in_0_q1,
        accum_out_address0,
        accum_out_ce0,
        accum_out_we0,
        accum_out_d0,
        accum_out_address1,
        accum_out_ce1,
        accum_out_we1,
        accum_out_d1
);

parameter    ap_ST_fsm_state1 = 8'd1;
parameter    ap_ST_fsm_pp0_stage0 = 8'd2;
parameter    ap_ST_fsm_pp0_stage1 = 8'd4;
parameter    ap_ST_fsm_pp0_stage2 = 8'd8;
parameter    ap_ST_fsm_pp0_stage3 = 8'd16;
parameter    ap_ST_fsm_state12 = 8'd32;
parameter    ap_ST_fsm_state13 = 8'd64;
parameter    ap_ST_fsm_state14 = 8'd128;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [9:0] accum_in_0_address0;
output   accum_in_0_ce0;
input  [15:0] accum_in_0_q0;
output  [9:0] accum_in_0_address1;
output   accum_in_0_ce1;
input  [15:0] accum_in_0_q1;
output  [2:0] accum_out_address0;
output   accum_out_ce0;
output   accum_out_we0;
output  [15:0] accum_out_d0;
output  [2:0] accum_out_address1;
output   accum_out_ce1;
output   accum_out_we1;
output  [15:0] accum_out_d1;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg[9:0] accum_in_0_address0;
reg accum_in_0_ce0;
reg[9:0] accum_in_0_address1;
reg accum_in_0_ce1;
reg accum_out_ce0;
reg accum_out_we0;
reg accum_out_ce1;
reg accum_out_we1;

reg    ap_done_reg;
  reg   [7:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg   [9:0] x_reg_168;
reg   [15:0] psum_7_08_reg_180;
reg   [15:0] psum_6_07_reg_192;
reg   [15:0] psum_5_06_reg_204;
reg   [15:0] psum_4_05_reg_216;
reg   [15:0] psum_3_04_reg_228;
reg   [15:0] psum_2_03_reg_240;
reg   [15:0] psum_1_02_reg_252;
reg   [15:0] psum_0_01_reg_264;
wire   [0:0] icmp_ln132_fu_321_p2;
reg   [0:0] icmp_ln132_reg_492;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state6_pp0_stage0_iter1;
wire    ap_block_state10_pp0_stage0_iter2;
wire    ap_block_pp0_stage0_11001;
reg   [0:0] icmp_ln132_reg_492_pp0_iter1_reg;
reg   [0:0] icmp_ln132_reg_492_pp0_iter2_reg;
reg   [15:0] accum_in_0_load_reg_506;
wire    ap_CS_fsm_pp0_stage1;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_state3_pp0_stage1_iter0;
wire    ap_block_state7_pp0_stage1_iter1;
wire    ap_block_state11_pp0_stage1_iter2;
wire    ap_block_pp0_stage1_11001;
reg   [15:0] accum_in_0_load_65_reg_511;
reg   [15:0] accum_in_0_load_66_reg_526;
wire    ap_CS_fsm_pp0_stage2;
wire    ap_block_state4_pp0_stage2_iter0;
wire    ap_block_state8_pp0_stage2_iter1;
wire    ap_block_pp0_stage2_11001;
reg   [15:0] accum_in_0_load_67_reg_531;
wire   [9:0] add_ln132_fu_387_p2;
reg   [9:0] add_ln132_reg_546;
wire    ap_CS_fsm_pp0_stage3;
wire    ap_block_state5_pp0_stage3_iter0;
wire    ap_block_state9_pp0_stage3_iter1;
wire    ap_block_pp0_stage3_11001;
reg   [15:0] accum_in_0_load_68_reg_551;
reg   [15:0] accum_in_0_load_69_reg_556;
reg   [15:0] accum_in_0_load_70_reg_571;
reg    ap_enable_reg_pp0_iter1;
reg   [15:0] accum_in_0_load_71_reg_576;
wire   [15:0] grp_fu_305_p2;
wire   [15:0] grp_fu_310_p2;
reg    ap_enable_reg_pp0_iter2;
wire   [3:0] add_ln140_fu_432_p2;
wire    ap_CS_fsm_state13;
wire   [0:0] tmp_fu_415_p3;
reg    ap_block_state1;
wire    ap_block_pp0_stage2_subdone;
reg    ap_condition_pp0_exit_iter0_state4;
wire    ap_block_pp0_stage3_subdone;
wire    ap_block_pp0_stage1_subdone;
reg   [9:0] ap_phi_mux_x_phi_fu_172_p4;
wire    ap_block_pp0_stage0;
wire   [15:0] ap_phi_mux_psum_7_08_phi_fu_184_p4;
wire    ap_block_pp0_stage1;
wire   [15:0] ap_phi_mux_psum_6_07_phi_fu_196_p4;
wire   [15:0] ap_phi_mux_psum_5_06_phi_fu_208_p4;
wire   [15:0] ap_phi_mux_psum_4_05_phi_fu_220_p4;
wire   [15:0] ap_phi_mux_psum_3_04_phi_fu_232_p4;
wire    ap_block_pp0_stage3;
wire   [15:0] ap_phi_mux_psum_2_03_phi_fu_244_p4;
wire    ap_block_pp0_stage2;
reg   [3:0] q_reg_276;
wire    ap_CS_fsm_state12;
reg   [15:0] ap_phi_mux_phi_ln152_phi_fu_290_p8;
wire   [2:0] trunc_ln140_fu_428_p1;
wire   [63:0] zext_ln132_fu_327_p1;
wire   [63:0] zext_ln136_fu_338_p1;
wire   [63:0] zext_ln136_13_fu_349_p1;
wire   [63:0] zext_ln136_14_fu_360_p1;
wire   [63:0] zext_ln136_15_fu_371_p1;
wire   [63:0] zext_ln136_16_fu_382_p1;
wire   [63:0] zext_ln136_17_fu_399_p1;
wire   [63:0] zext_ln136_18_fu_410_p1;
wire   [63:0] zext_ln140_fu_423_p1;
wire   [63:0] zext_ln140_3_fu_444_p1;
reg   [15:0] grp_fu_305_p0;
reg   [15:0] grp_fu_305_p1;
reg   [15:0] grp_fu_310_p0;
reg   [15:0] grp_fu_310_p1;
wire   [9:0] or_ln136_fu_332_p2;
wire   [9:0] or_ln136_13_fu_343_p2;
wire   [9:0] or_ln136_14_fu_354_p2;
wire   [9:0] or_ln136_15_fu_365_p2;
wire   [9:0] or_ln136_16_fu_376_p2;
wire   [9:0] or_ln136_17_fu_393_p2;
wire   [9:0] or_ln136_18_fu_404_p2;
wire   [2:0] or_ln140_fu_438_p2;
wire   [0:0] icmp_ln152_fu_449_p2;
wire   [0:0] icmp_ln152_5_fu_463_p2;
wire   [15:0] select_ln152_fu_455_p3;
wire   [0:0] icmp_ln152_6_fu_477_p2;
wire   [15:0] select_ln152_5_fu_469_p3;
wire    ap_CS_fsm_state14;
reg   [7:0] ap_NS_fsm;
wire    ap_block_pp0_stage0_subdone;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
reg    ap_condition_514;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 8'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
end

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U699(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(grp_fu_305_p0),
    .din1(grp_fu_305_p1),
    .dout(grp_fu_305_p2)
);

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U700(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(grp_fu_310_p0),
    .din1(grp_fu_310_p1),
    .dout(grp_fu_310_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state14)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage2_subdone) & (1'b1 == ap_condition_pp0_exit_iter0_state4) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage3_subdone) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b0)) | ((1'b0 == ap_block_pp0_stage3_subdone) & (1'b1 == ap_CS_fsm_pp0_stage3)))) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end else if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter2 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state12)) begin
        q_reg_276 <= 4'd0;
    end else if (((tmp_fu_415_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state13))) begin
        q_reg_276 <= add_ln140_fu_432_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln132_reg_492 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        x_reg_168 <= add_ln132_reg_546;
    end else if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        x_reg_168 <= 10'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage1_11001) & (icmp_ln132_reg_492 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
        accum_in_0_load_65_reg_511 <= accum_in_0_q0;
        accum_in_0_load_reg_506 <= accum_in_0_q1;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2_11001) & (icmp_ln132_reg_492 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
        accum_in_0_load_66_reg_526 <= accum_in_0_q1;
        accum_in_0_load_67_reg_531 <= accum_in_0_q0;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage3_11001) & (icmp_ln132_reg_492 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
        accum_in_0_load_68_reg_551 <= accum_in_0_q1;
        accum_in_0_load_69_reg_556 <= accum_in_0_q0;
        add_ln132_reg_546 <= add_ln132_fu_387_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln132_reg_492 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        accum_in_0_load_70_reg_571 <= accum_in_0_q1;
        accum_in_0_load_71_reg_576 <= accum_in_0_q0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln132_reg_492 <= icmp_ln132_fu_321_p2;
        icmp_ln132_reg_492_pp0_iter1_reg <= icmp_ln132_reg_492;
        icmp_ln132_reg_492_pp0_iter2_reg <= icmp_ln132_reg_492_pp0_iter1_reg;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln132_reg_492_pp0_iter1_reg == 1'd1) & (1'b0 == ap_block_pp0_stage2_11001) & (1'b1 == ap_CS_fsm_pp0_stage2) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        psum_0_01_reg_264 <= grp_fu_305_p2;
        psum_1_02_reg_252 <= grp_fu_310_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln132_reg_492_pp0_iter1_reg == 1'd1) & (1'b0 == ap_block_pp0_stage3_11001) & (1'b1 == ap_CS_fsm_pp0_stage3) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        psum_2_03_reg_240 <= grp_fu_305_p2;
        psum_3_04_reg_228 <= grp_fu_310_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln132_reg_492_pp0_iter1_reg == 1'd1) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        psum_4_05_reg_216 <= grp_fu_305_p2;
        psum_5_06_reg_204 <= grp_fu_310_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln132_reg_492_pp0_iter2_reg == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        psum_6_07_reg_192 <= grp_fu_305_p2;
        psum_7_08_reg_180 <= grp_fu_310_p2;
    end
end

always @ (*) begin
    if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
        if (((1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            accum_in_0_address0 = zext_ln136_18_fu_410_p1;
        end else if (((1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            accum_in_0_address0 = zext_ln136_16_fu_382_p1;
        end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            accum_in_0_address0 = zext_ln136_14_fu_360_p1;
        end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            accum_in_0_address0 = zext_ln136_fu_338_p1;
        end else begin
            accum_in_0_address0 = 'bx;
        end
    end else begin
        accum_in_0_address0 = 'bx;
    end
end

always @ (*) begin
    if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
        if (((1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            accum_in_0_address1 = zext_ln136_17_fu_399_p1;
        end else if (((1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            accum_in_0_address1 = zext_ln136_15_fu_371_p1;
        end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            accum_in_0_address1 = zext_ln136_13_fu_349_p1;
        end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            accum_in_0_address1 = zext_ln132_fu_327_p1;
        end else begin
            accum_in_0_address1 = 'bx;
        end
    end else begin
        accum_in_0_address1 = 'bx;
    end
end

always @ (*) begin
    if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage3_11001) & (1'b1 == ap_CS_fsm_pp0_stage3)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2_11001) & (1'b1 == ap_CS_fsm_pp0_stage2)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1)))) begin
        accum_in_0_ce0 = 1'b1;
    end else begin
        accum_in_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage3_11001) & (1'b1 == ap_CS_fsm_pp0_stage3)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2_11001) & (1'b1 == ap_CS_fsm_pp0_stage2)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1)))) begin
        accum_in_0_ce1 = 1'b1;
    end else begin
        accum_in_0_ce1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state13)) begin
        accum_out_ce0 = 1'b1;
    end else begin
        accum_out_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state13)) begin
        accum_out_ce1 = 1'b1;
    end else begin
        accum_out_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((tmp_fu_415_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state13))) begin
        accum_out_we0 = 1'b1;
    end else begin
        accum_out_we0 = 1'b0;
    end
end

always @ (*) begin
    if (((tmp_fu_415_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state13))) begin
        accum_out_we1 = 1'b1;
    end else begin
        accum_out_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((icmp_ln132_reg_492 == 1'd0)) begin
        ap_condition_pp0_exit_iter0_state4 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state4 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state14)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((tmp_fu_415_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state13))) begin
        if ((trunc_ln140_fu_428_p1 == 3'd0)) begin
            ap_phi_mux_phi_ln152_phi_fu_290_p8 = psum_0_01_reg_264;
        end else if ((1'b1 == ap_condition_514)) begin
            ap_phi_mux_phi_ln152_phi_fu_290_p8 = psum_6_07_reg_192;
        end else if ((trunc_ln140_fu_428_p1 == 3'd4)) begin
            ap_phi_mux_phi_ln152_phi_fu_290_p8 = psum_4_05_reg_216;
        end else if ((trunc_ln140_fu_428_p1 == 3'd2)) begin
            ap_phi_mux_phi_ln152_phi_fu_290_p8 = psum_2_03_reg_240;
        end else begin
            ap_phi_mux_phi_ln152_phi_fu_290_p8 = 'bx;
        end
    end else begin
        ap_phi_mux_phi_ln152_phi_fu_290_p8 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0) & (icmp_ln132_reg_492 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_x_phi_fu_172_p4 = add_ln132_reg_546;
    end else begin
        ap_phi_mux_x_phi_fu_172_p4 = x_reg_168;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state14)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_305_p0 = ap_phi_mux_psum_6_07_phi_fu_196_p4;
    end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_305_p0 = ap_phi_mux_psum_4_05_phi_fu_220_p4;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
        grp_fu_305_p0 = ap_phi_mux_psum_2_03_phi_fu_244_p4;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
        grp_fu_305_p0 = grp_fu_305_p2;
    end else begin
        grp_fu_305_p0 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_305_p1 = accum_in_0_load_70_reg_571;
    end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_305_p1 = accum_in_0_load_68_reg_551;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
        grp_fu_305_p1 = accum_in_0_load_66_reg_526;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
        grp_fu_305_p1 = accum_in_0_load_reg_506;
    end else begin
        grp_fu_305_p1 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_310_p0 = ap_phi_mux_psum_7_08_phi_fu_184_p4;
    end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_310_p0 = ap_phi_mux_psum_5_06_phi_fu_208_p4;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
        grp_fu_310_p0 = ap_phi_mux_psum_3_04_phi_fu_232_p4;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
        grp_fu_310_p0 = grp_fu_310_p2;
    end else begin
        grp_fu_310_p0 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_310_p1 = accum_in_0_load_71_reg_576;
    end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_310_p1 = accum_in_0_load_69_reg_556;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
        grp_fu_310_p1 = accum_in_0_load_67_reg_531;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
        grp_fu_310_p1 = accum_in_0_load_65_reg_511;
    end else begin
        grp_fu_310_p1 = 'bx;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_pp0_stage1 : begin
            if ((~((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter2 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0)) & (1'b0 == ap_block_pp0_stage1_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage2;
            end else if (((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter2 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
                ap_NS_fsm = ap_ST_fsm_state12;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end
        end
        ap_ST_fsm_pp0_stage2 : begin
            if ((~((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2_subdone) & (icmp_ln132_reg_492 == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b0)) & (1'b0 == ap_block_pp0_stage2_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage3;
            end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2_subdone) & (icmp_ln132_reg_492 == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
                ap_NS_fsm = ap_ST_fsm_state12;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage2;
            end
        end
        ap_ST_fsm_pp0_stage3 : begin
            if ((1'b0 == ap_block_pp0_stage3_subdone)) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage3;
            end
        end
        ap_ST_fsm_state12 : begin
            ap_NS_fsm = ap_ST_fsm_state13;
        end
        ap_ST_fsm_state13 : begin
            if (((tmp_fu_415_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state13))) begin
                ap_NS_fsm = ap_ST_fsm_state13;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state14;
            end
        end
        ap_ST_fsm_state14 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign accum_out_address0 = zext_ln140_3_fu_444_p1;

assign accum_out_address1 = zext_ln140_fu_423_p1;

assign accum_out_d0 = ((icmp_ln152_6_fu_477_p2[0:0] == 1'b1) ? psum_5_06_reg_204 : select_ln152_5_fu_469_p3);

assign accum_out_d1 = ap_phi_mux_phi_ln152_phi_fu_290_p8;

assign add_ln132_fu_387_p2 = (x_reg_168 + 10'd8);

assign add_ln140_fu_432_p2 = (q_reg_276 + 4'd2);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_pp0_stage1 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_pp0_stage2 = ap_CS_fsm[32'd3];

assign ap_CS_fsm_pp0_stage3 = ap_CS_fsm[32'd4];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state12 = ap_CS_fsm[32'd5];

assign ap_CS_fsm_state13 = ap_CS_fsm[32'd6];

assign ap_CS_fsm_state14 = ap_CS_fsm[32'd7];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1_subdone = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage2 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage2_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage2_subdone = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage3 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage3_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage3_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((ap_done_reg == 1'b1) | (ap_start == 1'b0));
end

assign ap_block_state10_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state11_pp0_stage1_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage1_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage2_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage3_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage1_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage2_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state9_pp0_stage3_iter1 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_condition_514 = (~(trunc_ln140_fu_428_p1 == 3'd0) & ~(trunc_ln140_fu_428_p1 == 3'd4) & ~(trunc_ln140_fu_428_p1 == 3'd2));
end

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign ap_phi_mux_psum_2_03_phi_fu_244_p4 = grp_fu_305_p2;

assign ap_phi_mux_psum_3_04_phi_fu_232_p4 = grp_fu_310_p2;

assign ap_phi_mux_psum_4_05_phi_fu_220_p4 = grp_fu_305_p2;

assign ap_phi_mux_psum_5_06_phi_fu_208_p4 = grp_fu_310_p2;

assign ap_phi_mux_psum_6_07_phi_fu_196_p4 = grp_fu_305_p2;

assign ap_phi_mux_psum_7_08_phi_fu_184_p4 = grp_fu_310_p2;

assign icmp_ln132_fu_321_p2 = ((ap_phi_mux_x_phi_fu_172_p4 < 10'd576) ? 1'b1 : 1'b0);

assign icmp_ln152_5_fu_463_p2 = ((or_ln140_fu_438_p2 == 3'd3) ? 1'b1 : 1'b0);

assign icmp_ln152_6_fu_477_p2 = ((or_ln140_fu_438_p2 == 3'd5) ? 1'b1 : 1'b0);

assign icmp_ln152_fu_449_p2 = ((or_ln140_fu_438_p2 == 3'd1) ? 1'b1 : 1'b0);

assign or_ln136_13_fu_343_p2 = (x_reg_168 | 10'd2);

assign or_ln136_14_fu_354_p2 = (x_reg_168 | 10'd3);

assign or_ln136_15_fu_365_p2 = (x_reg_168 | 10'd4);

assign or_ln136_16_fu_376_p2 = (x_reg_168 | 10'd5);

assign or_ln136_17_fu_393_p2 = (x_reg_168 | 10'd6);

assign or_ln136_18_fu_404_p2 = (x_reg_168 | 10'd7);

assign or_ln136_fu_332_p2 = (ap_phi_mux_x_phi_fu_172_p4 | 10'd1);

assign or_ln140_fu_438_p2 = (trunc_ln140_fu_428_p1 | 3'd1);

assign select_ln152_5_fu_469_p3 = ((icmp_ln152_5_fu_463_p2[0:0] == 1'b1) ? psum_3_04_reg_228 : select_ln152_fu_455_p3);

assign select_ln152_fu_455_p3 = ((icmp_ln152_fu_449_p2[0:0] == 1'b1) ? psum_1_02_reg_252 : psum_7_08_reg_180);

assign tmp_fu_415_p3 = q_reg_276[32'd3];

assign trunc_ln140_fu_428_p1 = q_reg_276[2:0];

assign zext_ln132_fu_327_p1 = ap_phi_mux_x_phi_fu_172_p4;

assign zext_ln136_13_fu_349_p1 = or_ln136_13_fu_343_p2;

assign zext_ln136_14_fu_360_p1 = or_ln136_14_fu_354_p2;

assign zext_ln136_15_fu_371_p1 = or_ln136_15_fu_365_p2;

assign zext_ln136_16_fu_382_p1 = or_ln136_16_fu_376_p2;

assign zext_ln136_17_fu_399_p1 = or_ln136_17_fu_393_p2;

assign zext_ln136_18_fu_410_p1 = or_ln136_18_fu_404_p2;

assign zext_ln136_fu_338_p1 = or_ln136_fu_332_p2;

assign zext_ln140_3_fu_444_p1 = or_ln140_fu_438_p2;

assign zext_ln140_fu_423_p1 = q_reg_276;

endmodule //td_fused_top_tdf11_accum_1
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf11_accum_2 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        accum_in_22,
        accum_in_22_ap_vld,
        accum_in_address0,
        accum_in_ce0,
        accum_in_q0
);

parameter    ap_ST_fsm_state1 = 7'd1;
parameter    ap_ST_fsm_state2 = 7'd2;
parameter    ap_ST_fsm_state3 = 7'd4;
parameter    ap_ST_fsm_state4 = 7'd8;
parameter    ap_ST_fsm_state5 = 7'd16;
parameter    ap_ST_fsm_state6 = 7'd32;
parameter    ap_ST_fsm_state7 = 7'd64;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [15:0] accum_in_22;
output   accum_in_22_ap_vld;
output  [2:0] accum_in_address0;
output   accum_in_ce0;
input  [15:0] accum_in_q0;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg[15:0] accum_in_22;
reg accum_in_22_ap_vld;
reg accum_in_ce0;

reg    ap_done_reg;
  reg   [6:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
wire   [3:0] add_ln164_fu_74_p2;
reg   [3:0] add_ln164_reg_91;
wire    ap_CS_fsm_state2;
wire   [0:0] icmp_ln164_fu_85_p2;
wire    ap_CS_fsm_state3;
wire   [15:0] grp_fu_68_p2;
wire    ap_CS_fsm_state7;
reg   [3:0] i_1_1_reg_44;
reg    ap_block_state1;
reg   [15:0] sum_01_reg_55;
wire   [63:0] zext_ln164_fu_80_p1;
reg   [15:0] accum_in_22_preg;
reg   [6:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 7'd1;
#0 accum_in_22_preg = 16'd0;
end

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U703(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(sum_01_reg_55),
    .din1(accum_in_q0),
    .dout(grp_fu_68_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        accum_in_22_preg <= 16'd0;
    end else begin
        if (((icmp_ln164_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
            accum_in_22_preg <= sum_01_reg_55;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if (((icmp_ln164_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        i_1_1_reg_44 <= 4'd0;
    end else if ((1'b1 == ap_CS_fsm_state7)) begin
        i_1_1_reg_44 <= add_ln164_reg_91;
    end
end

always @ (posedge ap_clk) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        sum_01_reg_55 <= 16'd0;
    end else if ((1'b1 == ap_CS_fsm_state7)) begin
        sum_01_reg_55 <= grp_fu_68_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        add_ln164_reg_91 <= add_ln164_fu_74_p2;
    end
end

always @ (*) begin
    if (((icmp_ln164_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        accum_in_22 = sum_01_reg_55;
    end else begin
        accum_in_22 = accum_in_22_preg;
    end
end

always @ (*) begin
    if (((icmp_ln164_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        accum_in_22_ap_vld = 1'b1;
    end else begin
        accum_in_22_ap_vld = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        accum_in_ce0 = 1'b1;
    end else begin
        accum_in_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln164_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln164_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_state2 : begin
            if (((icmp_ln164_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end
        end
        ap_ST_fsm_state3 : begin
            ap_NS_fsm = ap_ST_fsm_state4;
        end
        ap_ST_fsm_state4 : begin
            ap_NS_fsm = ap_ST_fsm_state5;
        end
        ap_ST_fsm_state5 : begin
            ap_NS_fsm = ap_ST_fsm_state6;
        end
        ap_ST_fsm_state6 : begin
            ap_NS_fsm = ap_ST_fsm_state7;
        end
        ap_ST_fsm_state7 : begin
            ap_NS_fsm = ap_ST_fsm_state2;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign accum_in_address0 = zext_ln164_fu_80_p1;

assign add_ln164_fu_74_p2 = (i_1_1_reg_44 + 4'd1);

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state7 = ap_CS_fsm[32'd6];

always @ (*) begin
    ap_block_state1 = ((ap_done_reg == 1'b1) | (ap_start == 1'b0));
end

assign icmp_ln164_fu_85_p2 = ((i_1_1_reg_44 == 4'd8) ? 1'b1 : 1'b0);

assign zext_ln164_fu_80_p1 = i_1_1_reg_44;

endmodule //td_fused_top_tdf11_accum_2
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf11_adjust (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        sums_read,
        adjustments_address0,
        adjustments_ce0,
        adjustments_q0,
        indices_23_dout,
        indices_23_empty_n,
        indices_23_read,
        indices_23_out_din,
        indices_23_out_full_n,
        indices_23_out_write,
        ap_return
);

parameter    ap_ST_fsm_state1 = 17'd1;
parameter    ap_ST_fsm_state2 = 17'd2;
parameter    ap_ST_fsm_state3 = 17'd4;
parameter    ap_ST_fsm_state4 = 17'd8;
parameter    ap_ST_fsm_state5 = 17'd16;
parameter    ap_ST_fsm_state6 = 17'd32;
parameter    ap_ST_fsm_state7 = 17'd64;
parameter    ap_ST_fsm_state8 = 17'd128;
parameter    ap_ST_fsm_state9 = 17'd256;
parameter    ap_ST_fsm_state10 = 17'd512;
parameter    ap_ST_fsm_state11 = 17'd1024;
parameter    ap_ST_fsm_state12 = 17'd2048;
parameter    ap_ST_fsm_state13 = 17'd4096;
parameter    ap_ST_fsm_state14 = 17'd8192;
parameter    ap_ST_fsm_state15 = 17'd16384;
parameter    ap_ST_fsm_state16 = 17'd32768;
parameter    ap_ST_fsm_state17 = 17'd65536;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
input  [15:0] sums_read;
output  [8:0] adjustments_address0;
output   adjustments_ce0;
input  [47:0] adjustments_q0;
input  [8:0] indices_23_dout;
input   indices_23_empty_n;
output   indices_23_read;
output  [8:0] indices_23_out_din;
input   indices_23_out_full_n;
output   indices_23_out_write;
output  [15:0] ap_return;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg adjustments_ce0;
reg indices_23_read;
reg indices_23_out_write;

reg    ap_done_reg;
  reg   [16:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    indices_23_blk_n;
reg    indices_23_out_blk_n;
wire    ap_CS_fsm_state4;
reg   [15:0] tmp_96_i_i_reg_179;
reg   [15:0] tmp_97_i_i_reg_184;
wire   [15:0] grp_fu_93_p2;
reg   [15:0] sub_i_i_i_reg_189;
wire    ap_CS_fsm_state8;
wire    ap_CS_fsm_state9;
wire   [15:0] grp_fu_98_p2;
reg   [15:0] mul_i_i_i_reg_199;
wire    ap_CS_fsm_state12;
wire    ap_CS_fsm_state13;
wire   [63:0] zext_ln220_fu_102_p1;
reg    ap_block_state1;
wire    ap_CS_fsm_state2;
wire    ap_CS_fsm_state3;
wire   [15:0] grp_fu_89_p1;
wire   [15:0] grp_fu_93_p1;
wire   [15:0] grp_fu_98_p1;
wire   [15:0] trunc_ln220_fu_107_p1;
wire   [15:0] grp_fu_89_p2;
wire    ap_CS_fsm_state17;
wire   [15:0] bitcast_ln648_fu_144_p1;
wire   [0:0] tmp_fu_148_p3;
reg   [16:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 17'd1;
end

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U707(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(mul_i_i_i_reg_199),
    .din1(grp_fu_89_p1),
    .dout(grp_fu_89_p2)
);

td_fused_top_hsub_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hsub_16ns_16ns_16_5_full_dsp_1_U708(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(sums_read),
    .din1(grp_fu_93_p1),
    .dout(grp_fu_93_p2)
);

td_fused_top_hmul_16ns_16ns_16_4_max_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hmul_16ns_16ns_16_4_max_dsp_1_U709(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(sub_i_i_i_reg_189),
    .din1(grp_fu_98_p1),
    .dout(grp_fu_98_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state17)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state12)) begin
        mul_i_i_i_reg_199 <= grp_fu_98_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state8)) begin
        sub_i_i_i_reg_189 <= grp_fu_93_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        tmp_96_i_i_reg_179 <= {{adjustments_q0[31:16]}};
        tmp_97_i_i_reg_184 <= {{adjustments_q0[47:32]}};
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state2) | (~((indices_23_out_full_n == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1)))) begin
        adjustments_ce0 = 1'b1;
    end else begin
        adjustments_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state17)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state17)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_23_blk_n = indices_23_empty_n;
    end else begin
        indices_23_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_23_out_blk_n = indices_23_out_full_n;
    end else begin
        indices_23_out_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((indices_23_out_full_n == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_23_out_write = 1'b1;
    end else begin
        indices_23_out_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((indices_23_out_full_n == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_23_read = 1'b1;
    end else begin
        indices_23_read = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((indices_23_out_full_n == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_state2 : begin
            ap_NS_fsm = ap_ST_fsm_state3;
        end
        ap_ST_fsm_state3 : begin
            ap_NS_fsm = ap_ST_fsm_state4;
        end
        ap_ST_fsm_state4 : begin
            ap_NS_fsm = ap_ST_fsm_state5;
        end
        ap_ST_fsm_state5 : begin
            ap_NS_fsm = ap_ST_fsm_state6;
        end
        ap_ST_fsm_state6 : begin
            ap_NS_fsm = ap_ST_fsm_state7;
        end
        ap_ST_fsm_state7 : begin
            ap_NS_fsm = ap_ST_fsm_state8;
        end
        ap_ST_fsm_state8 : begin
            ap_NS_fsm = ap_ST_fsm_state9;
        end
        ap_ST_fsm_state9 : begin
            ap_NS_fsm = ap_ST_fsm_state10;
        end
        ap_ST_fsm_state10 : begin
            ap_NS_fsm = ap_ST_fsm_state11;
        end
        ap_ST_fsm_state11 : begin
            ap_NS_fsm = ap_ST_fsm_state12;
        end
        ap_ST_fsm_state12 : begin
            ap_NS_fsm = ap_ST_fsm_state13;
        end
        ap_ST_fsm_state13 : begin
            ap_NS_fsm = ap_ST_fsm_state14;
        end
        ap_ST_fsm_state14 : begin
            ap_NS_fsm = ap_ST_fsm_state15;
        end
        ap_ST_fsm_state15 : begin
            ap_NS_fsm = ap_ST_fsm_state16;
        end
        ap_ST_fsm_state16 : begin
            ap_NS_fsm = ap_ST_fsm_state17;
        end
        ap_ST_fsm_state17 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign adjustments_address0 = zext_ln220_fu_102_p1;

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state12 = ap_CS_fsm[32'd11];

assign ap_CS_fsm_state13 = ap_CS_fsm[32'd12];

assign ap_CS_fsm_state17 = ap_CS_fsm[32'd16];

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

assign ap_CS_fsm_state8 = ap_CS_fsm[32'd7];

assign ap_CS_fsm_state9 = ap_CS_fsm[32'd8];

always @ (*) begin
    ap_block_state1 = ((indices_23_out_full_n == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0));
end

assign ap_return = ((tmp_fu_148_p3[0:0] == 1'b1) ? 16'd0 : grp_fu_89_p2);

assign bitcast_ln648_fu_144_p1 = grp_fu_89_p2;

assign grp_fu_89_p1 = tmp_97_i_i_reg_184;

assign grp_fu_93_p1 = trunc_ln220_fu_107_p1;

assign grp_fu_98_p1 = tmp_96_i_i_reg_179;

assign indices_23_out_din = indices_23_dout;

assign tmp_fu_148_p3 = bitcast_ln648_fu_144_p1[32'd15];

assign trunc_ln220_fu_107_p1 = adjustments_q0[15:0];

assign zext_ln220_fu_102_p1 = indices_23_dout;

endmodule //td_fused_top_tdf11_adjust
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf11_dot_product (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        ifmap_vec_address0,
        ifmap_vec_ce0,
        ifmap_vec_q0,
        weight_vecs_0_address0,
        weight_vecs_0_ce0,
        weight_vecs_0_q0,
        products_0_address0,
        products_0_ce0,
        products_0_we0,
        products_0_d0
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state10 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [9:0] ifmap_vec_address0;
output   ifmap_vec_ce0;
input  [15:0] ifmap_vec_q0;
output  [9:0] weight_vecs_0_address0;
output   weight_vecs_0_ce0;
input  [15:0] weight_vecs_0_q0;
output  [9:0] products_0_address0;
output   products_0_ce0;
output   products_0_we0;
output  [15:0] products_0_d0;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg ifmap_vec_ce0;
reg weight_vecs_0_ce0;
reg products_0_ce0;
reg products_0_we0;

reg    ap_done_reg;
  reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg   [9:0] indvar_flatten17_reg_97;
reg   [8:0] indvar_flatten_reg_108;
reg   [1:0] jj_reg_119;
reg   [6:0] ic_reg_131;
reg   [1:0] ii_reg_142;
wire   [9:0] add_ln147_7_fu_157_p2;
wire    ap_CS_fsm_pp0_stage0;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
wire    ap_block_state4_pp0_stage0_iter2;
wire    ap_block_state5_pp0_stage0_iter3;
wire    ap_block_state6_pp0_stage0_iter4;
wire    ap_block_state7_pp0_stage0_iter5;
wire    ap_block_state8_pp0_stage0_iter6;
wire    ap_block_state9_pp0_stage0_iter7;
wire    ap_block_pp0_stage0_11001;
wire   [0:0] icmp_ln147_fu_163_p2;
reg   [0:0] icmp_ln147_reg_408;
reg   [0:0] icmp_ln147_reg_408_pp0_iter1_reg;
reg   [0:0] icmp_ln147_reg_408_pp0_iter2_reg;
reg   [0:0] icmp_ln147_reg_408_pp0_iter3_reg;
reg   [0:0] icmp_ln147_reg_408_pp0_iter4_reg;
reg   [0:0] icmp_ln147_reg_408_pp0_iter5_reg;
reg   [0:0] icmp_ln147_reg_408_pp0_iter6_reg;
wire   [0:0] icmp_ln148_fu_169_p2;
reg   [0:0] icmp_ln148_reg_412;
wire   [0:0] and_ln147_fu_195_p2;
reg   [0:0] and_ln147_reg_419;
wire   [1:0] add_ln148_fu_201_p2;
reg   [1:0] add_ln148_reg_424;
wire   [6:0] select_ln148_fu_213_p3;
reg   [6:0] select_ln148_reg_429;
wire   [1:0] select_ln148_19_fu_221_p3;
reg   [1:0] select_ln148_19_reg_434;
wire   [5:0] trunc_ln150_fu_229_p1;
reg   [5:0] trunc_ln150_reg_440;
reg   [5:0] trunc_ln150_reg_440_pp0_iter1_reg;
reg   [5:0] trunc_ln150_reg_440_pp0_iter2_reg;
reg   [5:0] trunc_ln150_reg_440_pp0_iter3_reg;
reg   [5:0] trunc_ln150_reg_440_pp0_iter4_reg;
reg   [5:0] trunc_ln150_reg_440_pp0_iter5_reg;
reg   [5:0] trunc_ln150_reg_440_pp0_iter6_reg;
wire   [6:0] add_ln149_fu_233_p2;
wire   [8:0] select_ln148_21_fu_245_p3;
wire   [1:0] select_ln147_20_fu_287_p3;
reg   [1:0] select_ln147_20_reg_455;
reg    ap_enable_reg_pp0_iter1;
wire   [3:0] select_ln148_20_fu_370_p3;
reg   [3:0] select_ln148_20_reg_460;
reg   [3:0] select_ln148_20_reg_460_pp0_iter2_reg;
reg   [3:0] select_ln148_20_reg_460_pp0_iter3_reg;
reg   [3:0] select_ln148_20_reg_460_pp0_iter4_reg;
reg   [3:0] select_ln148_20_reg_460_pp0_iter5_reg;
reg   [3:0] select_ln148_20_reg_460_pp0_iter6_reg;
reg   [15:0] ifmap_vec_load_reg_475;
reg   [15:0] weight_vecs_0_load_reg_480;
wire   [15:0] grp_fu_153_p2;
reg   [15:0] mul_reg_485;
reg    ap_block_state1;
wire    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_flush_enable;
reg    ap_enable_reg_pp0_iter2;
reg    ap_condition_pp0_exit_iter1_state3;
reg    ap_enable_reg_pp0_iter3;
reg    ap_enable_reg_pp0_iter4;
reg    ap_enable_reg_pp0_iter5;
reg    ap_enable_reg_pp0_iter6;
reg    ap_enable_reg_pp0_iter7;
reg   [1:0] ap_phi_mux_jj_phi_fu_123_p4;
wire    ap_block_pp0_stage0;
reg   [1:0] ap_phi_mux_ii_phi_fu_146_p4;
wire   [63:0] p_cast25_fu_386_p1;
wire   [63:0] idxprom30_fu_398_p1;
wire   [0:0] icmp_ln149_fu_189_p2;
wire   [0:0] xor_ln147_fu_183_p2;
wire   [1:0] select_ln147_fu_175_p3;
wire   [0:0] or_ln148_fu_207_p2;
wire   [8:0] add_ln148_7_fu_239_p2;
wire   [3:0] shl_ln_fu_257_p3;
wire   [3:0] zext_ln150_fu_253_p1;
wire   [3:0] sub_ln150_fu_265_p2;
wire   [3:0] zext_ln150_10_fu_271_p1;
wire   [1:0] add_ln147_fu_281_p2;
wire   [3:0] tmp_fu_298_p3;
wire   [3:0] select_ln147_26_cast_fu_294_p1;
wire   [3:0] shl_ln150_mid1_fu_316_p3;
wire   [3:0] zext_ln150_15_fu_312_p1;
wire   [3:0] sub_ln150_9_fu_324_p2;
wire   [3:0] add_ln150_fu_275_p2;
wire   [3:0] empty_139_fu_306_p2;
wire   [3:0] select_ln148_25_cast_fu_344_p1;
wire   [3:0] empty_140_fu_347_p2;
wire   [3:0] select_ln147_21_fu_330_p3;
wire   [3:0] zext_ln150_16_fu_361_p1;
wire   [3:0] add_ln150_8_fu_364_p2;
wire   [3:0] select_ln147_22_fu_337_p3;
wire   [9:0] tmp_178_cast_fu_353_p3;
wire   [9:0] select_ln148_cast_fu_377_p1;
wire   [9:0] empty_141_fu_380_p2;
wire   [9:0] p_fu_392_p3;
wire    ap_CS_fsm_state10;
reg   [2:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
#0 ap_enable_reg_pp0_iter4 = 1'b0;
#0 ap_enable_reg_pp0_iter5 = 1'b0;
#0 ap_enable_reg_pp0_iter6 = 1'b0;
#0 ap_enable_reg_pp0_iter7 = 1'b0;
end

td_fused_top_hmul_16ns_16ns_16_4_max_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hmul_16ns_16ns_16_4_max_dsp_1_U695(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(ifmap_vec_load_reg_475),
    .din1(weight_vecs_0_load_reg_480),
    .dout(grp_fu_153_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state10)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if ((1'b1 == ap_condition_pp0_flush_enable)) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            if ((1'b1 == ap_condition_pp0_exit_iter1_state3)) begin
                ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter0;
            end else if ((1'b1 == 1'b1)) begin
                ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
            end
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter4 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter5 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter5 <= ap_enable_reg_pp0_iter4;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter6 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter6 <= ap_enable_reg_pp0_iter5;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter7 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter7 <= ap_enable_reg_pp0_iter6;
        end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter7 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_fu_163_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ic_reg_131 <= add_ln149_fu_233_p2;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ic_reg_131 <= 7'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_reg_408_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        ii_reg_142 <= select_ln147_20_reg_455;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ii_reg_142 <= 2'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_fu_163_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        indvar_flatten17_reg_97 <= add_ln147_7_fu_157_p2;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indvar_flatten17_reg_97 <= 10'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_fu_163_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        indvar_flatten_reg_108 <= select_ln148_21_fu_245_p3;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indvar_flatten_reg_108 <= 9'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_reg_408 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        jj_reg_119 <= select_ln148_19_reg_434;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        jj_reg_119 <= 2'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_fu_163_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        add_ln148_reg_424 <= add_ln148_fu_201_p2;
        and_ln147_reg_419 <= and_ln147_fu_195_p2;
        icmp_ln148_reg_412 <= icmp_ln148_fu_169_p2;
        select_ln148_reg_429 <= select_ln148_fu_213_p3;
        trunc_ln150_reg_440 <= trunc_ln150_fu_229_p1;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln147_reg_408 <= icmp_ln147_fu_163_p2;
        icmp_ln147_reg_408_pp0_iter1_reg <= icmp_ln147_reg_408;
        trunc_ln150_reg_440_pp0_iter1_reg <= trunc_ln150_reg_440;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        icmp_ln147_reg_408_pp0_iter2_reg <= icmp_ln147_reg_408_pp0_iter1_reg;
        icmp_ln147_reg_408_pp0_iter3_reg <= icmp_ln147_reg_408_pp0_iter2_reg;
        icmp_ln147_reg_408_pp0_iter4_reg <= icmp_ln147_reg_408_pp0_iter3_reg;
        icmp_ln147_reg_408_pp0_iter5_reg <= icmp_ln147_reg_408_pp0_iter4_reg;
        icmp_ln147_reg_408_pp0_iter6_reg <= icmp_ln147_reg_408_pp0_iter5_reg;
        select_ln148_20_reg_460_pp0_iter2_reg <= select_ln148_20_reg_460;
        select_ln148_20_reg_460_pp0_iter3_reg <= select_ln148_20_reg_460_pp0_iter2_reg;
        select_ln148_20_reg_460_pp0_iter4_reg <= select_ln148_20_reg_460_pp0_iter3_reg;
        select_ln148_20_reg_460_pp0_iter5_reg <= select_ln148_20_reg_460_pp0_iter4_reg;
        select_ln148_20_reg_460_pp0_iter6_reg <= select_ln148_20_reg_460_pp0_iter5_reg;
        trunc_ln150_reg_440_pp0_iter2_reg <= trunc_ln150_reg_440_pp0_iter1_reg;
        trunc_ln150_reg_440_pp0_iter3_reg <= trunc_ln150_reg_440_pp0_iter2_reg;
        trunc_ln150_reg_440_pp0_iter4_reg <= trunc_ln150_reg_440_pp0_iter3_reg;
        trunc_ln150_reg_440_pp0_iter5_reg <= trunc_ln150_reg_440_pp0_iter4_reg;
        trunc_ln150_reg_440_pp0_iter6_reg <= trunc_ln150_reg_440_pp0_iter5_reg;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_reg_408_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        ifmap_vec_load_reg_475 <= ifmap_vec_q0;
        weight_vecs_0_load_reg_480 <= weight_vecs_0_q0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_reg_408_pp0_iter5_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        mul_reg_485 <= grp_fu_153_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_reg_408 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        select_ln147_20_reg_455 <= select_ln147_20_fu_287_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_fu_163_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        select_ln148_19_reg_434 <= select_ln148_19_fu_221_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_reg_408 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        select_ln148_20_reg_460 <= select_ln148_20_fu_370_p3;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_condition_pp0_exit_iter1_state3 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter1_state3 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln147_fu_163_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_condition_pp0_flush_enable = 1'b1;
    end else begin
        ap_condition_pp0_flush_enable = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state10)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter7 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln147_reg_408_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        ap_phi_mux_ii_phi_fu_146_p4 = select_ln147_20_reg_455;
    end else begin
        ap_phi_mux_ii_phi_fu_146_p4 = ii_reg_142;
    end
end

always @ (*) begin
    if (((icmp_ln147_reg_408 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_jj_phi_fu_123_p4 = select_ln148_19_reg_434;
    end else begin
        ap_phi_mux_jj_phi_fu_123_p4 = jj_reg_119;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state10)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ifmap_vec_ce0 = 1'b1;
    end else begin
        ifmap_vec_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter7 == 1'b1))) begin
        products_0_ce0 = 1'b1;
    end else begin
        products_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln147_reg_408_pp0_iter6_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter7 == 1'b1))) begin
        products_0_we0 = 1'b1;
    end else begin
        products_0_we0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        weight_vecs_0_ce0 = 1'b1;
    end else begin
        weight_vecs_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((~((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b1)) & ~((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter7 == 1'b1) & (ap_enable_reg_pp0_iter6 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if ((((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter7 == 1'b1) & (ap_enable_reg_pp0_iter6 == 1'b0)) | ((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b1)))) begin
                ap_NS_fsm = ap_ST_fsm_state10;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state10 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln147_7_fu_157_p2 = (indvar_flatten17_reg_97 + 10'd1);

assign add_ln147_fu_281_p2 = (ap_phi_mux_ii_phi_fu_146_p4 + 2'd1);

assign add_ln148_7_fu_239_p2 = (indvar_flatten_reg_108 + 9'd1);

assign add_ln148_fu_201_p2 = (select_ln147_fu_175_p3 + 2'd1);

assign add_ln149_fu_233_p2 = (select_ln148_fu_213_p3 + 7'd1);

assign add_ln150_8_fu_364_p2 = (select_ln147_21_fu_330_p3 + zext_ln150_16_fu_361_p1);

assign add_ln150_fu_275_p2 = (sub_ln150_fu_265_p2 + zext_ln150_10_fu_271_p1);

assign and_ln147_fu_195_p2 = (xor_ln147_fu_183_p2 & icmp_ln149_fu_189_p2);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state10 = ap_CS_fsm[32'd2];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (ap_done_reg == 1'b1));
end

assign ap_block_state2_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter4 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage0_iter5 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage0_iter6 = ~(1'b1 == 1'b1);

assign ap_block_state9_pp0_stage0_iter7 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign empty_139_fu_306_p2 = (tmp_fu_298_p3 - select_ln147_26_cast_fu_294_p1);

assign empty_140_fu_347_p2 = (empty_139_fu_306_p2 + select_ln148_25_cast_fu_344_p1);

assign empty_141_fu_380_p2 = (tmp_178_cast_fu_353_p3 + select_ln148_cast_fu_377_p1);

assign icmp_ln147_fu_163_p2 = ((indvar_flatten17_reg_97 == 10'd576) ? 1'b1 : 1'b0);

assign icmp_ln148_fu_169_p2 = ((indvar_flatten_reg_108 == 9'd192) ? 1'b1 : 1'b0);

assign icmp_ln149_fu_189_p2 = ((ic_reg_131 == 7'd64) ? 1'b1 : 1'b0);

assign idxprom30_fu_398_p1 = p_fu_392_p3;

assign ifmap_vec_address0 = p_cast25_fu_386_p1;

assign or_ln148_fu_207_p2 = (icmp_ln148_fu_169_p2 | and_ln147_fu_195_p2);

assign p_cast25_fu_386_p1 = empty_141_fu_380_p2;

assign p_fu_392_p3 = {{select_ln148_20_reg_460_pp0_iter6_reg}, {trunc_ln150_reg_440_pp0_iter6_reg}};

assign products_0_address0 = idxprom30_fu_398_p1;

assign products_0_d0 = mul_reg_485;

assign select_ln147_20_fu_287_p3 = ((icmp_ln148_reg_412[0:0] == 1'b1) ? add_ln147_fu_281_p2 : ap_phi_mux_ii_phi_fu_146_p4);

assign select_ln147_21_fu_330_p3 = ((icmp_ln148_reg_412[0:0] == 1'b1) ? sub_ln150_9_fu_324_p2 : sub_ln150_fu_265_p2);

assign select_ln147_22_fu_337_p3 = ((icmp_ln148_reg_412[0:0] == 1'b1) ? sub_ln150_9_fu_324_p2 : add_ln150_fu_275_p2);

assign select_ln147_26_cast_fu_294_p1 = select_ln147_20_fu_287_p3;

assign select_ln147_fu_175_p3 = ((icmp_ln148_fu_169_p2[0:0] == 1'b1) ? 2'd0 : ap_phi_mux_jj_phi_fu_123_p4);

assign select_ln148_19_fu_221_p3 = ((and_ln147_fu_195_p2[0:0] == 1'b1) ? add_ln148_fu_201_p2 : select_ln147_fu_175_p3);

assign select_ln148_20_fu_370_p3 = ((and_ln147_reg_419[0:0] == 1'b1) ? add_ln150_8_fu_364_p2 : select_ln147_22_fu_337_p3);

assign select_ln148_21_fu_245_p3 = ((icmp_ln148_fu_169_p2[0:0] == 1'b1) ? 9'd1 : add_ln148_7_fu_239_p2);

assign select_ln148_25_cast_fu_344_p1 = select_ln148_19_reg_434;

assign select_ln148_cast_fu_377_p1 = select_ln148_reg_429;

assign select_ln148_fu_213_p3 = ((or_ln148_fu_207_p2[0:0] == 1'b1) ? 7'd0 : ic_reg_131);

assign shl_ln150_mid1_fu_316_p3 = {{add_ln147_fu_281_p2}, {2'd0}};

assign shl_ln_fu_257_p3 = {{ap_phi_mux_ii_phi_fu_146_p4}, {2'd0}};

assign sub_ln150_9_fu_324_p2 = (shl_ln150_mid1_fu_316_p3 - zext_ln150_15_fu_312_p1);

assign sub_ln150_fu_265_p2 = (shl_ln_fu_257_p3 - zext_ln150_fu_253_p1);

assign tmp_178_cast_fu_353_p3 = {{empty_140_fu_347_p2}, {6'd0}};

assign tmp_fu_298_p3 = {{select_ln147_20_fu_287_p3}, {2'd0}};

assign trunc_ln150_fu_229_p1 = select_ln148_fu_213_p3[5:0];

assign weight_vecs_0_address0 = p_cast25_fu_386_p1;

assign xor_ln147_fu_183_p2 = (icmp_ln148_fu_169_p2 ^ 1'd1);

assign zext_ln150_10_fu_271_p1 = jj_reg_119;

assign zext_ln150_15_fu_312_p1 = add_ln147_fu_281_p2;

assign zext_ln150_16_fu_361_p1 = add_ln148_reg_424;

assign zext_ln150_fu_253_p1 = ap_phi_mux_ii_phi_fu_146_p4;

endmodule //td_fused_top_tdf11_dot_product
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf11_get_next_ijk (
        ap_clk,
        ap_rst,
        ap_start,
        start_full_n,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        start_out,
        start_write,
        indices_0_din,
        indices_0_full_n,
        indices_0_write,
        indices_1_din,
        indices_1_full_n,
        indices_1_write,
        indices_2_out_din,
        indices_2_out_full_n,
        indices_2_out_write,
        indices_2_out1_din,
        indices_2_out1_full_n,
        indices_2_out1_write,
        write_r_din,
        write_r_full_n,
        write_r_write
);

parameter    ap_ST_fsm_state1 = 1'd1;

input   ap_clk;
input   ap_rst;
input   ap_start;
input   start_full_n;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output   start_out;
output   start_write;
output  [15:0] indices_0_din;
input   indices_0_full_n;
output   indices_0_write;
output  [15:0] indices_1_din;
input   indices_1_full_n;
output   indices_1_write;
output  [8:0] indices_2_out_din;
input   indices_2_out_full_n;
output   indices_2_out_write;
output  [8:0] indices_2_out1_din;
input   indices_2_out1_full_n;
output   indices_2_out1_write;
output   write_r_din;
input   write_r_full_n;
output   write_r_write;

reg ap_done;
reg ap_idle;
reg start_write;
reg indices_0_write;
reg indices_1_write;
reg indices_2_out_write;
reg indices_2_out1_write;
reg write_r_write;

reg    real_start;
reg    start_once_reg;
reg    ap_done_reg;
  reg   [0:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    internal_ap_ready;
reg   [15:0] i_9;
reg   [15:0] j_9;
reg   [15:0] k_9;
reg    indices_0_blk_n;
reg    indices_1_blk_n;
reg    indices_2_out_blk_n;
reg    indices_2_out1_blk_n;
reg    write_r_blk_n;
reg   [0:0] ap_phi_mux_j_20_flag_0_i_phi_fu_90_p6;
reg    ap_block_state1;
wire   [0:0] icmp_ln188_fu_161_p2;
wire   [0:0] icmp_ln191_fu_174_p2;
reg   [15:0] ap_phi_mux_j_20_new_0_i_phi_fu_104_p6;
wire   [15:0] add_ln190_fu_167_p2;
reg   [15:0] ap_phi_mux_k_20_new_0_i_phi_fu_117_p6;
wire   [15:0] add_ln187_fu_154_p2;
wire   [15:0] select_ln194_fu_192_p3;
wire   [8:0] trunc_ln185_fu_141_p1;
wire   [15:0] add_ln193_fu_180_p2;
wire   [0:0] icmp_ln194_fu_186_p2;
reg   [0:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 start_once_reg = 1'b0;
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 1'd1;
#0 i_9 = 16'd0;
#0 j_9 = 16'd0;
#0 k_9 = 16'd0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((~((real_start == 1'b0) | (write_r_full_n == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        start_once_reg <= 1'b0;
    end else begin
        if (((real_start == 1'b1) & (internal_ap_ready == 1'b0))) begin
            start_once_reg <= 1'b1;
        end else if ((internal_ap_ready == 1'b1)) begin
            start_once_reg <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((~((real_start == 1'b0) | (write_r_full_n == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (icmp_ln191_fu_174_p2 == 1'd1) & (icmp_ln188_fu_161_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1))) begin
        i_9 <= select_ln194_fu_192_p3;
    end
end

always @ (posedge ap_clk) begin
    if ((~((real_start == 1'b0) | (write_r_full_n == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (ap_phi_mux_j_20_flag_0_i_phi_fu_90_p6 == 1'd1) & (1'b1 == ap_CS_fsm_state1))) begin
        j_9 <= ap_phi_mux_j_20_new_0_i_phi_fu_104_p6;
    end
end

always @ (posedge ap_clk) begin
    if ((~((real_start == 1'b0) | (write_r_full_n == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        k_9 <= ap_phi_mux_k_20_new_0_i_phi_fu_117_p6;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (write_r_full_n == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((real_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln188_fu_161_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_phi_mux_j_20_flag_0_i_phi_fu_90_p6 = 1'd0;
    end else if ((((icmp_ln191_fu_174_p2 == 1'd0) & (icmp_ln188_fu_161_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1)) | ((icmp_ln191_fu_174_p2 == 1'd1) & (icmp_ln188_fu_161_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1)))) begin
        ap_phi_mux_j_20_flag_0_i_phi_fu_90_p6 = 1'd1;
    end else begin
        ap_phi_mux_j_20_flag_0_i_phi_fu_90_p6 = 'bx;
    end
end

always @ (*) begin
    if (((icmp_ln188_fu_161_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1))) begin
        if ((icmp_ln191_fu_174_p2 == 1'd0)) begin
            ap_phi_mux_j_20_new_0_i_phi_fu_104_p6 = add_ln190_fu_167_p2;
        end else if ((icmp_ln191_fu_174_p2 == 1'd1)) begin
            ap_phi_mux_j_20_new_0_i_phi_fu_104_p6 = 16'd0;
        end else begin
            ap_phi_mux_j_20_new_0_i_phi_fu_104_p6 = 'bx;
        end
    end else begin
        ap_phi_mux_j_20_new_0_i_phi_fu_104_p6 = 'bx;
    end
end

always @ (*) begin
    if (((icmp_ln188_fu_161_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_phi_mux_k_20_new_0_i_phi_fu_117_p6 = add_ln187_fu_154_p2;
    end else if ((((icmp_ln191_fu_174_p2 == 1'd0) & (icmp_ln188_fu_161_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1)) | ((icmp_ln191_fu_174_p2 == 1'd1) & (icmp_ln188_fu_161_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1)))) begin
        ap_phi_mux_k_20_new_0_i_phi_fu_117_p6 = 16'd0;
    end else begin
        ap_phi_mux_k_20_new_0_i_phi_fu_117_p6 = 'bx;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_0_blk_n = indices_0_full_n;
    end else begin
        indices_0_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (write_r_full_n == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_0_write = 1'b1;
    end else begin
        indices_0_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_1_blk_n = indices_1_full_n;
    end else begin
        indices_1_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (write_r_full_n == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_1_write = 1'b1;
    end else begin
        indices_1_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_2_out1_blk_n = indices_2_out1_full_n;
    end else begin
        indices_2_out1_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (write_r_full_n == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_2_out1_write = 1'b1;
    end else begin
        indices_2_out1_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_2_out_blk_n = indices_2_out_full_n;
    end else begin
        indices_2_out_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (write_r_full_n == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_2_out_write = 1'b1;
    end else begin
        indices_2_out_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (write_r_full_n == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        internal_ap_ready = 1'b1;
    end else begin
        internal_ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((start_full_n == 1'b0) & (start_once_reg == 1'b0))) begin
        real_start = 1'b0;
    end else begin
        real_start = ap_start;
    end
end

always @ (*) begin
    if (((real_start == 1'b1) & (start_once_reg == 1'b0))) begin
        start_write = 1'b1;
    end else begin
        start_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        write_r_blk_n = write_r_full_n;
    end else begin
        write_r_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (write_r_full_n == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        write_r_write = 1'b1;
    end else begin
        write_r_write = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln187_fu_154_p2 = (k_9 + 16'd1);

assign add_ln190_fu_167_p2 = (j_9 + 16'd1);

assign add_ln193_fu_180_p2 = (i_9 + 16'd1);

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

always @ (*) begin
    ap_block_state1 = ((real_start == 1'b0) | (write_r_full_n == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1));
end

assign ap_ready = internal_ap_ready;

assign icmp_ln188_fu_161_p2 = ((add_ln187_fu_154_p2 == 16'd512) ? 1'b1 : 1'b0);

assign icmp_ln191_fu_174_p2 = ((add_ln190_fu_167_p2 == 16'd14) ? 1'b1 : 1'b0);

assign icmp_ln194_fu_186_p2 = ((add_ln193_fu_180_p2 == 16'd14) ? 1'b1 : 1'b0);

assign indices_0_din = i_9;

assign indices_1_din = j_9;

assign indices_2_out1_din = trunc_ln185_fu_141_p1;

assign indices_2_out_din = trunc_ln185_fu_141_p1;

assign select_ln194_fu_192_p3 = ((icmp_ln194_fu_186_p2[0:0] == 1'b1) ? 16'd0 : add_ln193_fu_180_p2);

assign start_out = real_start;

assign trunc_ln185_fu_141_p1 = k_9[8:0];

assign write_r_din = ((k_9 == 16'd511) ? 1'b1 : 1'b0);

endmodule //td_fused_top_tdf11_get_next_ijk
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_tdf11_l2_filters_ram (addr0, ce0, q0, addr1, ce1, d1, we1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 16;
parameter MEM_SIZE = 65536;

input[AWIDTH-1:0] addr0;
input ce0;
output wire[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
input clk;

 reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];
wire [AWIDTH-1:0] addr0_t0; 
reg [AWIDTH-1:0] addr0_t1; 
reg [DWIDTH-1:0] q0_t0;
reg [DWIDTH-1:0] q0_t1;
wire [AWIDTH-1:0] addr1_t0; 
reg [AWIDTH-1:0] addr1_t1; 
wire [DWIDTH-1:0] d1_t0; 
wire we1_t0; 
reg [DWIDTH-1:0] d1_t1; 
reg we1_t1; 


assign addr0_t0 = addr0;
assign q0 = q0_t1;
assign addr1_t0 = addr1;
assign d1_t0 = d1;
assign we1_t0 = we1;

always @(posedge clk)  
begin
    if (ce0) 
    begin
        addr0_t1 <= addr0_t0; 
        q0_t1 <= q0_t0;
    end
    if (ce1) 
    begin
        addr1_t1 <= addr1_t0; 
        d1_t1 <= d1_t0;
        we1_t1 <= we1_t0;
    end
end


always @(posedge clk)  
begin 
    if (ce0) begin
        q0_t0 <= ram[addr0_t1];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1_t1) 
            ram[addr1_t1] <= d1_t1; 
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_tdf11_l2_filters(
    reset,
    clk,
    address0,
    ce0,
    q0,
    address1,
    ce1,
    we1,
    d1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd65536;
parameter AddressWidth = 32'd16;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;



td_fused_top_tdf11_l2_filters_ram td_fused_top_tdf11_l2_filters_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 )
);

endmodule

// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf11_l2_multiply72 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        intermediate_fmaps_read,
        l2_filter_data_address0,
        l2_filter_data_ce0,
        l2_filter_data_q0,
        l2_products_address0,
        l2_products_ce0,
        l2_products_we0,
        l2_products_d0,
        indices_23_dout,
        indices_23_empty_n,
        indices_23_read
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state10 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
input  [15:0] intermediate_fmaps_read;
output  [15:0] l2_filter_data_address0;
output   l2_filter_data_ce0;
input  [15:0] l2_filter_data_q0;
output  [6:0] l2_products_address0;
output   l2_products_ce0;
output   l2_products_we0;
output  [15:0] l2_products_d0;
input  [8:0] indices_23_dout;
input   indices_23_empty_n;
output   indices_23_read;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg l2_filter_data_ce0;
reg l2_products_ce0;
reg l2_products_we0;
reg indices_23_read;

reg    ap_done_reg;
  reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    indices_23_blk_n;
reg   [7:0] i_1_1_reg_106;
reg   [7:0] i_1_1_reg_106_pp0_iter1_reg;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
wire    ap_block_state4_pp0_stage0_iter2;
wire    ap_block_state5_pp0_stage0_iter3;
wire    ap_block_state6_pp0_stage0_iter4;
wire    ap_block_state7_pp0_stage0_iter5;
wire    ap_block_state8_pp0_stage0_iter6;
wire    ap_block_state9_pp0_stage0_iter7;
wire    ap_block_pp0_stage0_11001;
reg   [7:0] i_1_1_reg_106_pp0_iter2_reg;
reg   [7:0] i_1_1_reg_106_pp0_iter3_reg;
reg   [7:0] i_1_1_reg_106_pp0_iter4_reg;
reg   [7:0] i_1_1_reg_106_pp0_iter5_reg;
reg   [7:0] i_1_1_reg_106_pp0_iter6_reg;
reg   [8:0] indices_23_read_reg_167;
wire   [7:0] i_12_fu_123_p2;
reg   [7:0] i_12_reg_172;
reg    ap_enable_reg_pp0_iter0;
wire   [0:0] icmp_ln20_fu_129_p2;
reg   [0:0] icmp_ln20_reg_177;
reg   [0:0] icmp_ln20_reg_177_pp0_iter1_reg;
reg   [0:0] icmp_ln20_reg_177_pp0_iter2_reg;
reg   [0:0] icmp_ln20_reg_177_pp0_iter3_reg;
reg   [0:0] icmp_ln20_reg_177_pp0_iter4_reg;
reg   [0:0] icmp_ln20_reg_177_pp0_iter5_reg;
reg   [0:0] icmp_ln20_reg_177_pp0_iter6_reg;
wire   [15:0] grp_fu_118_p2;
reg   [15:0] mul_i_i_reg_191;
reg    ap_block_state1;
wire    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_exit_iter0_state2;
reg    ap_enable_reg_pp0_iter1;
reg    ap_enable_reg_pp0_iter2;
reg    ap_enable_reg_pp0_iter3;
reg    ap_enable_reg_pp0_iter4;
reg    ap_enable_reg_pp0_iter5;
reg    ap_enable_reg_pp0_iter6;
reg    ap_enable_reg_pp0_iter7;
reg   [7:0] ap_phi_mux_i_1_1_phi_fu_110_p4;
wire    ap_block_pp0_stage0;
wire   [63:0] zext_ln29_25_fu_152_p1;
wire   [63:0] zext_ln29_fu_157_p1;
wire   [6:0] trunc_ln29_fu_140_p1;
wire   [8:0] l2_ichan_fu_135_p2;
wire   [15:0] tmp_s_fu_144_p3;
wire    ap_CS_fsm_state10;
reg   [2:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
#0 ap_enable_reg_pp0_iter4 = 1'b0;
#0 ap_enable_reg_pp0_iter5 = 1'b0;
#0 ap_enable_reg_pp0_iter6 = 1'b0;
#0 ap_enable_reg_pp0_iter7 = 1'b0;
end

td_fused_top_hmul_16ns_16ns_16_4_max_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hmul_16ns_16ns_16_4_max_dsp_1_U714(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(l2_filter_data_q0),
    .din1(intermediate_fmaps_read),
    .dout(grp_fu_118_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state10)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b1 == ap_condition_pp0_exit_iter0_state2))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            if ((1'b1 == ap_condition_pp0_exit_iter0_state2)) begin
                ap_enable_reg_pp0_iter1 <= (1'b1 ^ ap_condition_pp0_exit_iter0_state2);
            end else if ((1'b1 == 1'b1)) begin
                ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
            end
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter4 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter5 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter5 <= ap_enable_reg_pp0_iter4;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter6 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter6 <= ap_enable_reg_pp0_iter5;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter7 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter7 <= ap_enable_reg_pp0_iter6;
        end else if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter7 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln20_reg_177 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        i_1_1_reg_106 <= i_12_reg_172;
    end else if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        i_1_1_reg_106 <= 8'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        i_12_reg_172 <= i_12_fu_123_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        i_1_1_reg_106_pp0_iter1_reg <= i_1_1_reg_106;
        icmp_ln20_reg_177 <= icmp_ln20_fu_129_p2;
        icmp_ln20_reg_177_pp0_iter1_reg <= icmp_ln20_reg_177;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        i_1_1_reg_106_pp0_iter2_reg <= i_1_1_reg_106_pp0_iter1_reg;
        i_1_1_reg_106_pp0_iter3_reg <= i_1_1_reg_106_pp0_iter2_reg;
        i_1_1_reg_106_pp0_iter4_reg <= i_1_1_reg_106_pp0_iter3_reg;
        i_1_1_reg_106_pp0_iter5_reg <= i_1_1_reg_106_pp0_iter4_reg;
        i_1_1_reg_106_pp0_iter6_reg <= i_1_1_reg_106_pp0_iter5_reg;
        icmp_ln20_reg_177_pp0_iter2_reg <= icmp_ln20_reg_177_pp0_iter1_reg;
        icmp_ln20_reg_177_pp0_iter3_reg <= icmp_ln20_reg_177_pp0_iter2_reg;
        icmp_ln20_reg_177_pp0_iter4_reg <= icmp_ln20_reg_177_pp0_iter3_reg;
        icmp_ln20_reg_177_pp0_iter5_reg <= icmp_ln20_reg_177_pp0_iter4_reg;
        icmp_ln20_reg_177_pp0_iter6_reg <= icmp_ln20_reg_177_pp0_iter5_reg;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state1)) begin
        indices_23_read_reg_167 <= indices_23_dout;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln20_reg_177_pp0_iter5_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        mul_i_i_reg_191 <= grp_fu_118_p2;
    end
end

always @ (*) begin
    if ((icmp_ln20_fu_129_p2 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state2 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state2 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state10)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter7 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln20_reg_177 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_i_1_1_phi_fu_110_p4 = i_12_reg_172;
    end else begin
        ap_phi_mux_i_1_1_phi_fu_110_p4 = i_1_1_reg_106;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state10)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_23_blk_n = indices_23_empty_n;
    end else begin
        indices_23_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_23_read = 1'b1;
    end else begin
        indices_23_read = 1'b0;
    end
end

always @ (*) begin
    if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter3 == 1'b1)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1)))) begin
        l2_filter_data_ce0 = 1'b1;
    end else begin
        l2_filter_data_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter7 == 1'b1))) begin
        l2_products_ce0 = 1'b1;
    end else begin
        l2_products_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln20_reg_177_pp0_iter6_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter7 == 1'b1))) begin
        l2_products_we0 = 1'b1;
    end else begin
        l2_products_we0 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((~((icmp_ln20_fu_129_p2 == 1'd1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter1 == 1'b0)) & ~((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter7 == 1'b1) & (ap_enable_reg_pp0_iter6 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if ((((icmp_ln20_fu_129_p2 == 1'd1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter1 == 1'b0)) | ((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter7 == 1'b1) & (ap_enable_reg_pp0_iter6 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_state10;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state10 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state10 = ap_CS_fsm[32'd2];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1));
end

assign ap_block_state2_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter4 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage0_iter5 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage0_iter6 = ~(1'b1 == 1'b1);

assign ap_block_state9_pp0_stage0_iter7 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign i_12_fu_123_p2 = (ap_phi_mux_i_1_1_phi_fu_110_p4 + 8'd1);

assign icmp_ln20_fu_129_p2 = ((ap_phi_mux_i_1_1_phi_fu_110_p4 == 8'd128) ? 1'b1 : 1'b0);

assign l2_filter_data_address0 = zext_ln29_25_fu_152_p1;

assign l2_ichan_fu_135_p2 = (indices_23_read_reg_167 + 9'd0);

assign l2_products_address0 = zext_ln29_fu_157_p1;

assign l2_products_d0 = mul_i_i_reg_191;

assign tmp_s_fu_144_p3 = {{trunc_ln29_fu_140_p1}, {l2_ichan_fu_135_p2}};

assign trunc_ln29_fu_140_p1 = ap_phi_mux_i_1_1_phi_fu_110_p4[6:0];

assign zext_ln29_25_fu_152_p1 = tmp_s_fu_144_p3;

assign zext_ln29_fu_157_p1 = i_1_1_reg_106_pp0_iter6_reg;

endmodule //td_fused_top_tdf11_l2_multiply72
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_tdf11_l2_writeOutputs_171_running_sums_2_ram (addr0, ce0, d0, we0, addr1, ce1, q1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
input[AWIDTH-1:0] addr1;
input ce1;
output reg[DWIDTH-1:0] q1;
input clk;

 reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];

//initial begin
//    $readmemh("./td_fused_top_tdf11_l2_writeOutputs_171_running_sums_2_ram.dat", ram);
//end



always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        q1 <= ram[addr1];
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_tdf11_l2_writeOutputs_171_running_sums_2(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    address1,
    ce1,
    q1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
input[AddressWidth - 1:0] address1;
input ce1;
output[DataWidth - 1:0] q1;



td_fused_top_tdf11_l2_writeOutputs_171_running_sums_2_ram td_fused_top_tdf11_l2_writeOutputs_171_running_sums_2_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .q1( q1 )
);

endmodule

// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf11_l2_writeOutputs_171 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        indices_01_dout,
        indices_01_empty_n,
        indices_01_read,
        indices_12_dout,
        indices_12_empty_n,
        indices_12_read,
        write4_dout,
        write4_empty_n,
        write4_read,
        l2_partial_sums_address0,
        l2_partial_sums_ce0,
        l2_partial_sums_q0,
        out_data_address1,
        out_data_ce1,
        out_data_we1,
        out_data_d1,
        l2_adjustments_address0,
        l2_adjustments_ce0,
        l2_adjustments_q0
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state25 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
input  [3:0] indices_01_dout;
input   indices_01_empty_n;
output   indices_01_read;
input  [7:0] indices_12_dout;
input   indices_12_empty_n;
output   indices_12_read;
input  [0:0] write4_dout;
input   write4_empty_n;
output   write4_read;
output  [6:0] l2_partial_sums_address0;
output   l2_partial_sums_ce0;
input  [15:0] l2_partial_sums_q0;
output  [12:0] out_data_address1;
output   out_data_ce1;
output   out_data_we1;
output  [63:0] out_data_d1;
output  [6:0] l2_adjustments_address0;
output   l2_adjustments_ce0;
input  [47:0] l2_adjustments_q0;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg indices_01_read;
reg indices_12_read;
reg write4_read;
reg l2_partial_sums_ce0;
reg out_data_ce1;
reg out_data_we1;
reg l2_adjustments_ce0;

reg    ap_done_reg;
  reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    running_sums_2_ce0;
reg    running_sums_2_we0;
wire   [15:0] running_sums_2_d0;
wire   [6:0] running_sums_2_address1;
reg    running_sums_2_ce1;
wire   [15:0] running_sums_2_q1;
reg    indices_01_blk_n;
reg    indices_12_blk_n;
reg    write4_blk_n;
reg   [7:0] ochan_reg_208;
reg   [0:0] write4_read_reg_567;
wire   [9:0] add_ln109_fu_273_p2;
reg   [9:0] add_ln109_reg_573;
wire   [7:0] ochan_1_fu_279_p2;
wire    ap_CS_fsm_pp0_stage0;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
wire    ap_block_state4_pp0_stage0_iter2;
wire    ap_block_state5_pp0_stage0_iter3;
wire    ap_block_state6_pp0_stage0_iter4;
wire    ap_block_state7_pp0_stage0_iter5;
wire    ap_block_state8_pp0_stage0_iter6;
wire    ap_block_state9_pp0_stage0_iter7;
wire    ap_block_state10_pp0_stage0_iter8;
wire    ap_block_state11_pp0_stage0_iter9;
wire    ap_block_state12_pp0_stage0_iter10;
wire    ap_block_state13_pp0_stage0_iter11;
wire    ap_block_state14_pp0_stage0_iter12;
wire    ap_block_state15_pp0_stage0_iter13;
wire    ap_block_state16_pp0_stage0_iter14;
wire    ap_block_state17_pp0_stage0_iter15;
wire    ap_block_state18_pp0_stage0_iter16;
wire    ap_block_state19_pp0_stage0_iter17;
wire    ap_block_state20_pp0_stage0_iter18;
wire    ap_block_state21_pp0_stage0_iter19;
wire    ap_block_state22_pp0_stage0_iter20;
wire    ap_block_state23_pp0_stage0_iter21;
wire    ap_block_state24_pp0_stage0_iter22;
wire    ap_block_pp0_stage0_11001;
wire   [0:0] icmp_ln86_fu_285_p2;
wire   [1:0] trunc_ln86_fu_291_p1;
reg   [1:0] trunc_ln86_reg_587;
reg   [1:0] trunc_ln86_reg_587_pp0_iter1_reg;
reg   [1:0] trunc_ln86_reg_587_pp0_iter2_reg;
reg   [1:0] trunc_ln86_reg_587_pp0_iter3_reg;
reg   [1:0] trunc_ln86_reg_587_pp0_iter4_reg;
reg   [1:0] trunc_ln86_reg_587_pp0_iter5_reg;
reg   [1:0] trunc_ln86_reg_587_pp0_iter6_reg;
reg   [1:0] trunc_ln86_reg_587_pp0_iter7_reg;
reg   [1:0] trunc_ln86_reg_587_pp0_iter8_reg;
reg   [1:0] trunc_ln86_reg_587_pp0_iter9_reg;
reg   [1:0] trunc_ln86_reg_587_pp0_iter10_reg;
reg   [1:0] trunc_ln86_reg_587_pp0_iter11_reg;
reg   [1:0] trunc_ln86_reg_587_pp0_iter12_reg;
reg   [1:0] trunc_ln86_reg_587_pp0_iter13_reg;
reg   [1:0] trunc_ln86_reg_587_pp0_iter14_reg;
reg   [1:0] trunc_ln86_reg_587_pp0_iter15_reg;
reg   [1:0] trunc_ln86_reg_587_pp0_iter16_reg;
reg   [1:0] trunc_ln86_reg_587_pp0_iter17_reg;
reg   [1:0] trunc_ln86_reg_587_pp0_iter18_reg;
reg   [1:0] trunc_ln86_reg_587_pp0_iter19_reg;
reg   [1:0] trunc_ln86_reg_587_pp0_iter20_reg;
wire   [63:0] zext_ln89_fu_295_p1;
reg   [63:0] zext_ln89_reg_594;
reg   [63:0] zext_ln89_reg_594_pp0_iter1_reg;
reg   [63:0] zext_ln89_reg_594_pp0_iter2_reg;
reg   [63:0] zext_ln89_reg_594_pp0_iter3_reg;
reg   [6:0] running_sums_2_addr_reg_604;
reg   [6:0] running_sums_2_addr_reg_604_pp0_iter1_reg;
reg   [6:0] running_sums_2_addr_reg_604_pp0_iter2_reg;
reg   [6:0] running_sums_2_addr_reg_604_pp0_iter3_reg;
reg   [6:0] running_sums_2_addr_reg_604_pp0_iter4_reg;
reg   [6:0] running_sums_2_addr_reg_604_pp0_iter5_reg;
reg   [6:0] running_sums_2_addr_reg_604_pp0_iter6_reg;
wire   [0:0] and_ln103_fu_307_p2;
reg   [0:0] and_ln103_reg_610;
reg   [0:0] and_ln103_reg_610_pp0_iter1_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter2_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter3_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter4_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter5_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter6_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter7_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter8_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter9_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter10_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter11_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter12_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter13_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter14_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter15_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter16_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter17_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter18_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter19_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter20_reg;
reg   [4:0] lshr_ln_reg_614;
reg   [4:0] lshr_ln_reg_614_pp0_iter1_reg;
reg   [4:0] lshr_ln_reg_614_pp0_iter2_reg;
reg   [4:0] lshr_ln_reg_614_pp0_iter3_reg;
reg   [4:0] lshr_ln_reg_614_pp0_iter4_reg;
reg   [4:0] lshr_ln_reg_614_pp0_iter5_reg;
reg   [4:0] lshr_ln_reg_614_pp0_iter6_reg;
reg   [4:0] lshr_ln_reg_614_pp0_iter7_reg;
reg   [4:0] lshr_ln_reg_614_pp0_iter8_reg;
reg   [4:0] lshr_ln_reg_614_pp0_iter9_reg;
reg   [4:0] lshr_ln_reg_614_pp0_iter10_reg;
reg   [4:0] lshr_ln_reg_614_pp0_iter11_reg;
reg   [4:0] lshr_ln_reg_614_pp0_iter12_reg;
reg   [4:0] lshr_ln_reg_614_pp0_iter13_reg;
reg   [4:0] lshr_ln_reg_614_pp0_iter14_reg;
reg   [4:0] lshr_ln_reg_614_pp0_iter15_reg;
reg   [4:0] lshr_ln_reg_614_pp0_iter16_reg;
reg   [4:0] lshr_ln_reg_614_pp0_iter17_reg;
reg   [4:0] lshr_ln_reg_614_pp0_iter18_reg;
reg   [4:0] lshr_ln_reg_614_pp0_iter19_reg;
reg   [4:0] lshr_ln_reg_614_pp0_iter20_reg;
reg   [15:0] val_reg_619;
reg   [15:0] running_sums_2_load_reg_624;
reg    ap_enable_reg_pp0_iter1;
wire   [15:0] grp_fu_219_p2;
reg   [15:0] sum_reg_634;
reg   [15:0] tmp_90_i_i_reg_645;
reg   [15:0] tmp_90_i_i_reg_645_pp0_iter8_reg;
reg   [15:0] tmp_90_i_i_reg_645_pp0_iter9_reg;
reg   [15:0] tmp_90_i_i_reg_645_pp0_iter10_reg;
reg   [15:0] tmp_90_i_i_reg_645_pp0_iter11_reg;
reg   [15:0] tmp_91_i_i_reg_650;
reg   [15:0] tmp_91_i_i_reg_650_pp0_iter8_reg;
reg   [15:0] tmp_91_i_i_reg_650_pp0_iter9_reg;
reg   [15:0] tmp_91_i_i_reg_650_pp0_iter10_reg;
reg   [15:0] tmp_91_i_i_reg_650_pp0_iter11_reg;
reg   [15:0] tmp_91_i_i_reg_650_pp0_iter12_reg;
reg   [15:0] tmp_91_i_i_reg_650_pp0_iter13_reg;
reg   [15:0] tmp_91_i_i_reg_650_pp0_iter14_reg;
reg   [15:0] tmp_91_i_i_reg_650_pp0_iter15_reg;
wire   [15:0] grp_fu_227_p2;
reg   [15:0] sub_i_i_i_reg_655;
wire   [15:0] grp_fu_231_p2;
reg   [15:0] normalized_reg_665;
wire   [15:0] grp_fu_223_p2;
reg   [15:0] biased_reg_675;
reg    ap_block_state1;
wire    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_exit_iter0_state2;
reg    ap_enable_reg_pp0_iter2;
reg    ap_enable_reg_pp0_iter3;
reg    ap_enable_reg_pp0_iter4;
reg    ap_enable_reg_pp0_iter5;
reg    ap_enable_reg_pp0_iter6;
reg    ap_enable_reg_pp0_iter7;
reg    ap_enable_reg_pp0_iter8;
reg    ap_enable_reg_pp0_iter9;
reg    ap_enable_reg_pp0_iter10;
reg    ap_enable_reg_pp0_iter11;
reg    ap_enable_reg_pp0_iter12;
reg    ap_enable_reg_pp0_iter13;
reg    ap_enable_reg_pp0_iter14;
reg    ap_enable_reg_pp0_iter15;
reg    ap_enable_reg_pp0_iter16;
reg    ap_enable_reg_pp0_iter17;
reg    ap_enable_reg_pp0_iter18;
reg    ap_enable_reg_pp0_iter19;
reg    ap_enable_reg_pp0_iter20;
reg    ap_enable_reg_pp0_iter21;
reg    ap_enable_reg_pp0_iter22;
wire    ap_block_pp0_stage0;
wire   [63:0] sext_ln109_fu_509_p1;
reg   [15:0] quad_3_27_fu_114;
wire   [15:0] quad_3_38_fu_475_p3;
reg   [15:0] quad_3_26_fu_118;
wire   [15:0] quad_3_37_fu_467_p3;
reg   [15:0] quad_3_28_fu_122;
wire   [15:0] quad_3_35_fu_451_p3;
reg   [15:0] quad_3_29_fu_126;
wire   [15:0] quad_3_32_fu_427_p3;
wire   [15:0] grp_fu_223_p1;
wire   [15:0] grp_fu_227_p1;
wire   [15:0] grp_fu_231_p1;
wire   [7:0] tmp_fu_235_p3;
wire   [4:0] tmp_s_fu_247_p3;
wire   [8:0] zext_ln109_fu_243_p1;
wire   [8:0] zext_ln109_5_fu_255_p1;
wire   [8:0] sub_ln109_fu_259_p2;
wire   [9:0] sub_ln109_cast_fu_265_p1;
wire   [9:0] zext_ln109_6_fu_269_p1;
wire   [0:0] icmp_ln103_fu_301_p2;
wire   [15:0] trunc_ln95_fu_329_p1;
wire   [15:0] data_V_fu_378_p1;
wire   [0:0] p_Result_s_fu_381_p3;
wire   [0:0] icmp_ln99_fu_396_p2;
wire   [15:0] quad_0_fu_389_p3;
wire   [0:0] icmp_ln99_5_fu_409_p2;
wire   [15:0] quad_3_fu_401_p3;
wire   [0:0] icmp_ln99_6_fu_422_p2;
wire   [15:0] quad_3_31_fu_414_p3;
wire   [15:0] quad_3_33_fu_435_p3;
wire   [15:0] quad_3_34_fu_443_p3;
wire   [15:0] quad_3_36_fu_459_p3;
wire   [14:0] tmp_61_fu_503_p3;
wire   [15:0] bitcast_ln109_9_fu_526_p1;
wire   [15:0] bitcast_ln109_8_fu_522_p1;
wire   [15:0] bitcast_ln109_7_fu_518_p1;
wire   [15:0] bitcast_ln109_fu_514_p1;
wire    ap_CS_fsm_state25;
reg   [2:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
#0 ap_enable_reg_pp0_iter4 = 1'b0;
#0 ap_enable_reg_pp0_iter5 = 1'b0;
#0 ap_enable_reg_pp0_iter6 = 1'b0;
#0 ap_enable_reg_pp0_iter7 = 1'b0;
#0 ap_enable_reg_pp0_iter8 = 1'b0;
#0 ap_enable_reg_pp0_iter9 = 1'b0;
#0 ap_enable_reg_pp0_iter10 = 1'b0;
#0 ap_enable_reg_pp0_iter11 = 1'b0;
#0 ap_enable_reg_pp0_iter12 = 1'b0;
#0 ap_enable_reg_pp0_iter13 = 1'b0;
#0 ap_enable_reg_pp0_iter14 = 1'b0;
#0 ap_enable_reg_pp0_iter15 = 1'b0;
#0 ap_enable_reg_pp0_iter16 = 1'b0;
#0 ap_enable_reg_pp0_iter17 = 1'b0;
#0 ap_enable_reg_pp0_iter18 = 1'b0;
#0 ap_enable_reg_pp0_iter19 = 1'b0;
#0 ap_enable_reg_pp0_iter20 = 1'b0;
#0 ap_enable_reg_pp0_iter21 = 1'b0;
#0 ap_enable_reg_pp0_iter22 = 1'b0;
end

td_fused_top_tdf11_l2_writeOutputs_171_running_sums_2 #(
    .DataWidth( 16 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
running_sums_2_U(
    .reset(ap_rst),
    .clk(ap_clk),
    .address0(running_sums_2_addr_reg_604_pp0_iter6_reg),
    .ce0(running_sums_2_ce0),
    .we0(running_sums_2_we0),
    .d0(running_sums_2_d0),
    .address1(running_sums_2_address1),
    .ce1(running_sums_2_ce1),
    .q1(running_sums_2_q1)
);

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U719(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(running_sums_2_load_reg_624),
    .din1(val_reg_619),
    .dout(grp_fu_219_p2)
);

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U720(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(normalized_reg_665),
    .din1(grp_fu_223_p1),
    .dout(grp_fu_223_p2)
);

td_fused_top_hsub_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hsub_16ns_16ns_16_5_full_dsp_1_U721(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(sum_reg_634),
    .din1(grp_fu_227_p1),
    .dout(grp_fu_227_p2)
);

td_fused_top_hmul_16ns_16ns_16_4_max_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hmul_16ns_16ns_16_4_max_dsp_1_U722(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(sub_i_i_i_reg_655),
    .din1(grp_fu_231_p1),
    .dout(grp_fu_231_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state25)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b1 == ap_condition_pp0_exit_iter0_state2) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((~((ap_start == 1'b0) | (write4_empty_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            if ((1'b1 == ap_condition_pp0_exit_iter0_state2)) begin
                ap_enable_reg_pp0_iter1 <= (1'b1 ^ ap_condition_pp0_exit_iter0_state2);
            end else if ((1'b1 == 1'b1)) begin
                ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
            end
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter10 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter10 <= ap_enable_reg_pp0_iter9;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter11 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter11 <= ap_enable_reg_pp0_iter10;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter12 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter12 <= ap_enable_reg_pp0_iter11;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter13 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter13 <= ap_enable_reg_pp0_iter12;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter14 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter14 <= ap_enable_reg_pp0_iter13;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter15 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter15 <= ap_enable_reg_pp0_iter14;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter16 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter16 <= ap_enable_reg_pp0_iter15;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter17 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter17 <= ap_enable_reg_pp0_iter16;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter18 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter18 <= ap_enable_reg_pp0_iter17;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter19 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter19 <= ap_enable_reg_pp0_iter18;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter20 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter20 <= ap_enable_reg_pp0_iter19;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter21 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter21 <= ap_enable_reg_pp0_iter20;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter22 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter22 <= ap_enable_reg_pp0_iter21;
        end else if ((~((ap_start == 1'b0) | (write4_empty_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter22 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter4 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter5 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter5 <= ap_enable_reg_pp0_iter4;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter6 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter6 <= ap_enable_reg_pp0_iter5;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter7 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter7 <= ap_enable_reg_pp0_iter6;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter8 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter8 <= ap_enable_reg_pp0_iter7;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter9 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter9 <= ap_enable_reg_pp0_iter8;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (icmp_ln86_fu_285_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        ochan_reg_208 <= ochan_1_fu_279_p2;
    end else if ((~((ap_start == 1'b0) | (write4_empty_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ochan_reg_208 <= 8'd0;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state1)) begin
        add_ln109_reg_573 <= add_ln109_fu_273_p2;
        write4_read_reg_567 <= write4_dout;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (icmp_ln86_fu_285_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        and_ln103_reg_610 <= and_ln103_fu_307_p2;
        running_sums_2_addr_reg_604 <= zext_ln89_fu_295_p1;
        trunc_ln86_reg_587 <= trunc_ln86_fu_291_p1;
        zext_ln89_reg_594[7 : 0] <= zext_ln89_fu_295_p1[7 : 0];
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        and_ln103_reg_610_pp0_iter10_reg <= and_ln103_reg_610_pp0_iter9_reg;
        and_ln103_reg_610_pp0_iter11_reg <= and_ln103_reg_610_pp0_iter10_reg;
        and_ln103_reg_610_pp0_iter12_reg <= and_ln103_reg_610_pp0_iter11_reg;
        and_ln103_reg_610_pp0_iter13_reg <= and_ln103_reg_610_pp0_iter12_reg;
        and_ln103_reg_610_pp0_iter14_reg <= and_ln103_reg_610_pp0_iter13_reg;
        and_ln103_reg_610_pp0_iter15_reg <= and_ln103_reg_610_pp0_iter14_reg;
        and_ln103_reg_610_pp0_iter16_reg <= and_ln103_reg_610_pp0_iter15_reg;
        and_ln103_reg_610_pp0_iter17_reg <= and_ln103_reg_610_pp0_iter16_reg;
        and_ln103_reg_610_pp0_iter18_reg <= and_ln103_reg_610_pp0_iter17_reg;
        and_ln103_reg_610_pp0_iter19_reg <= and_ln103_reg_610_pp0_iter18_reg;
        and_ln103_reg_610_pp0_iter20_reg <= and_ln103_reg_610_pp0_iter19_reg;
        and_ln103_reg_610_pp0_iter2_reg <= and_ln103_reg_610_pp0_iter1_reg;
        and_ln103_reg_610_pp0_iter3_reg <= and_ln103_reg_610_pp0_iter2_reg;
        and_ln103_reg_610_pp0_iter4_reg <= and_ln103_reg_610_pp0_iter3_reg;
        and_ln103_reg_610_pp0_iter5_reg <= and_ln103_reg_610_pp0_iter4_reg;
        and_ln103_reg_610_pp0_iter6_reg <= and_ln103_reg_610_pp0_iter5_reg;
        and_ln103_reg_610_pp0_iter7_reg <= and_ln103_reg_610_pp0_iter6_reg;
        and_ln103_reg_610_pp0_iter8_reg <= and_ln103_reg_610_pp0_iter7_reg;
        and_ln103_reg_610_pp0_iter9_reg <= and_ln103_reg_610_pp0_iter8_reg;
        biased_reg_675 <= grp_fu_223_p2;
        lshr_ln_reg_614_pp0_iter10_reg <= lshr_ln_reg_614_pp0_iter9_reg;
        lshr_ln_reg_614_pp0_iter11_reg <= lshr_ln_reg_614_pp0_iter10_reg;
        lshr_ln_reg_614_pp0_iter12_reg <= lshr_ln_reg_614_pp0_iter11_reg;
        lshr_ln_reg_614_pp0_iter13_reg <= lshr_ln_reg_614_pp0_iter12_reg;
        lshr_ln_reg_614_pp0_iter14_reg <= lshr_ln_reg_614_pp0_iter13_reg;
        lshr_ln_reg_614_pp0_iter15_reg <= lshr_ln_reg_614_pp0_iter14_reg;
        lshr_ln_reg_614_pp0_iter16_reg <= lshr_ln_reg_614_pp0_iter15_reg;
        lshr_ln_reg_614_pp0_iter17_reg <= lshr_ln_reg_614_pp0_iter16_reg;
        lshr_ln_reg_614_pp0_iter18_reg <= lshr_ln_reg_614_pp0_iter17_reg;
        lshr_ln_reg_614_pp0_iter19_reg <= lshr_ln_reg_614_pp0_iter18_reg;
        lshr_ln_reg_614_pp0_iter20_reg <= lshr_ln_reg_614_pp0_iter19_reg;
        lshr_ln_reg_614_pp0_iter2_reg <= lshr_ln_reg_614_pp0_iter1_reg;
        lshr_ln_reg_614_pp0_iter3_reg <= lshr_ln_reg_614_pp0_iter2_reg;
        lshr_ln_reg_614_pp0_iter4_reg <= lshr_ln_reg_614_pp0_iter3_reg;
        lshr_ln_reg_614_pp0_iter5_reg <= lshr_ln_reg_614_pp0_iter4_reg;
        lshr_ln_reg_614_pp0_iter6_reg <= lshr_ln_reg_614_pp0_iter5_reg;
        lshr_ln_reg_614_pp0_iter7_reg <= lshr_ln_reg_614_pp0_iter6_reg;
        lshr_ln_reg_614_pp0_iter8_reg <= lshr_ln_reg_614_pp0_iter7_reg;
        lshr_ln_reg_614_pp0_iter9_reg <= lshr_ln_reg_614_pp0_iter8_reg;
        normalized_reg_665 <= grp_fu_231_p2;
        running_sums_2_addr_reg_604_pp0_iter2_reg <= running_sums_2_addr_reg_604_pp0_iter1_reg;
        running_sums_2_addr_reg_604_pp0_iter3_reg <= running_sums_2_addr_reg_604_pp0_iter2_reg;
        running_sums_2_addr_reg_604_pp0_iter4_reg <= running_sums_2_addr_reg_604_pp0_iter3_reg;
        running_sums_2_addr_reg_604_pp0_iter5_reg <= running_sums_2_addr_reg_604_pp0_iter4_reg;
        running_sums_2_addr_reg_604_pp0_iter6_reg <= running_sums_2_addr_reg_604_pp0_iter5_reg;
        sub_i_i_i_reg_655 <= grp_fu_227_p2;
        sum_reg_634 <= grp_fu_219_p2;
        tmp_90_i_i_reg_645 <= {{l2_adjustments_q0[31:16]}};
        tmp_90_i_i_reg_645_pp0_iter10_reg <= tmp_90_i_i_reg_645_pp0_iter9_reg;
        tmp_90_i_i_reg_645_pp0_iter11_reg <= tmp_90_i_i_reg_645_pp0_iter10_reg;
        tmp_90_i_i_reg_645_pp0_iter8_reg <= tmp_90_i_i_reg_645;
        tmp_90_i_i_reg_645_pp0_iter9_reg <= tmp_90_i_i_reg_645_pp0_iter8_reg;
        tmp_91_i_i_reg_650 <= {{l2_adjustments_q0[47:32]}};
        tmp_91_i_i_reg_650_pp0_iter10_reg <= tmp_91_i_i_reg_650_pp0_iter9_reg;
        tmp_91_i_i_reg_650_pp0_iter11_reg <= tmp_91_i_i_reg_650_pp0_iter10_reg;
        tmp_91_i_i_reg_650_pp0_iter12_reg <= tmp_91_i_i_reg_650_pp0_iter11_reg;
        tmp_91_i_i_reg_650_pp0_iter13_reg <= tmp_91_i_i_reg_650_pp0_iter12_reg;
        tmp_91_i_i_reg_650_pp0_iter14_reg <= tmp_91_i_i_reg_650_pp0_iter13_reg;
        tmp_91_i_i_reg_650_pp0_iter15_reg <= tmp_91_i_i_reg_650_pp0_iter14_reg;
        tmp_91_i_i_reg_650_pp0_iter8_reg <= tmp_91_i_i_reg_650;
        tmp_91_i_i_reg_650_pp0_iter9_reg <= tmp_91_i_i_reg_650_pp0_iter8_reg;
        trunc_ln86_reg_587_pp0_iter10_reg <= trunc_ln86_reg_587_pp0_iter9_reg;
        trunc_ln86_reg_587_pp0_iter11_reg <= trunc_ln86_reg_587_pp0_iter10_reg;
        trunc_ln86_reg_587_pp0_iter12_reg <= trunc_ln86_reg_587_pp0_iter11_reg;
        trunc_ln86_reg_587_pp0_iter13_reg <= trunc_ln86_reg_587_pp0_iter12_reg;
        trunc_ln86_reg_587_pp0_iter14_reg <= trunc_ln86_reg_587_pp0_iter13_reg;
        trunc_ln86_reg_587_pp0_iter15_reg <= trunc_ln86_reg_587_pp0_iter14_reg;
        trunc_ln86_reg_587_pp0_iter16_reg <= trunc_ln86_reg_587_pp0_iter15_reg;
        trunc_ln86_reg_587_pp0_iter17_reg <= trunc_ln86_reg_587_pp0_iter16_reg;
        trunc_ln86_reg_587_pp0_iter18_reg <= trunc_ln86_reg_587_pp0_iter17_reg;
        trunc_ln86_reg_587_pp0_iter19_reg <= trunc_ln86_reg_587_pp0_iter18_reg;
        trunc_ln86_reg_587_pp0_iter20_reg <= trunc_ln86_reg_587_pp0_iter19_reg;
        trunc_ln86_reg_587_pp0_iter2_reg <= trunc_ln86_reg_587_pp0_iter1_reg;
        trunc_ln86_reg_587_pp0_iter3_reg <= trunc_ln86_reg_587_pp0_iter2_reg;
        trunc_ln86_reg_587_pp0_iter4_reg <= trunc_ln86_reg_587_pp0_iter3_reg;
        trunc_ln86_reg_587_pp0_iter5_reg <= trunc_ln86_reg_587_pp0_iter4_reg;
        trunc_ln86_reg_587_pp0_iter6_reg <= trunc_ln86_reg_587_pp0_iter5_reg;
        trunc_ln86_reg_587_pp0_iter7_reg <= trunc_ln86_reg_587_pp0_iter6_reg;
        trunc_ln86_reg_587_pp0_iter8_reg <= trunc_ln86_reg_587_pp0_iter7_reg;
        trunc_ln86_reg_587_pp0_iter9_reg <= trunc_ln86_reg_587_pp0_iter8_reg;
        zext_ln89_reg_594_pp0_iter2_reg[7 : 0] <= zext_ln89_reg_594_pp0_iter1_reg[7 : 0];
        zext_ln89_reg_594_pp0_iter3_reg[7 : 0] <= zext_ln89_reg_594_pp0_iter2_reg[7 : 0];
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        and_ln103_reg_610_pp0_iter1_reg <= and_ln103_reg_610;
        lshr_ln_reg_614_pp0_iter1_reg <= lshr_ln_reg_614;
        running_sums_2_addr_reg_604_pp0_iter1_reg <= running_sums_2_addr_reg_604;
        trunc_ln86_reg_587_pp0_iter1_reg <= trunc_ln86_reg_587;
        val_reg_619 <= l2_partial_sums_q0;
        zext_ln89_reg_594_pp0_iter1_reg[7 : 0] <= zext_ln89_reg_594[7 : 0];
    end
end

always @ (posedge ap_clk) begin
    if (((1'd1 == and_ln103_fu_307_p2) & (1'b1 == ap_CS_fsm_pp0_stage0) & (icmp_ln86_fu_285_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        lshr_ln_reg_614 <= {{ochan_reg_208[6:2]}};
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        quad_3_26_fu_118 <= quad_3_37_fu_467_p3;
        quad_3_27_fu_114 <= quad_3_38_fu_475_p3;
        quad_3_28_fu_122 <= quad_3_35_fu_451_p3;
        quad_3_29_fu_126 <= quad_3_32_fu_427_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        running_sums_2_load_reg_624 <= running_sums_2_q1;
    end
end

always @ (*) begin
    if ((icmp_ln86_fu_285_p2 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state2 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state2 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state25)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter22 == 1'b0) & (ap_enable_reg_pp0_iter21 == 1'b0) & (ap_enable_reg_pp0_iter20 == 1'b0) & (ap_enable_reg_pp0_iter19 == 1'b0) & (ap_enable_reg_pp0_iter18 == 1'b0) & (ap_enable_reg_pp0_iter17 == 1'b0) & (ap_enable_reg_pp0_iter16 == 1'b0) & (ap_enable_reg_pp0_iter15 == 1'b0) & (ap_enable_reg_pp0_iter14 == 1'b0) & (ap_enable_reg_pp0_iter13 == 1'b0) & (ap_enable_reg_pp0_iter12 == 1'b0) & (ap_enable_reg_pp0_iter11 == 1'b0) & (ap_enable_reg_pp0_iter10 == 1'b0) & (ap_enable_reg_pp0_iter9 == 1'b0) & (ap_enable_reg_pp0_iter8 == 1'b0) & (ap_enable_reg_pp0_iter7 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state25)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_01_blk_n = indices_01_empty_n;
    end else begin
        indices_01_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (write4_empty_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_01_read = 1'b1;
    end else begin
        indices_01_read = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_12_blk_n = indices_12_empty_n;
    end else begin
        indices_12_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (write4_empty_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_12_read = 1'b1;
    end else begin
        indices_12_read = 1'b0;
    end
end

always @ (*) begin
    if ((((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001)) | ((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001)) | ((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001)) | ((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
        l2_adjustments_ce0 = 1'b1;
    end else begin
        l2_adjustments_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        l2_partial_sums_ce0 = 1'b1;
    end else begin
        l2_partial_sums_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001)) | ((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
        out_data_ce1 = 1'b1;
    end else begin
        out_data_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'd1 == and_ln103_reg_610_pp0_iter20_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        out_data_we1 = 1'b1;
    end else begin
        out_data_we1 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        running_sums_2_ce0 = 1'b1;
    end else begin
        running_sums_2_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        running_sums_2_ce1 = 1'b1;
    end else begin
        running_sums_2_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        running_sums_2_we0 = 1'b1;
    end else begin
        running_sums_2_we0 = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        write4_blk_n = write4_empty_n;
    end else begin
        write4_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (write4_empty_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        write4_read = 1'b1;
    end else begin
        write4_read = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_start == 1'b0) | (write4_empty_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((~((ap_enable_reg_pp0_iter0 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0) & (icmp_ln86_fu_285_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone)) & ~((ap_enable_reg_pp0_iter22 == 1'b1) & (ap_enable_reg_pp0_iter21 == 1'b0) & (1'b0 == ap_block_pp0_stage0_subdone)))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0) & (icmp_ln86_fu_285_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone)) | ((ap_enable_reg_pp0_iter22 == 1'b1) & (ap_enable_reg_pp0_iter21 == 1'b0) & (1'b0 == ap_block_pp0_stage0_subdone)))) begin
                ap_NS_fsm = ap_ST_fsm_state25;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state25 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln109_fu_273_p2 = ((sub_ln109_cast_fu_265_p1) + (zext_ln109_6_fu_269_p1));

assign and_ln103_fu_307_p2 = (write4_read_reg_567 & icmp_ln103_fu_301_p2);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state25 = ap_CS_fsm[32'd2];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (write4_empty_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1));
end

assign ap_block_state10_pp0_stage0_iter8 = ~(1'b1 == 1'b1);

assign ap_block_state11_pp0_stage0_iter9 = ~(1'b1 == 1'b1);

assign ap_block_state12_pp0_stage0_iter10 = ~(1'b1 == 1'b1);

assign ap_block_state13_pp0_stage0_iter11 = ~(1'b1 == 1'b1);

assign ap_block_state14_pp0_stage0_iter12 = ~(1'b1 == 1'b1);

assign ap_block_state15_pp0_stage0_iter13 = ~(1'b1 == 1'b1);

assign ap_block_state16_pp0_stage0_iter14 = ~(1'b1 == 1'b1);

assign ap_block_state17_pp0_stage0_iter15 = ~(1'b1 == 1'b1);

assign ap_block_state18_pp0_stage0_iter16 = ~(1'b1 == 1'b1);

assign ap_block_state19_pp0_stage0_iter17 = ~(1'b1 == 1'b1);

assign ap_block_state20_pp0_stage0_iter18 = ~(1'b1 == 1'b1);

assign ap_block_state21_pp0_stage0_iter19 = ~(1'b1 == 1'b1);

assign ap_block_state22_pp0_stage0_iter20 = ~(1'b1 == 1'b1);

assign ap_block_state23_pp0_stage0_iter21 = ~(1'b1 == 1'b1);

assign ap_block_state24_pp0_stage0_iter22 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter4 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage0_iter5 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage0_iter6 = ~(1'b1 == 1'b1);

assign ap_block_state9_pp0_stage0_iter7 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign bitcast_ln109_7_fu_518_p1 = quad_3_37_fu_467_p3;

assign bitcast_ln109_8_fu_522_p1 = quad_3_35_fu_451_p3;

assign bitcast_ln109_9_fu_526_p1 = quad_3_32_fu_427_p3;

assign bitcast_ln109_fu_514_p1 = quad_3_38_fu_475_p3;

assign data_V_fu_378_p1 = biased_reg_675;

assign grp_fu_223_p1 = tmp_91_i_i_reg_650_pp0_iter15_reg;

assign grp_fu_227_p1 = trunc_ln95_fu_329_p1;

assign grp_fu_231_p1 = tmp_90_i_i_reg_645_pp0_iter11_reg;

assign icmp_ln103_fu_301_p2 = ((trunc_ln86_fu_291_p1 == 2'd3) ? 1'b1 : 1'b0);

assign icmp_ln86_fu_285_p2 = ((ochan_reg_208 == 8'd128) ? 1'b1 : 1'b0);

assign icmp_ln99_5_fu_409_p2 = ((trunc_ln86_reg_587_pp0_iter20_reg == 2'd1) ? 1'b1 : 1'b0);

assign icmp_ln99_6_fu_422_p2 = ((trunc_ln86_reg_587_pp0_iter20_reg == 2'd0) ? 1'b1 : 1'b0);

assign icmp_ln99_fu_396_p2 = ((trunc_ln86_reg_587_pp0_iter20_reg == 2'd2) ? 1'b1 : 1'b0);

assign l2_adjustments_address0 = zext_ln89_reg_594_pp0_iter3_reg;

assign l2_partial_sums_address0 = zext_ln89_fu_295_p1;

assign ochan_1_fu_279_p2 = (ochan_reg_208 + 8'd1);

assign out_data_address1 = sext_ln109_fu_509_p1;

assign out_data_d1 = {{{{bitcast_ln109_9_fu_526_p1}, {bitcast_ln109_8_fu_522_p1}}, {bitcast_ln109_7_fu_518_p1}}, {bitcast_ln109_fu_514_p1}};

assign p_Result_s_fu_381_p3 = data_V_fu_378_p1[32'd15];

assign quad_0_fu_389_p3 = ((p_Result_s_fu_381_p3[0:0] == 1'b1) ? 16'd0 : biased_reg_675);

assign quad_3_31_fu_414_p3 = ((icmp_ln99_5_fu_409_p2[0:0] == 1'b1) ? quad_3_29_fu_126 : quad_3_fu_401_p3);

assign quad_3_32_fu_427_p3 = ((icmp_ln99_6_fu_422_p2[0:0] == 1'b1) ? quad_3_29_fu_126 : quad_3_31_fu_414_p3);

assign quad_3_33_fu_435_p3 = ((icmp_ln99_fu_396_p2[0:0] == 1'b1) ? quad_0_fu_389_p3 : quad_3_28_fu_122);

assign quad_3_34_fu_443_p3 = ((icmp_ln99_5_fu_409_p2[0:0] == 1'b1) ? quad_3_28_fu_122 : quad_3_33_fu_435_p3);

assign quad_3_35_fu_451_p3 = ((icmp_ln99_6_fu_422_p2[0:0] == 1'b1) ? quad_3_28_fu_122 : quad_3_34_fu_443_p3);

assign quad_3_36_fu_459_p3 = ((icmp_ln99_5_fu_409_p2[0:0] == 1'b1) ? quad_0_fu_389_p3 : quad_3_26_fu_118);

assign quad_3_37_fu_467_p3 = ((icmp_ln99_6_fu_422_p2[0:0] == 1'b1) ? quad_3_26_fu_118 : quad_3_36_fu_459_p3);

assign quad_3_38_fu_475_p3 = ((icmp_ln99_6_fu_422_p2[0:0] == 1'b1) ? quad_0_fu_389_p3 : quad_3_27_fu_114);

assign quad_3_fu_401_p3 = ((icmp_ln99_fu_396_p2[0:0] == 1'b1) ? quad_3_29_fu_126 : quad_0_fu_389_p3);

assign running_sums_2_address1 = zext_ln89_fu_295_p1;

assign running_sums_2_d0 = ((write4_read_reg_567[0:0] == 1'b1) ? 16'd0 : sum_reg_634);

assign sext_ln109_fu_509_p1 = (tmp_61_fu_503_p3);

assign sub_ln109_cast_fu_265_p1 = (sub_ln109_fu_259_p2);

assign sub_ln109_fu_259_p2 = (zext_ln109_fu_243_p1 - zext_ln109_5_fu_255_p1);

assign tmp_61_fu_503_p3 = {{add_ln109_reg_573}, {lshr_ln_reg_614_pp0_iter20_reg}};

assign tmp_fu_235_p3 = {{indices_01_dout}, {4'd0}};

assign tmp_s_fu_247_p3 = {{indices_01_dout}, {1'd0}};

assign trunc_ln86_fu_291_p1 = ochan_reg_208[1:0];

assign trunc_ln95_fu_329_p1 = l2_adjustments_q0[15:0];

assign zext_ln109_5_fu_255_p1 = tmp_s_fu_247_p3;

assign zext_ln109_6_fu_269_p1 = indices_12_dout;

assign zext_ln109_fu_243_p1 = tmp_fu_235_p3;

assign zext_ln89_fu_295_p1 = ochan_reg_208;

always @ (posedge ap_clk) begin
    zext_ln89_reg_594[63:8] <= 56'b00000000000000000000000000000000000000000000000000000000;
    zext_ln89_reg_594_pp0_iter1_reg[63:8] <= 56'b00000000000000000000000000000000000000000000000000000000;
    zext_ln89_reg_594_pp0_iter2_reg[63:8] <= 56'b00000000000000000000000000000000000000000000000000000000;
    zext_ln89_reg_594_pp0_iter3_reg[63:8] <= 56'b00000000000000000000000000000000000000000000000000000000;
end

endmodule //td_fused_top_tdf11_l2_writeOutputs_171
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf11_readFilters74 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        filter_data_address0,
        filter_data_ce0,
        filter_data_q0,
        indices_23_dout,
        indices_23_empty_n,
        indices_23_read,
        weight_vecs_0_address0,
        weight_vecs_0_ce0,
        weight_vecs_0_we0,
        weight_vecs_0_d0,
        weight_vecs_0_address1,
        weight_vecs_0_ce1,
        weight_vecs_0_we1,
        weight_vecs_0_d1
);

parameter    ap_ST_fsm_state1 = 4'd1;
parameter    ap_ST_fsm_pp0_stage0 = 4'd2;
parameter    ap_ST_fsm_pp0_stage1 = 4'd4;
parameter    ap_ST_fsm_state7 = 4'd8;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [16:0] filter_data_address0;
output   filter_data_ce0;
input  [63:0] filter_data_q0;
input  [8:0] indices_23_dout;
input   indices_23_empty_n;
output   indices_23_read;
output  [9:0] weight_vecs_0_address0;
output   weight_vecs_0_ce0;
output   weight_vecs_0_we0;
output  [15:0] weight_vecs_0_d0;
output  [9:0] weight_vecs_0_address1;
output   weight_vecs_0_ce1;
output   weight_vecs_0_we1;
output  [15:0] weight_vecs_0_d1;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg filter_data_ce0;
reg indices_23_read;
reg[9:0] weight_vecs_0_address0;
reg weight_vecs_0_ce0;
reg weight_vecs_0_we0;
reg[15:0] weight_vecs_0_d0;
reg[9:0] weight_vecs_0_address1;
reg weight_vecs_0_ce1;
reg weight_vecs_0_we1;
reg[15:0] weight_vecs_0_d1;

reg    ap_done_reg;
  reg   [3:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    indices_23_blk_n;
reg   [7:0] indvar_flatten13_reg_174;
reg   [1:0] ii_reg_185;
reg   [6:0] indvar_flatten_reg_196;
reg   [1:0] jj_reg_207;
reg   [6:0] kk_0_i_i_reg_218;
wire   [12:0] sext_ln47_fu_251_p1;
reg   [12:0] sext_ln47_reg_583;
wire   [7:0] add_ln47_7_fu_255_p2;
reg   [7:0] add_ln47_7_reg_588;
wire    ap_CS_fsm_pp0_stage0;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state4_pp0_stage0_iter1;
wire    ap_block_state6_pp0_stage0_iter2;
wire    ap_block_pp0_stage0_11001;
wire   [0:0] icmp_ln47_fu_261_p2;
reg   [0:0] icmp_ln47_reg_593;
reg   [0:0] icmp_ln47_reg_593_pp0_iter1_reg;
wire   [0:0] icmp_ln48_fu_273_p2;
reg   [0:0] icmp_ln48_reg_597;
wire   [1:0] select_ln47_7_fu_287_p3;
reg   [1:0] select_ln47_7_reg_602;
wire   [6:0] select_ln48_fu_356_p3;
reg   [6:0] select_ln48_reg_609;
wire   [1:0] select_ln48_13_fu_364_p3;
reg   [1:0] select_ln48_13_reg_615;
wire   [5:0] empty_138_fu_382_p1;
reg   [5:0] empty_138_reg_621;
reg   [5:0] empty_138_reg_621_pp0_iter1_reg;
wire   [6:0] add_ln48_7_fu_405_p2;
reg   [6:0] add_ln48_7_reg_633;
wire   [6:0] add_ln49_fu_411_p2;
reg   [6:0] add_ln49_reg_638;
wire    ap_CS_fsm_pp0_stage1;
wire    ap_block_state3_pp0_stage1_iter0;
wire    ap_block_state5_pp0_stage1_iter1;
wire    ap_block_pp0_stage1_11001;
wire   [6:0] select_ln48_14_fu_416_p3;
reg   [6:0] select_ln48_14_reg_643;
wire   [5:0] add_ln55_26_fu_449_p2;
reg   [5:0] add_ln55_26_reg_648;
wire   [9:0] add_ln55_27_fu_470_p2;
reg   [9:0] add_ln55_27_reg_655;
reg   [15:0] tmp_88_i_i_reg_660;
reg   [15:0] tmp_89_i_i_reg_665;
reg    ap_block_state1;
wire    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_exit_iter0_state2;
reg    ap_enable_reg_pp0_iter1;
wire    ap_block_pp0_stage1_subdone;
reg    ap_enable_reg_pp0_iter2;
reg   [7:0] ap_phi_mux_indvar_flatten13_phi_fu_178_p4;
wire    ap_block_pp0_stage0;
reg   [1:0] ap_phi_mux_ii_phi_fu_189_p4;
reg   [6:0] ap_phi_mux_indvar_flatten_phi_fu_200_p4;
reg   [1:0] ap_phi_mux_jj_phi_fu_211_p4;
reg   [6:0] ap_phi_mux_kk_0_i_i_phi_fu_222_p4;
wire   [63:0] tmp_17_fu_396_p3;
wire   [63:0] zext_ln55_67_fu_476_p1;
wire    ap_block_pp0_stage1;
wire   [63:0] sext_ln55_3_fu_501_p1;
wire   [63:0] sext_ln55_4_fu_553_p1;
wire   [63:0] sext_ln55_5_fu_574_p1;
wire   [15:0] bitcast_ln55_fu_484_p1;
wire   [15:0] bitcast_ln55_1_fu_516_p1;
wire   [15:0] bitcast_ln55_2_fu_558_p1;
wire   [15:0] bitcast_ln55_3_fu_579_p1;
wire   [10:0] tmp_fu_233_p3;
wire   [11:0] zext_ln55_60_fu_241_p1;
wire   [11:0] zext_ln55_fu_229_p1;
wire   [11:0] sub_ln55_fu_245_p2;
wire   [1:0] add_ln47_fu_267_p2;
wire   [12:0] zext_ln55_62_fu_295_p1;
wire   [12:0] add_ln55_fu_299_p2;
wire   [14:0] tmp_56_fu_308_p3;
wire   [59:0] sext_ln55_2_fu_316_p1;
wire   [59:0] sext_ln55_fu_304_p1;
wire   [0:0] icmp_ln49_fu_332_p2;
wire   [0:0] xor_ln47_fu_326_p2;
wire   [1:0] select_ln47_fu_279_p3;
wire   [0:0] and_ln47_fu_338_p2;
wire   [0:0] or_ln48_fu_350_p2;
wire   [1:0] add_ln48_fu_344_p2;
wire   [59:0] sub_ln55_15_fu_320_p2;
wire   [59:0] zext_ln55_65_fu_372_p1;
wire   [59:0] add_ln55_25_fu_376_p2;
wire   [3:0] lshr_ln_fu_386_p4;
wire   [3:0] tmp_s_fu_425_p3;
wire   [4:0] zext_ln55_63_fu_432_p1;
wire   [4:0] zext_ln55_61_fu_422_p1;
wire   [4:0] sub_ln55_16_fu_436_p2;
wire   [5:0] sext_ln48_fu_442_p1;
wire   [5:0] zext_ln55_64_fu_446_p1;
wire   [3:0] trunc_ln55_fu_455_p1;
wire   [9:0] tmp_166_cast_fu_459_p3;
wire   [9:0] zext_ln55_66_fu_467_p1;
wire   [15:0] trunc_ln55_4_fu_480_p1;
wire   [5:0] or_ln49_fu_489_p2;
wire   [11:0] tmp_57_fu_494_p3;
wire   [15:0] tmp_87_i_i_fu_506_p4;
wire   [5:0] or_ln49_1_fu_541_p2;
wire   [11:0] tmp_58_fu_546_p3;
wire   [5:0] or_ln49_2_fu_562_p2;
wire   [11:0] tmp_59_fu_567_p3;
wire    ap_CS_fsm_state7;
reg   [3:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 4'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state7)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b1 == ap_condition_pp0_exit_iter0_state2))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1)) | ((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b0)))) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end else if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter2 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_reg_593 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ii_reg_185 <= select_ln47_7_reg_602;
    end else if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ii_reg_185 <= 2'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_reg_593 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        indvar_flatten13_reg_174 <= add_ln47_7_reg_588;
    end else if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indvar_flatten13_reg_174 <= 8'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_reg_593 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        indvar_flatten_reg_196 <= select_ln48_14_reg_643;
    end else if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indvar_flatten_reg_196 <= 7'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_reg_593 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        jj_reg_207 <= select_ln48_13_reg_615;
    end else if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        jj_reg_207 <= 2'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_reg_593 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        kk_0_i_i_reg_218 <= add_ln49_reg_638;
    end else if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        kk_0_i_i_reg_218 <= 7'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        add_ln47_7_reg_588 <= add_ln47_7_fu_255_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_fu_261_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        add_ln48_7_reg_633 <= add_ln48_7_fu_405_p2;
        empty_138_reg_621 <= empty_138_fu_382_p1;
        icmp_ln48_reg_597 <= icmp_ln48_fu_273_p2;
        select_ln48_reg_609 <= select_ln48_fu_356_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_reg_593 == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
        add_ln49_reg_638 <= add_ln49_fu_411_p2;
        select_ln48_14_reg_643 <= select_ln48_14_fu_416_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_reg_593 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        add_ln55_26_reg_648 <= add_ln55_26_fu_449_p2;
        add_ln55_27_reg_655 <= add_ln55_27_fu_470_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        empty_138_reg_621_pp0_iter1_reg <= empty_138_reg_621;
        icmp_ln47_reg_593 <= icmp_ln47_fu_261_p2;
        icmp_ln47_reg_593_pp0_iter1_reg <= icmp_ln47_reg_593;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_fu_261_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        select_ln47_7_reg_602 <= select_ln47_7_fu_287_p3;
        select_ln48_13_reg_615 <= select_ln48_13_fu_364_p3;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state1)) begin
        sext_ln47_reg_583 <= sext_ln47_fu_251_p1;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_reg_593_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
        tmp_88_i_i_reg_660 <= {{filter_data_q0[47:32]}};
        tmp_89_i_i_reg_665 <= {{filter_data_q0[63:48]}};
    end
end

always @ (*) begin
    if ((icmp_ln47_fu_261_p2 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state2 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state2 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state7)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln47_reg_593 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_ii_phi_fu_189_p4 = select_ln47_7_reg_602;
    end else begin
        ap_phi_mux_ii_phi_fu_189_p4 = ii_reg_185;
    end
end

always @ (*) begin
    if (((icmp_ln47_reg_593 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_indvar_flatten13_phi_fu_178_p4 = add_ln47_7_reg_588;
    end else begin
        ap_phi_mux_indvar_flatten13_phi_fu_178_p4 = indvar_flatten13_reg_174;
    end
end

always @ (*) begin
    if (((icmp_ln47_reg_593 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_indvar_flatten_phi_fu_200_p4 = select_ln48_14_reg_643;
    end else begin
        ap_phi_mux_indvar_flatten_phi_fu_200_p4 = indvar_flatten_reg_196;
    end
end

always @ (*) begin
    if (((icmp_ln47_reg_593 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_jj_phi_fu_211_p4 = select_ln48_13_reg_615;
    end else begin
        ap_phi_mux_jj_phi_fu_211_p4 = jj_reg_207;
    end
end

always @ (*) begin
    if (((icmp_ln47_reg_593 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_kk_0_i_i_phi_fu_222_p4 = add_ln49_reg_638;
    end else begin
        ap_phi_mux_kk_0_i_i_phi_fu_222_p4 = kk_0_i_i_reg_218;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state7)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1)) | ((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)) | ((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1)))) begin
        filter_data_ce0 = 1'b1;
    end else begin
        filter_data_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_23_blk_n = indices_23_empty_n;
    end else begin
        indices_23_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_23_read = 1'b1;
    end else begin
        indices_23_read = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        weight_vecs_0_address0 = sext_ln55_5_fu_574_p1;
    end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        weight_vecs_0_address0 = sext_ln55_3_fu_501_p1;
    end else begin
        weight_vecs_0_address0 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        weight_vecs_0_address1 = sext_ln55_4_fu_553_p1;
    end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        weight_vecs_0_address1 = zext_ln55_67_fu_476_p1;
    end else begin
        weight_vecs_0_address1 = 'bx;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1)) | ((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1)))) begin
        weight_vecs_0_ce0 = 1'b1;
    end else begin
        weight_vecs_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1)) | ((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1)))) begin
        weight_vecs_0_ce1 = 1'b1;
    end else begin
        weight_vecs_0_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        weight_vecs_0_d0 = bitcast_ln55_3_fu_579_p1;
    end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        weight_vecs_0_d0 = bitcast_ln55_1_fu_516_p1;
    end else begin
        weight_vecs_0_d0 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        weight_vecs_0_d1 = bitcast_ln55_2_fu_558_p1;
    end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        weight_vecs_0_d1 = bitcast_ln55_fu_484_p1;
    end else begin
        weight_vecs_0_d1 = 'bx;
    end
end

always @ (*) begin
    if ((((icmp_ln47_reg_593_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1)) | ((icmp_ln47_reg_593_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1)))) begin
        weight_vecs_0_we0 = 1'b1;
    end else begin
        weight_vecs_0_we0 = 1'b0;
    end
end

always @ (*) begin
    if ((((icmp_ln47_reg_593_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1)) | ((icmp_ln47_reg_593_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1)))) begin
        weight_vecs_0_we1 = 1'b1;
    end else begin
        weight_vecs_0_we1 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((~((icmp_ln47_fu_261_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0)) & ~((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0)) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end else if ((((icmp_ln47_fu_261_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0)) | ((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_state7;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_pp0_stage1 : begin
            if ((1'b0 == ap_block_pp0_stage1_subdone)) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end
        end
        ap_ST_fsm_state7 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln47_7_fu_255_p2 = (ap_phi_mux_indvar_flatten13_phi_fu_178_p4 + 8'd1);

assign add_ln47_fu_267_p2 = (ap_phi_mux_ii_phi_fu_189_p4 + 2'd1);

assign add_ln48_7_fu_405_p2 = (ap_phi_mux_indvar_flatten_phi_fu_200_p4 + 7'd1);

assign add_ln48_fu_344_p2 = (select_ln47_fu_279_p3 + 2'd1);

assign add_ln49_fu_411_p2 = (select_ln48_reg_609 + 7'd4);

assign add_ln55_25_fu_376_p2 = (sub_ln55_15_fu_320_p2 + zext_ln55_65_fu_372_p1);

assign add_ln55_26_fu_449_p2 = ((sext_ln48_fu_442_p1) + (zext_ln55_64_fu_446_p1));

assign add_ln55_27_fu_470_p2 = (tmp_166_cast_fu_459_p3 + zext_ln55_66_fu_467_p1);

assign add_ln55_fu_299_p2 = ((sext_ln47_reg_583) + (zext_ln55_62_fu_295_p1));

assign and_ln47_fu_338_p2 = (xor_ln47_fu_326_p2 & icmp_ln49_fu_332_p2);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_pp0_stage1 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state7 = ap_CS_fsm[32'd3];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1));
end

assign ap_block_state2_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage1_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage1_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign bitcast_ln55_1_fu_516_p1 = tmp_87_i_i_fu_506_p4;

assign bitcast_ln55_2_fu_558_p1 = tmp_88_i_i_reg_660;

assign bitcast_ln55_3_fu_579_p1 = tmp_89_i_i_reg_665;

assign bitcast_ln55_fu_484_p1 = trunc_ln55_4_fu_480_p1;

assign empty_138_fu_382_p1 = select_ln48_fu_356_p3[5:0];

assign filter_data_address0 = tmp_17_fu_396_p3;

assign icmp_ln47_fu_261_p2 = ((ap_phi_mux_indvar_flatten13_phi_fu_178_p4 == 8'd144) ? 1'b1 : 1'b0);

assign icmp_ln48_fu_273_p2 = ((ap_phi_mux_indvar_flatten_phi_fu_200_p4 == 7'd48) ? 1'b1 : 1'b0);

assign icmp_ln49_fu_332_p2 = ((ap_phi_mux_kk_0_i_i_phi_fu_222_p4 == 7'd64) ? 1'b1 : 1'b0);

assign lshr_ln_fu_386_p4 = {{select_ln48_fu_356_p3[5:2]}};

assign or_ln48_fu_350_p2 = (icmp_ln48_fu_273_p2 | and_ln47_fu_338_p2);

assign or_ln49_1_fu_541_p2 = (empty_138_reg_621_pp0_iter1_reg | 6'd2);

assign or_ln49_2_fu_562_p2 = (empty_138_reg_621_pp0_iter1_reg | 6'd3);

assign or_ln49_fu_489_p2 = (empty_138_reg_621_pp0_iter1_reg | 6'd1);

assign select_ln47_7_fu_287_p3 = ((icmp_ln48_fu_273_p2[0:0] == 1'b1) ? add_ln47_fu_267_p2 : ap_phi_mux_ii_phi_fu_189_p4);

assign select_ln47_fu_279_p3 = ((icmp_ln48_fu_273_p2[0:0] == 1'b1) ? 2'd0 : ap_phi_mux_jj_phi_fu_211_p4);

assign select_ln48_13_fu_364_p3 = ((and_ln47_fu_338_p2[0:0] == 1'b1) ? add_ln48_fu_344_p2 : select_ln47_fu_279_p3);

assign select_ln48_14_fu_416_p3 = ((icmp_ln48_reg_597[0:0] == 1'b1) ? 7'd1 : add_ln48_7_reg_633);

assign select_ln48_fu_356_p3 = ((or_ln48_fu_350_p2[0:0] == 1'b1) ? 7'd0 : ap_phi_mux_kk_0_i_i_phi_fu_222_p4);

assign sext_ln47_fu_251_p1 = (sub_ln55_fu_245_p2);

assign sext_ln48_fu_442_p1 = (sub_ln55_16_fu_436_p2);

assign sext_ln55_2_fu_316_p1 = (tmp_56_fu_308_p3);

assign sext_ln55_3_fu_501_p1 = (tmp_57_fu_494_p3);

assign sext_ln55_4_fu_553_p1 = (tmp_58_fu_546_p3);

assign sext_ln55_5_fu_574_p1 = (tmp_59_fu_567_p3);

assign sext_ln55_fu_304_p1 = add_ln55_fu_299_p2;

assign sub_ln55_15_fu_320_p2 = ((sext_ln55_2_fu_316_p1) - (sext_ln55_fu_304_p1));

assign sub_ln55_16_fu_436_p2 = (zext_ln55_63_fu_432_p1 - zext_ln55_61_fu_422_p1);

assign sub_ln55_fu_245_p2 = (zext_ln55_60_fu_241_p1 - zext_ln55_fu_229_p1);

assign tmp_166_cast_fu_459_p3 = {{trunc_ln55_fu_455_p1}, {6'd0}};

assign tmp_17_fu_396_p3 = {{add_ln55_25_fu_376_p2}, {lshr_ln_fu_386_p4}};

assign tmp_56_fu_308_p3 = {{add_ln55_fu_299_p2}, {2'd0}};

assign tmp_57_fu_494_p3 = {{add_ln55_26_reg_648}, {or_ln49_fu_489_p2}};

assign tmp_58_fu_546_p3 = {{add_ln55_26_reg_648}, {or_ln49_1_fu_541_p2}};

assign tmp_59_fu_567_p3 = {{add_ln55_26_reg_648}, {or_ln49_2_fu_562_p2}};

assign tmp_87_i_i_fu_506_p4 = {{filter_data_q0[31:16]}};

assign tmp_fu_233_p3 = {{indices_23_dout}, {2'd0}};

assign tmp_s_fu_425_p3 = {{select_ln47_7_reg_602}, {2'd0}};

assign trunc_ln55_4_fu_480_p1 = filter_data_q0[15:0];

assign trunc_ln55_fu_455_p1 = add_ln55_26_fu_449_p2[3:0];

assign xor_ln47_fu_326_p2 = (icmp_ln48_fu_273_p2 ^ 1'd1);

assign zext_ln55_60_fu_241_p1 = tmp_fu_233_p3;

assign zext_ln55_61_fu_422_p1 = select_ln47_7_reg_602;

assign zext_ln55_62_fu_295_p1 = select_ln47_7_fu_287_p3;

assign zext_ln55_63_fu_432_p1 = tmp_s_fu_425_p3;

assign zext_ln55_64_fu_446_p1 = select_ln48_13_reg_615;

assign zext_ln55_65_fu_372_p1 = select_ln48_13_fu_364_p3;

assign zext_ln55_66_fu_467_p1 = select_ln48_reg_609;

assign zext_ln55_67_fu_476_p1 = add_ln55_27_reg_655;

assign zext_ln55_fu_229_p1 = indices_23_dout;

endmodule //td_fused_top_tdf11_readFilters74
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf11_readInputs75 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        in_data_address0,
        in_data_ce0,
        in_data_q0,
        indices_01_dout,
        indices_01_empty_n,
        indices_01_read,
        indices_12_dout,
        indices_12_empty_n,
        indices_12_read,
        ifmap_vec_address0,
        ifmap_vec_ce0,
        ifmap_vec_we0,
        ifmap_vec_d0,
        ifmap_vec_address1,
        ifmap_vec_ce1,
        ifmap_vec_we1,
        ifmap_vec_d1,
        indices_01_out_din,
        indices_01_out_full_n,
        indices_01_out_write,
        indices_12_out_din,
        indices_12_out_full_n,
        indices_12_out_write
);

parameter    ap_ST_fsm_state1 = 5'd1;
parameter    ap_ST_fsm_state2 = 5'd2;
parameter    ap_ST_fsm_pp0_stage0 = 5'd4;
parameter    ap_ST_fsm_pp0_stage1 = 5'd8;
parameter    ap_ST_fsm_state9 = 5'd16;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [11:0] in_data_address0;
output   in_data_ce0;
input  [63:0] in_data_q0;
input  [15:0] indices_01_dout;
input   indices_01_empty_n;
output   indices_01_read;
input  [15:0] indices_12_dout;
input   indices_12_empty_n;
output   indices_12_read;
output  [9:0] ifmap_vec_address0;
output   ifmap_vec_ce0;
output   ifmap_vec_we0;
output  [15:0] ifmap_vec_d0;
output  [9:0] ifmap_vec_address1;
output   ifmap_vec_ce1;
output   ifmap_vec_we1;
output  [15:0] ifmap_vec_d1;
output  [3:0] indices_01_out_din;
input   indices_01_out_full_n;
output   indices_01_out_write;
output  [7:0] indices_12_out_din;
input   indices_12_out_full_n;
output   indices_12_out_write;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg in_data_ce0;
reg indices_01_read;
reg indices_12_read;
reg[9:0] ifmap_vec_address0;
reg ifmap_vec_ce0;
reg ifmap_vec_we0;
reg[15:0] ifmap_vec_d0;
reg[9:0] ifmap_vec_address1;
reg ifmap_vec_ce1;
reg ifmap_vec_we1;
reg[15:0] ifmap_vec_d1;
reg indices_01_out_write;
reg indices_12_out_write;

reg    ap_done_reg;
  reg   [4:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    indices_01_blk_n;
reg    indices_12_blk_n;
reg    indices_01_out_blk_n;
reg    indices_12_out_blk_n;
reg   [7:0] indvar_flatten47_reg_224;
reg   [1:0] ii_reg_236;
reg   [6:0] indvar_flatten_reg_248;
reg   [1:0] jj_reg_259;
reg   [6:0] kk_0_i_i_reg_271;
reg   [15:0] indices_01_read_reg_960;
wire   [3:0] trunc_ln250_fu_282_p1;
reg   [3:0] trunc_ln250_reg_965;
reg   [15:0] indices_12_read_reg_970;
wire   [7:0] empty_fu_287_p1;
reg   [7:0] empty_reg_975;
wire   [17:0] p_cast_i_i_fu_304_p1;
reg   [17:0] p_cast_i_i_reg_982;
wire    ap_CS_fsm_state2;
wire   [17:0] sext_ln22_fu_314_p1;
reg   [17:0] sext_ln22_reg_988;
wire   [3:0] p_cast_fu_318_p2;
reg   [3:0] p_cast_reg_994;
wire   [0:0] or_ln23_31_fu_337_p2;
reg   [0:0] or_ln23_31_reg_1000;
wire   [7:0] p_mid137_fu_343_p2;
reg   [7:0] p_mid137_reg_1005;
wire   [3:0] p_cast5_i_i_fu_361_p2;
reg   [3:0] p_cast5_i_i_reg_1010;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_block_state3_pp0_stage0_iter0;
wire    ap_block_state5_pp0_stage0_iter1;
wire    ap_block_state7_pp0_stage0_iter2;
wire    ap_block_pp0_stage0_11001;
wire   [0:0] is_padding_fu_401_p2;
reg   [0:0] is_padding_reg_1016;
wire   [0:0] icmp_ln19_fu_407_p2;
reg   [0:0] icmp_ln19_reg_1023;
reg   [0:0] icmp_ln19_reg_1023_pp0_iter1_reg;
reg   [0:0] icmp_ln19_reg_1023_pp0_iter2_reg;
wire   [1:0] add_ln19_fu_413_p2;
reg   [1:0] add_ln19_reg_1027;
wire   [0:0] icmp_ln20_fu_419_p2;
reg   [0:0] icmp_ln20_reg_1033;
wire   [1:0] select_ln19_fu_425_p3;
reg   [1:0] select_ln19_reg_1045;
wire   [0:0] or_ln23_33_fu_456_p2;
reg   [0:0] or_ln23_33_reg_1050;
wire   [1:0] add_ln20_fu_461_p2;
reg   [1:0] add_ln20_reg_1057;
wire   [0:0] or_ln23_35_fu_496_p2;
reg   [0:0] or_ln23_35_reg_1063;
wire   [6:0] add_ln20_7_fu_502_p2;
reg   [6:0] add_ln20_7_reg_1070;
wire   [7:0] add_ln19_7_fu_508_p2;
reg   [7:0] add_ln19_7_reg_1075;
wire    ap_CS_fsm_pp0_stage1;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_state4_pp0_stage1_iter0;
wire    ap_block_state6_pp0_stage1_iter1;
wire    ap_block_state8_pp0_stage1_iter2;
wire    ap_block_pp0_stage1_11001;
wire   [1:0] select_ln19_36_fu_546_p3;
reg   [1:0] select_ln19_36_reg_1080;
wire   [6:0] select_ln20_fu_620_p3;
reg   [6:0] select_ln20_reg_1087;
wire   [1:0] select_ln20_30_fu_628_p3;
reg   [1:0] select_ln20_30_reg_1093;
wire   [0:0] select_ln20_31_fu_637_p3;
reg   [0:0] select_ln20_31_reg_1099;
reg   [0:0] select_ln20_31_reg_1099_pp0_iter1_reg;
wire   [5:0] empty_137_fu_733_p1;
reg   [5:0] empty_137_reg_1107;
reg   [5:0] empty_137_reg_1107_pp0_iter1_reg;
wire   [6:0] select_ln20_34_fu_760_p3;
reg   [6:0] select_ln20_34_reg_1119;
wire   [6:0] add_ln25_fu_766_p2;
reg   [6:0] add_ln25_reg_1124;
reg    ap_enable_reg_pp0_iter1;
wire   [5:0] add_ln33_fu_798_p2;
reg   [5:0] add_ln33_reg_1129;
wire   [9:0] add_ln33_7_fu_819_p2;
reg   [9:0] add_ln33_7_reg_1136;
wire   [15:0] select_ln33_29_fu_898_p3;
reg   [15:0] select_ln33_29_reg_1141;
wire   [15:0] select_ln33_30_fu_919_p3;
reg   [15:0] select_ln33_30_reg_1146;
wire    ap_block_pp0_stage1_subdone;
reg    ap_condition_pp0_exit_iter0_state4;
reg    ap_enable_reg_pp0_iter2;
reg   [7:0] ap_phi_mux_indvar_flatten47_phi_fu_228_p4;
wire    ap_block_pp0_stage0;
reg   [1:0] ap_phi_mux_ii_phi_fu_240_p4;
reg   [6:0] ap_phi_mux_indvar_flatten_phi_fu_252_p4;
reg   [1:0] ap_phi_mux_jj_phi_fu_263_p4;
reg   [6:0] ap_phi_mux_kk_0_i_i_phi_fu_275_p4;
wire    ap_block_pp0_stage1;
wire   [63:0] sext_ln32_fu_755_p1;
wire   [63:0] zext_ln33_29_fu_825_p1;
wire   [63:0] sext_ln33_fu_857_p1;
wire   [63:0] sext_ln33_11_fu_938_p1;
wire   [63:0] sext_ln33_12_fu_955_p1;
reg    ap_block_state1;
wire   [15:0] select_ln33_fu_837_p3;
wire   [15:0] select_ln33_28_fu_876_p3;
wire   [16:0] zext_ln19_fu_295_p1;
wire   [16:0] empty_132_fu_298_p2;
wire   [16:0] j_cast_i_i_fu_292_p1;
wire   [16:0] add_ln22_fu_308_p2;
wire   [0:0] tmp_49_fu_323_p3;
wire   [0:0] icmp_ln24_fu_331_p2;
wire   [17:0] ii_cast_i_i_fu_348_p1;
wire   [3:0] ii_cast_fu_352_p1;
wire   [17:0] empty_133_fu_356_p2;
wire   [17:0] zext_ln20_fu_372_p1;
wire   [17:0] add_ln22_7_fu_376_p2;
wire   [0:0] tmp_50_fu_381_p3;
wire   [0:0] icmp_ln24_7_fu_389_p2;
wire   [0:0] or_ln23_fu_395_p2;
wire   [0:0] empty_134_fu_366_p2;
wire   [17:0] ii_cast_i_i_mid1_fu_433_p1;
wire   [17:0] p_mid111_fu_437_p2;
wire   [0:0] p_mid113_fu_442_p2;
wire   [17:0] zext_ln20_7_fu_467_p1;
wire   [17:0] add_ln22_8_fu_471_p2;
wire   [0:0] tmp_51_fu_476_p3;
wire   [0:0] icmp_ln24_8_fu_484_p2;
wire   [0:0] or_ln23_34_fu_490_p2;
wire   [0:0] select_ln19_38_fu_448_p3;
wire   [2:0] zext_ln22_fu_514_p1;
wire   [2:0] tmp1_fu_524_p2;
wire   [7:0] tmp1_cast_fu_530_p1;
wire   [7:0] empty_135_fu_534_p2;
wire   [3:0] ii_cast_mid1_fu_552_p1;
wire   [3:0] p_cast5_i_i_mid1_fu_555_p2;
wire   [3:0] row_coord_int_mid131_fu_571_p3;
wire   [3:0] row_coord_int_fu_518_p3;
wire   [7:0] col_coord_int_mid139_fu_578_p3;
wire   [7:0] col_coord_int_fu_539_p3;
wire   [0:0] icmp_ln25_fu_603_p2;
wire   [0:0] xor_ln19_fu_598_p2;
wire   [0:0] and_ln19_fu_609_p2;
wire   [0:0] or_ln20_fu_615_p2;
wire   [0:0] select_ln19_39_fu_566_p3;
wire   [3:0] select_ln19_37_fu_560_p3;
wire   [2:0] zext_ln22_7_fu_634_p1;
wire   [2:0] tmp1_mid1_fu_651_p2;
wire   [7:0] tmp1_cast_mid1_fu_657_p1;
wire   [7:0] p_mid1_fu_661_p2;
wire   [3:0] row_coord_int_mid1_fu_644_p3;
wire   [3:0] select_ln19_40_fu_584_p3;
wire   [3:0] select_ln20_32_fu_673_p3;
wire   [7:0] tmp_s_fu_681_p3;
wire   [4:0] tmp_16_fu_693_p3;
wire   [8:0] zext_ln32_fu_689_p1;
wire   [8:0] zext_ln32_34_fu_701_p1;
wire   [8:0] sub_ln32_fu_705_p2;
wire   [7:0] col_coord_int_mid1_fu_666_p3;
wire   [7:0] select_ln19_41_fu_591_p3;
wire   [7:0] select_ln20_33_fu_715_p3;
wire   [9:0] sext_ln20_fu_711_p1;
wire   [9:0] zext_ln32_35_fu_723_p1;
wire   [9:0] add_ln32_fu_727_p2;
wire   [3:0] lshr_ln_fu_737_p4;
wire   [13:0] tmp_52_fu_747_p3;
wire   [3:0] tmp_fu_774_p3;
wire   [4:0] zext_ln33_26_fu_781_p1;
wire   [4:0] zext_ln33_fu_771_p1;
wire   [4:0] sub_ln33_fu_785_p2;
wire   [5:0] sub_ln33_cast_fu_791_p1;
wire   [5:0] zext_ln33_27_fu_795_p1;
wire   [3:0] trunc_ln33_fu_804_p1;
wire   [9:0] tmp_155_cast_fu_808_p3;
wire   [9:0] zext_ln33_28_fu_816_p1;
wire   [15:0] trunc_ln32_fu_829_p1;
wire   [15:0] bitcast_ln32_fu_833_p1;
wire   [5:0] or_ln25_fu_845_p2;
wire   [11:0] tmp_53_fu_850_p3;
wire   [15:0] tmp_84_i_i_fu_862_p4;
wire   [15:0] bitcast_ln32_28_fu_872_p1;
wire   [15:0] tmp_85_i_i_fu_884_p4;
wire   [15:0] bitcast_ln32_29_fu_894_p1;
wire   [15:0] tmp_86_i_i_fu_905_p4;
wire   [15:0] bitcast_ln32_30_fu_915_p1;
wire   [5:0] or_ln25_19_fu_926_p2;
wire   [11:0] tmp_54_fu_931_p3;
wire   [5:0] or_ln25_20_fu_943_p2;
wire   [11:0] tmp_55_fu_948_p3;
wire    ap_CS_fsm_state9;
reg   [4:0] ap_NS_fsm;
wire    ap_block_pp0_stage0_subdone;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 5'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b1 == ap_condition_pp0_exit_iter0_state4) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_subdone))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_subdone))) begin
            if ((1'b1 == ap_condition_pp0_exit_iter0_state4)) begin
                ap_enable_reg_pp0_iter1 <= (1'b1 ^ ap_condition_pp0_exit_iter0_state4);
            end else if ((1'b1 == 1'b1)) begin
                ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
            end
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_subdone))) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            ap_enable_reg_pp0_iter2 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln19_reg_1023 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        ii_reg_236 <= select_ln19_36_reg_1080;
    end else if ((1'b1 == ap_CS_fsm_state2)) begin
        ii_reg_236 <= 2'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln19_reg_1023 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        indvar_flatten47_reg_224 <= add_ln19_7_reg_1075;
    end else if ((1'b1 == ap_CS_fsm_state2)) begin
        indvar_flatten47_reg_224 <= 8'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln19_reg_1023 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        indvar_flatten_reg_248 <= select_ln20_34_reg_1119;
    end else if ((1'b1 == ap_CS_fsm_state2)) begin
        indvar_flatten_reg_248 <= 7'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln19_reg_1023 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        jj_reg_259 <= select_ln20_30_reg_1093;
    end else if ((1'b1 == ap_CS_fsm_state2)) begin
        jj_reg_259 <= 2'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln19_reg_1023_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001))) begin
        kk_0_i_i_reg_271 <= add_ln25_reg_1124;
    end else if ((1'b1 == ap_CS_fsm_state2)) begin
        kk_0_i_i_reg_271 <= 7'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
        add_ln19_7_reg_1075 <= add_ln19_7_fu_508_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (icmp_ln19_fu_407_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        add_ln19_reg_1027 <= add_ln19_fu_413_p2;
        add_ln20_7_reg_1070 <= add_ln20_7_fu_502_p2;
        add_ln20_reg_1057 <= add_ln20_fu_461_p2;
        icmp_ln20_reg_1033 <= icmp_ln20_fu_419_p2;
        or_ln23_33_reg_1050 <= or_ln23_33_fu_456_p2;
        or_ln23_35_reg_1063 <= or_ln23_35_fu_496_p2;
        select_ln19_reg_1045 <= select_ln19_fu_425_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln19_reg_1023 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        add_ln25_reg_1124 <= add_ln25_fu_766_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln19_reg_1023_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001))) begin
        add_ln33_7_reg_1136 <= add_ln33_7_fu_819_p2;
        add_ln33_reg_1129 <= add_ln33_fu_798_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln19_reg_1023 == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001))) begin
        empty_137_reg_1107 <= empty_137_fu_733_p1;
        select_ln20_31_reg_1099 <= select_ln20_31_fu_637_p3;
        select_ln20_reg_1087 <= select_ln20_fu_620_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
        empty_137_reg_1107_pp0_iter1_reg <= empty_137_reg_1107;
        select_ln20_31_reg_1099_pp0_iter1_reg <= select_ln20_31_reg_1099;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state1)) begin
        empty_reg_975 <= empty_fu_287_p1;
        indices_01_read_reg_960 <= indices_01_dout;
        indices_12_read_reg_970 <= indices_12_dout;
        trunc_ln250_reg_965 <= trunc_ln250_fu_282_p1;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        icmp_ln19_reg_1023 <= icmp_ln19_fu_407_p2;
        icmp_ln19_reg_1023_pp0_iter1_reg <= icmp_ln19_reg_1023;
        icmp_ln19_reg_1023_pp0_iter2_reg <= icmp_ln19_reg_1023_pp0_iter1_reg;
        is_padding_reg_1016 <= is_padding_fu_401_p2;
        p_cast5_i_i_reg_1010 <= p_cast5_i_i_fu_361_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        or_ln23_31_reg_1000 <= or_ln23_31_fu_337_p2;
        p_cast_i_i_reg_982 <= p_cast_i_i_fu_304_p1;
        p_cast_reg_994 <= p_cast_fu_318_p2;
        p_mid137_reg_1005 <= p_mid137_fu_343_p2;
        sext_ln22_reg_988 <= sext_ln22_fu_314_p1;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln19_reg_1023 == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001))) begin
        select_ln19_36_reg_1080 <= select_ln19_36_fu_546_p3;
        select_ln20_30_reg_1093 <= select_ln20_30_fu_628_p3;
        select_ln20_34_reg_1119 <= select_ln20_34_fu_760_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (icmp_ln19_reg_1023_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        select_ln33_29_reg_1141 <= select_ln33_29_fu_898_p3;
        select_ln33_30_reg_1146 <= select_ln33_30_fu_919_p3;
    end
end

always @ (*) begin
    if ((icmp_ln19_reg_1023 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state4 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state4 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state9)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln19_reg_1023 == 1'd0) & (1'b0 == ap_block_pp0_stage0))) begin
        ap_phi_mux_ii_phi_fu_240_p4 = select_ln19_36_reg_1080;
    end else begin
        ap_phi_mux_ii_phi_fu_240_p4 = ii_reg_236;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln19_reg_1023 == 1'd0) & (1'b0 == ap_block_pp0_stage0))) begin
        ap_phi_mux_indvar_flatten47_phi_fu_228_p4 = add_ln19_7_reg_1075;
    end else begin
        ap_phi_mux_indvar_flatten47_phi_fu_228_p4 = indvar_flatten47_reg_224;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln19_reg_1023 == 1'd0) & (1'b0 == ap_block_pp0_stage0))) begin
        ap_phi_mux_indvar_flatten_phi_fu_252_p4 = select_ln20_34_reg_1119;
    end else begin
        ap_phi_mux_indvar_flatten_phi_fu_252_p4 = indvar_flatten_reg_248;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln19_reg_1023 == 1'd0) & (1'b0 == ap_block_pp0_stage0))) begin
        ap_phi_mux_jj_phi_fu_263_p4 = select_ln20_30_reg_1093;
    end else begin
        ap_phi_mux_jj_phi_fu_263_p4 = jj_reg_259;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln19_reg_1023_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage1))) begin
        ap_phi_mux_kk_0_i_i_phi_fu_275_p4 = add_ln25_reg_1124;
    end else begin
        ap_phi_mux_kk_0_i_i_phi_fu_275_p4 = kk_0_i_i_reg_271;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state9)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((ap_enable_reg_pp0_iter2 == 1'b1)) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ifmap_vec_address0 = sext_ln33_12_fu_955_p1;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0))) begin
            ifmap_vec_address0 = sext_ln33_fu_857_p1;
        end else begin
            ifmap_vec_address0 = 'bx;
        end
    end else begin
        ifmap_vec_address0 = 'bx;
    end
end

always @ (*) begin
    if ((ap_enable_reg_pp0_iter2 == 1'b1)) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ifmap_vec_address1 = sext_ln33_11_fu_938_p1;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0))) begin
            ifmap_vec_address1 = zext_ln33_29_fu_825_p1;
        end else begin
            ifmap_vec_address1 = 'bx;
        end
    end else begin
        ifmap_vec_address1 = 'bx;
    end
end

always @ (*) begin
    if ((((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_11001)) | ((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
        ifmap_vec_ce0 = 1'b1;
    end else begin
        ifmap_vec_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_11001)) | ((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
        ifmap_vec_ce1 = 1'b1;
    end else begin
        ifmap_vec_ce1 = 1'b0;
    end
end

always @ (*) begin
    if ((ap_enable_reg_pp0_iter2 == 1'b1)) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ifmap_vec_d0 = select_ln33_30_reg_1146;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0))) begin
            ifmap_vec_d0 = select_ln33_28_fu_876_p3;
        end else begin
            ifmap_vec_d0 = 'bx;
        end
    end else begin
        ifmap_vec_d0 = 'bx;
    end
end

always @ (*) begin
    if ((ap_enable_reg_pp0_iter2 == 1'b1)) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ifmap_vec_d1 = select_ln33_29_reg_1141;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0))) begin
            ifmap_vec_d1 = select_ln33_fu_837_p3;
        end else begin
            ifmap_vec_d1 = 'bx;
        end
    end else begin
        ifmap_vec_d1 = 'bx;
    end
end

always @ (*) begin
    if ((((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln19_reg_1023_pp0_iter2_reg == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001)) | ((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (icmp_ln19_reg_1023_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
        ifmap_vec_we0 = 1'b1;
    end else begin
        ifmap_vec_we0 = 1'b0;
    end
end

always @ (*) begin
    if ((((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln19_reg_1023_pp0_iter2_reg == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001)) | ((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (icmp_ln19_reg_1023_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
        ifmap_vec_we1 = 1'b1;
    end else begin
        ifmap_vec_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001)) | ((1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b0 == ap_block_pp0_stage1_11001)) | ((1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage1_11001)) | ((1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
        in_data_ce0 = 1'b1;
    end else begin
        in_data_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_01_blk_n = indices_01_empty_n;
    end else begin
        indices_01_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_01_out_blk_n = indices_01_out_full_n;
    end else begin
        indices_01_out_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((indices_12_out_full_n == 1'b0) | (indices_01_out_full_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_01_out_write = 1'b1;
    end else begin
        indices_01_out_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((indices_12_out_full_n == 1'b0) | (indices_01_out_full_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_01_read = 1'b1;
    end else begin
        indices_01_read = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_12_blk_n = indices_12_empty_n;
    end else begin
        indices_12_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_12_out_blk_n = indices_12_out_full_n;
    end else begin
        indices_12_out_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((indices_12_out_full_n == 1'b0) | (indices_01_out_full_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_12_out_write = 1'b1;
    end else begin
        indices_12_out_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((indices_12_out_full_n == 1'b0) | (indices_01_out_full_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_12_read = 1'b1;
    end else begin
        indices_12_read = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((indices_12_out_full_n == 1'b0) | (indices_01_out_full_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_state2 : begin
            ap_NS_fsm = ap_ST_fsm_pp0_stage0;
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_pp0_stage1 : begin
            if ((~((ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln19_reg_1023 == 1'd1) & (1'b0 == ap_block_pp0_stage1_subdone)) & ~((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b0) & (1'b0 == ap_block_pp0_stage1_subdone)) & (1'b0 == ap_block_pp0_stage1_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if ((((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b0) & (1'b0 == ap_block_pp0_stage1_subdone)) | ((ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln19_reg_1023 == 1'd1) & (1'b0 == ap_block_pp0_stage1_subdone)))) begin
                ap_NS_fsm = ap_ST_fsm_state9;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end
        end
        ap_ST_fsm_state9 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln19_7_fu_508_p2 = (indvar_flatten47_reg_224 + 8'd1);

assign add_ln19_fu_413_p2 = (ap_phi_mux_ii_phi_fu_240_p4 + 2'd1);

assign add_ln20_7_fu_502_p2 = (ap_phi_mux_indvar_flatten_phi_fu_252_p4 + 7'd1);

assign add_ln20_fu_461_p2 = (select_ln19_fu_425_p3 + 2'd1);

assign add_ln22_7_fu_376_p2 = ((sext_ln22_reg_988) + (zext_ln20_fu_372_p1));

assign add_ln22_8_fu_471_p2 = ((sext_ln22_reg_988) + (zext_ln20_7_fu_467_p1));

assign add_ln22_fu_308_p2 = ((j_cast_i_i_fu_292_p1) + (17'd131071));

assign add_ln25_fu_766_p2 = (select_ln20_reg_1087 + 7'd4);

assign add_ln32_fu_727_p2 = ((sext_ln20_fu_711_p1) + (zext_ln32_35_fu_723_p1));

assign add_ln33_7_fu_819_p2 = (tmp_155_cast_fu_808_p3 + zext_ln33_28_fu_816_p1);

assign add_ln33_fu_798_p2 = ((sub_ln33_cast_fu_791_p1) + (zext_ln33_27_fu_795_p1));

assign and_ln19_fu_609_p2 = (xor_ln19_fu_598_p2 & icmp_ln25_fu_603_p2);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_pp0_stage1 = ap_CS_fsm[32'd3];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state9 = ap_CS_fsm[32'd4];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((indices_12_out_full_n == 1'b0) | (indices_01_out_full_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0));
end

assign ap_block_state3_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage1_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage1_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage1_iter2 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign bitcast_ln32_28_fu_872_p1 = tmp_84_i_i_fu_862_p4;

assign bitcast_ln32_29_fu_894_p1 = tmp_85_i_i_fu_884_p4;

assign bitcast_ln32_30_fu_915_p1 = tmp_86_i_i_fu_905_p4;

assign bitcast_ln32_fu_833_p1 = trunc_ln32_fu_829_p1;

assign col_coord_int_fu_539_p3 = ((is_padding_reg_1016[0:0] == 1'b1) ? 8'd0 : empty_135_fu_534_p2);

assign col_coord_int_mid139_fu_578_p3 = ((or_ln23_33_reg_1050[0:0] == 1'b1) ? 8'd0 : p_mid137_reg_1005);

assign col_coord_int_mid1_fu_666_p3 = ((or_ln23_35_reg_1063[0:0] == 1'b1) ? 8'd0 : p_mid1_fu_661_p2);

assign empty_132_fu_298_p2 = ((zext_ln19_fu_295_p1) + (17'd131071));

assign empty_133_fu_356_p2 = ((p_cast_i_i_reg_982) + (ii_cast_i_i_fu_348_p1));

assign empty_134_fu_366_p2 = ((empty_133_fu_356_p2 > 18'd13) ? 1'b1 : 1'b0);

assign empty_135_fu_534_p2 = ((tmp1_cast_fu_530_p1) + (empty_reg_975));

assign empty_137_fu_733_p1 = select_ln20_fu_620_p3[5:0];

assign empty_fu_287_p1 = indices_12_dout[7:0];

assign icmp_ln19_fu_407_p2 = ((ap_phi_mux_indvar_flatten47_phi_fu_228_p4 == 8'd144) ? 1'b1 : 1'b0);

assign icmp_ln20_fu_419_p2 = ((ap_phi_mux_indvar_flatten_phi_fu_252_p4 == 7'd48) ? 1'b1 : 1'b0);

assign icmp_ln24_7_fu_389_p2 = (((add_ln22_7_fu_376_p2) > (18'd13)) ? 1'b1 : 1'b0);

assign icmp_ln24_8_fu_484_p2 = (((add_ln22_8_fu_471_p2) > (18'd13)) ? 1'b1 : 1'b0);

assign icmp_ln24_fu_331_p2 = (((add_ln22_fu_308_p2) > (17'd13)) ? 1'b1 : 1'b0);

assign icmp_ln25_fu_603_p2 = ((ap_phi_mux_kk_0_i_i_phi_fu_275_p4 == 7'd64) ? 1'b1 : 1'b0);

assign ii_cast_fu_352_p1 = ap_phi_mux_ii_phi_fu_240_p4;

assign ii_cast_i_i_fu_348_p1 = ap_phi_mux_ii_phi_fu_240_p4;

assign ii_cast_i_i_mid1_fu_433_p1 = add_ln19_fu_413_p2;

assign ii_cast_mid1_fu_552_p1 = add_ln19_reg_1027;

assign in_data_address0 = sext_ln32_fu_755_p1;

assign indices_01_out_din = indices_01_dout[3:0];

assign indices_12_out_din = indices_12_dout[7:0];

assign is_padding_fu_401_p2 = (or_ln23_fu_395_p2 | empty_134_fu_366_p2);

assign j_cast_i_i_fu_292_p1 = indices_12_read_reg_970;

assign lshr_ln_fu_737_p4 = {{select_ln20_fu_620_p3[5:2]}};

assign or_ln20_fu_615_p2 = (icmp_ln20_reg_1033 | and_ln19_fu_609_p2);

assign or_ln23_31_fu_337_p2 = (tmp_49_fu_323_p3 | icmp_ln24_fu_331_p2);

assign or_ln23_33_fu_456_p2 = (p_mid113_fu_442_p2 | or_ln23_31_reg_1000);

assign or_ln23_34_fu_490_p2 = (tmp_51_fu_476_p3 | icmp_ln24_8_fu_484_p2);

assign or_ln23_35_fu_496_p2 = (select_ln19_38_fu_448_p3 | or_ln23_34_fu_490_p2);

assign or_ln23_fu_395_p2 = (tmp_50_fu_381_p3 | icmp_ln24_7_fu_389_p2);

assign or_ln25_19_fu_926_p2 = (empty_137_reg_1107_pp0_iter1_reg | 6'd2);

assign or_ln25_20_fu_943_p2 = (empty_137_reg_1107_pp0_iter1_reg | 6'd3);

assign or_ln25_fu_845_p2 = (empty_137_reg_1107_pp0_iter1_reg | 6'd1);

assign p_cast5_i_i_fu_361_p2 = (p_cast_reg_994 + ii_cast_fu_352_p1);

assign p_cast5_i_i_mid1_fu_555_p2 = (p_cast_reg_994 + ii_cast_mid1_fu_552_p1);

assign p_cast_fu_318_p2 = ((trunc_ln250_reg_965) + (4'd15));

assign p_cast_i_i_fu_304_p1 = (empty_132_fu_298_p2);

assign p_mid111_fu_437_p2 = ((p_cast_i_i_reg_982) + (ii_cast_i_i_mid1_fu_433_p1));

assign p_mid113_fu_442_p2 = ((p_mid111_fu_437_p2 > 18'd13) ? 1'b1 : 1'b0);

assign p_mid137_fu_343_p2 = ((empty_reg_975) + (8'd255));

assign p_mid1_fu_661_p2 = ((tmp1_cast_mid1_fu_657_p1) + (empty_reg_975));

assign row_coord_int_fu_518_p3 = ((is_padding_reg_1016[0:0] == 1'b1) ? 4'd0 : p_cast5_i_i_reg_1010);

assign row_coord_int_mid131_fu_571_p3 = ((or_ln23_33_reg_1050[0:0] == 1'b1) ? 4'd0 : p_cast5_i_i_mid1_fu_555_p2);

assign row_coord_int_mid1_fu_644_p3 = ((or_ln23_35_reg_1063[0:0] == 1'b1) ? 4'd0 : select_ln19_37_fu_560_p3);

assign select_ln19_36_fu_546_p3 = ((icmp_ln20_reg_1033[0:0] == 1'b1) ? add_ln19_reg_1027 : ii_reg_236);

assign select_ln19_37_fu_560_p3 = ((icmp_ln20_reg_1033[0:0] == 1'b1) ? p_cast5_i_i_mid1_fu_555_p2 : p_cast5_i_i_reg_1010);

assign select_ln19_38_fu_448_p3 = ((icmp_ln20_fu_419_p2[0:0] == 1'b1) ? p_mid113_fu_442_p2 : empty_134_fu_366_p2);

assign select_ln19_39_fu_566_p3 = ((icmp_ln20_reg_1033[0:0] == 1'b1) ? or_ln23_33_reg_1050 : is_padding_reg_1016);

assign select_ln19_40_fu_584_p3 = ((icmp_ln20_reg_1033[0:0] == 1'b1) ? row_coord_int_mid131_fu_571_p3 : row_coord_int_fu_518_p3);

assign select_ln19_41_fu_591_p3 = ((icmp_ln20_reg_1033[0:0] == 1'b1) ? col_coord_int_mid139_fu_578_p3 : col_coord_int_fu_539_p3);

assign select_ln19_fu_425_p3 = ((icmp_ln20_fu_419_p2[0:0] == 1'b1) ? 2'd0 : ap_phi_mux_jj_phi_fu_263_p4);

assign select_ln20_30_fu_628_p3 = ((and_ln19_fu_609_p2[0:0] == 1'b1) ? add_ln20_reg_1057 : select_ln19_reg_1045);

assign select_ln20_31_fu_637_p3 = ((and_ln19_fu_609_p2[0:0] == 1'b1) ? or_ln23_35_reg_1063 : select_ln19_39_fu_566_p3);

assign select_ln20_32_fu_673_p3 = ((and_ln19_fu_609_p2[0:0] == 1'b1) ? row_coord_int_mid1_fu_644_p3 : select_ln19_40_fu_584_p3);

assign select_ln20_33_fu_715_p3 = ((and_ln19_fu_609_p2[0:0] == 1'b1) ? col_coord_int_mid1_fu_666_p3 : select_ln19_41_fu_591_p3);

assign select_ln20_34_fu_760_p3 = ((icmp_ln20_reg_1033[0:0] == 1'b1) ? 7'd1 : add_ln20_7_reg_1070);

assign select_ln20_fu_620_p3 = ((or_ln20_fu_615_p2[0:0] == 1'b1) ? 7'd0 : ap_phi_mux_kk_0_i_i_phi_fu_275_p4);

assign select_ln33_28_fu_876_p3 = ((select_ln20_31_reg_1099_pp0_iter1_reg[0:0] == 1'b1) ? 16'd0 : bitcast_ln32_28_fu_872_p1);

assign select_ln33_29_fu_898_p3 = ((select_ln20_31_reg_1099_pp0_iter1_reg[0:0] == 1'b1) ? 16'd0 : bitcast_ln32_29_fu_894_p1);

assign select_ln33_30_fu_919_p3 = ((select_ln20_31_reg_1099_pp0_iter1_reg[0:0] == 1'b1) ? 16'd0 : bitcast_ln32_30_fu_915_p1);

assign select_ln33_fu_837_p3 = ((select_ln20_31_reg_1099_pp0_iter1_reg[0:0] == 1'b1) ? 16'd0 : bitcast_ln32_fu_833_p1);

assign sext_ln20_fu_711_p1 = (sub_ln32_fu_705_p2);

assign sext_ln22_fu_314_p1 = add_ln22_fu_308_p2;

assign sext_ln32_fu_755_p1 = (tmp_52_fu_747_p3);

assign sext_ln33_11_fu_938_p1 = (tmp_54_fu_931_p3);

assign sext_ln33_12_fu_955_p1 = (tmp_55_fu_948_p3);

assign sext_ln33_fu_857_p1 = (tmp_53_fu_850_p3);

assign sub_ln32_fu_705_p2 = (zext_ln32_fu_689_p1 - zext_ln32_34_fu_701_p1);

assign sub_ln33_cast_fu_791_p1 = (sub_ln33_fu_785_p2);

assign sub_ln33_fu_785_p2 = (zext_ln33_26_fu_781_p1 - zext_ln33_fu_771_p1);

assign tmp1_cast_fu_530_p1 = (tmp1_fu_524_p2);

assign tmp1_cast_mid1_fu_657_p1 = (tmp1_mid1_fu_651_p2);

assign tmp1_fu_524_p2 = ((zext_ln22_fu_514_p1) + (3'd7));

assign tmp1_mid1_fu_651_p2 = ((zext_ln22_7_fu_634_p1) + (3'd7));

assign tmp_155_cast_fu_808_p3 = {{trunc_ln33_fu_804_p1}, {6'd0}};

assign tmp_16_fu_693_p3 = {{select_ln20_32_fu_673_p3}, {1'd0}};

assign tmp_49_fu_323_p3 = add_ln22_fu_308_p2[32'd16];

assign tmp_50_fu_381_p3 = add_ln22_7_fu_376_p2[32'd17];

assign tmp_51_fu_476_p3 = add_ln22_8_fu_471_p2[32'd17];

assign tmp_52_fu_747_p3 = {{add_ln32_fu_727_p2}, {lshr_ln_fu_737_p4}};

assign tmp_53_fu_850_p3 = {{add_ln33_reg_1129}, {or_ln25_fu_845_p2}};

assign tmp_54_fu_931_p3 = {{add_ln33_reg_1129}, {or_ln25_19_fu_926_p2}};

assign tmp_55_fu_948_p3 = {{add_ln33_reg_1129}, {or_ln25_20_fu_943_p2}};

assign tmp_84_i_i_fu_862_p4 = {{in_data_q0[31:16]}};

assign tmp_85_i_i_fu_884_p4 = {{in_data_q0[47:32]}};

assign tmp_86_i_i_fu_905_p4 = {{in_data_q0[63:48]}};

assign tmp_fu_774_p3 = {{select_ln19_36_reg_1080}, {2'd0}};

assign tmp_s_fu_681_p3 = {{select_ln20_32_fu_673_p3}, {4'd0}};

assign trunc_ln250_fu_282_p1 = indices_01_dout[3:0];

assign trunc_ln32_fu_829_p1 = in_data_q0[15:0];

assign trunc_ln33_fu_804_p1 = add_ln33_fu_798_p2[3:0];

assign xor_ln19_fu_598_p2 = (icmp_ln20_reg_1033 ^ 1'd1);

assign zext_ln19_fu_295_p1 = indices_01_read_reg_960;

assign zext_ln20_7_fu_467_p1 = add_ln20_fu_461_p2;

assign zext_ln20_fu_372_p1 = ap_phi_mux_jj_phi_fu_263_p4;

assign zext_ln22_7_fu_634_p1 = add_ln20_reg_1057;

assign zext_ln22_fu_514_p1 = jj_reg_259;

assign zext_ln32_34_fu_701_p1 = tmp_16_fu_693_p3;

assign zext_ln32_35_fu_723_p1 = select_ln20_33_fu_715_p3;

assign zext_ln32_fu_689_p1 = tmp_s_fu_681_p3;

assign zext_ln33_26_fu_781_p1 = tmp_fu_774_p3;

assign zext_ln33_27_fu_795_p1 = select_ln20_30_reg_1093;

assign zext_ln33_28_fu_816_p1 = select_ln20_reg_1087;

assign zext_ln33_29_fu_825_p1 = add_ln33_7_reg_1136;

assign zext_ln33_fu_771_p1 = select_ln19_36_reg_1080;

endmodule //td_fused_top_tdf11_readInputs75
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf12_13 (
        in_data_address0,
        in_data_ce0,
        in_data_d0,
        in_data_q0,
        in_data_we0,
        in_data_address1,
        in_data_ce1,
        in_data_d1,
        in_data_q1,
        in_data_we1,
        out_data_address0,
        out_data_ce0,
        out_data_d0,
        out_data_q0,
        out_data_we0,
        out_data_address1,
        out_data_ce1,
        out_data_d1,
        out_data_q1,
        out_data_we1,
        filter_data_address0,
        filter_data_ce0,
        filter_data_d0,
        filter_data_q0,
        filter_data_we0,
        filter_data_address1,
        filter_data_ce1,
        filter_data_d1,
        filter_data_q1,
        filter_data_we1,
        adjustments_address0,
        adjustments_ce0,
        adjustments_d0,
        adjustments_q0,
        adjustments_we0,
        adjustments_address1,
        adjustments_ce1,
        adjustments_d1,
        adjustments_q1,
        adjustments_we1,
        ap_clk,
        ap_rst,
        in_data_empty_n,
        in_data_read,
        out_data_full_n,
        out_data_write,
        ap_start,
        ap_done,
        ap_ready,
        ap_idle,
        ap_continue
);


output  [12:0] in_data_address0;
output   in_data_ce0;
output  [63:0] in_data_d0;
input  [63:0] in_data_q0;
output   in_data_we0;
output  [12:0] in_data_address1;
output   in_data_ce1;
output  [63:0] in_data_d1;
input  [63:0] in_data_q1;
output   in_data_we1;
output  [15:0] out_data_address0;
output   out_data_ce0;
output  [63:0] out_data_d0;
input  [63:0] out_data_q0;
output   out_data_we0;
output  [15:0] out_data_address1;
output   out_data_ce1;
output  [63:0] out_data_d1;
input  [63:0] out_data_q1;
output   out_data_we1;
output  [16:0] filter_data_address0;
output   filter_data_ce0;
output  [15:0] filter_data_d0;
input  [15:0] filter_data_q0;
output   filter_data_we0;
output  [16:0] filter_data_address1;
output   filter_data_ce1;
output  [15:0] filter_data_d1;
input  [15:0] filter_data_q1;
output   filter_data_we1;
output  [9:0] adjustments_address0;
output   adjustments_ce0;
output  [47:0] adjustments_d0;
input  [47:0] adjustments_q0;
output   adjustments_we0;
output  [9:0] adjustments_address1;
output   adjustments_ce1;
output  [47:0] adjustments_d1;
input  [47:0] adjustments_q1;
output   adjustments_we1;
input   ap_clk;
input   ap_rst;
input   in_data_empty_n;
output   in_data_read;
input   out_data_full_n;
output   out_data_write;
input   ap_start;
output   ap_done;
output   ap_ready;
output   ap_idle;
input   ap_continue;

reg ap_done;
reg ap_ready;
reg ap_idle;

wire   [12:0] dataflow_in_loop_TOP_LOOP76_U0_in_data_address0;
wire    dataflow_in_loop_TOP_LOOP76_U0_in_data_ce0;
wire   [63:0] dataflow_in_loop_TOP_LOOP76_U0_in_data_d0;
wire    dataflow_in_loop_TOP_LOOP76_U0_in_data_we0;
wire   [12:0] dataflow_in_loop_TOP_LOOP76_U0_in_data_address1;
wire    dataflow_in_loop_TOP_LOOP76_U0_in_data_ce1;
wire   [63:0] dataflow_in_loop_TOP_LOOP76_U0_in_data_d1;
wire    dataflow_in_loop_TOP_LOOP76_U0_in_data_we1;
wire   [16:0] dataflow_in_loop_TOP_LOOP76_U0_filter_data_address0;
wire    dataflow_in_loop_TOP_LOOP76_U0_filter_data_ce0;
wire   [15:0] dataflow_in_loop_TOP_LOOP76_U0_filter_data_d0;
wire    dataflow_in_loop_TOP_LOOP76_U0_filter_data_we0;
wire   [16:0] dataflow_in_loop_TOP_LOOP76_U0_filter_data_address1;
wire    dataflow_in_loop_TOP_LOOP76_U0_filter_data_ce1;
wire   [15:0] dataflow_in_loop_TOP_LOOP76_U0_filter_data_d1;
wire    dataflow_in_loop_TOP_LOOP76_U0_filter_data_we1;
wire   [9:0] dataflow_in_loop_TOP_LOOP76_U0_adjustments_address0;
wire    dataflow_in_loop_TOP_LOOP76_U0_adjustments_ce0;
wire   [47:0] dataflow_in_loop_TOP_LOOP76_U0_adjustments_d0;
wire    dataflow_in_loop_TOP_LOOP76_U0_adjustments_we0;
wire   [9:0] dataflow_in_loop_TOP_LOOP76_U0_adjustments_address1;
wire    dataflow_in_loop_TOP_LOOP76_U0_adjustments_ce1;
wire   [47:0] dataflow_in_loop_TOP_LOOP76_U0_adjustments_d1;
wire    dataflow_in_loop_TOP_LOOP76_U0_adjustments_we1;
wire   [15:0] dataflow_in_loop_TOP_LOOP76_U0_out_data_address0;
wire    dataflow_in_loop_TOP_LOOP76_U0_out_data_ce0;
wire   [63:0] dataflow_in_loop_TOP_LOOP76_U0_out_data_d0;
wire    dataflow_in_loop_TOP_LOOP76_U0_out_data_we0;
wire   [15:0] dataflow_in_loop_TOP_LOOP76_U0_out_data_address1;
wire    dataflow_in_loop_TOP_LOOP76_U0_out_data_ce1;
wire   [63:0] dataflow_in_loop_TOP_LOOP76_U0_out_data_d1;
wire    dataflow_in_loop_TOP_LOOP76_U0_out_data_we1;
wire    dataflow_in_loop_TOP_LOOP76_U0_ap_start;
wire    dataflow_in_loop_TOP_LOOP76_U0_in_data_read;
wire    dataflow_in_loop_TOP_LOOP76_U0_out_data_write;
wire    dataflow_in_loop_TOP_LOOP76_U0_ap_done;
wire    dataflow_in_loop_TOP_LOOP76_U0_ap_ready;
wire    dataflow_in_loop_TOP_LOOP76_U0_ap_idle;
reg    dataflow_in_loop_TOP_LOOP76_U0_ap_continue;
wire    dataflow_in_loop_TOP_LOOP76_U0_in_data_full_n;
wire    dataflow_in_loop_TOP_LOOP76_U0_in_data_write;
wire    ap_sync_continue;
wire    ap_sync_done;
wire    ap_sync_ready;
reg   [17:0] loop_dataflow_input_count;
reg   [17:0] loop_dataflow_output_count;
wire   [17:0] bound_minus_1;
wire    dataflow_in_loop_TOP_LOOP76_U0_start_full_n;
wire    dataflow_in_loop_TOP_LOOP76_U0_start_write;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 loop_dataflow_input_count = 18'd0;
#0 loop_dataflow_output_count = 18'd0;
end

td_fused_top_dataflow_in_loop_TOP_LOOP76 dataflow_in_loop_TOP_LOOP76_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .in_data_address0(dataflow_in_loop_TOP_LOOP76_U0_in_data_address0),
    .in_data_ce0(dataflow_in_loop_TOP_LOOP76_U0_in_data_ce0),
    .in_data_d0(dataflow_in_loop_TOP_LOOP76_U0_in_data_d0),
    .in_data_q0(in_data_q0),
    .in_data_we0(dataflow_in_loop_TOP_LOOP76_U0_in_data_we0),
    .in_data_address1(dataflow_in_loop_TOP_LOOP76_U0_in_data_address1),
    .in_data_ce1(dataflow_in_loop_TOP_LOOP76_U0_in_data_ce1),
    .in_data_d1(dataflow_in_loop_TOP_LOOP76_U0_in_data_d1),
    .in_data_q1(64'd0),
    .in_data_we1(dataflow_in_loop_TOP_LOOP76_U0_in_data_we1),
    .filter_data_address0(dataflow_in_loop_TOP_LOOP76_U0_filter_data_address0),
    .filter_data_ce0(dataflow_in_loop_TOP_LOOP76_U0_filter_data_ce0),
    .filter_data_d0(dataflow_in_loop_TOP_LOOP76_U0_filter_data_d0),
    .filter_data_q0(filter_data_q0),
    .filter_data_we0(dataflow_in_loop_TOP_LOOP76_U0_filter_data_we0),
    .filter_data_address1(dataflow_in_loop_TOP_LOOP76_U0_filter_data_address1),
    .filter_data_ce1(dataflow_in_loop_TOP_LOOP76_U0_filter_data_ce1),
    .filter_data_d1(dataflow_in_loop_TOP_LOOP76_U0_filter_data_d1),
    .filter_data_q1(16'd0),
    .filter_data_we1(dataflow_in_loop_TOP_LOOP76_U0_filter_data_we1),
    .adjustments_address0(dataflow_in_loop_TOP_LOOP76_U0_adjustments_address0),
    .adjustments_ce0(dataflow_in_loop_TOP_LOOP76_U0_adjustments_ce0),
    .adjustments_d0(dataflow_in_loop_TOP_LOOP76_U0_adjustments_d0),
    .adjustments_q0(adjustments_q0),
    .adjustments_we0(dataflow_in_loop_TOP_LOOP76_U0_adjustments_we0),
    .adjustments_address1(dataflow_in_loop_TOP_LOOP76_U0_adjustments_address1),
    .adjustments_ce1(dataflow_in_loop_TOP_LOOP76_U0_adjustments_ce1),
    .adjustments_d1(dataflow_in_loop_TOP_LOOP76_U0_adjustments_d1),
    .adjustments_q1(48'd0),
    .adjustments_we1(dataflow_in_loop_TOP_LOOP76_U0_adjustments_we1),
    .out_data_address0(dataflow_in_loop_TOP_LOOP76_U0_out_data_address0),
    .out_data_ce0(dataflow_in_loop_TOP_LOOP76_U0_out_data_ce0),
    .out_data_d0(dataflow_in_loop_TOP_LOOP76_U0_out_data_d0),
    .out_data_q0(64'd0),
    .out_data_we0(dataflow_in_loop_TOP_LOOP76_U0_out_data_we0),
    .out_data_address1(dataflow_in_loop_TOP_LOOP76_U0_out_data_address1),
    .out_data_ce1(dataflow_in_loop_TOP_LOOP76_U0_out_data_ce1),
    .out_data_d1(dataflow_in_loop_TOP_LOOP76_U0_out_data_d1),
    .out_data_q1(64'd0),
    .out_data_we1(dataflow_in_loop_TOP_LOOP76_U0_out_data_we1),
    .ap_start(dataflow_in_loop_TOP_LOOP76_U0_ap_start),
    .in_data_empty_n(1'b0),
    .in_data_read(dataflow_in_loop_TOP_LOOP76_U0_in_data_read),
    .out_data_full_n(out_data_full_n),
    .out_data_write(dataflow_in_loop_TOP_LOOP76_U0_out_data_write),
    .ap_done(dataflow_in_loop_TOP_LOOP76_U0_ap_done),
    .ap_ready(dataflow_in_loop_TOP_LOOP76_U0_ap_ready),
    .ap_idle(dataflow_in_loop_TOP_LOOP76_U0_ap_idle),
    .ap_continue(dataflow_in_loop_TOP_LOOP76_U0_ap_continue)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        loop_dataflow_input_count <= 18'd0;
    end else begin
        if ((~(loop_dataflow_input_count == bound_minus_1) & (dataflow_in_loop_TOP_LOOP76_U0_ap_ready == 1'b1) & (ap_start == 1'b1))) begin
            loop_dataflow_input_count <= (loop_dataflow_input_count + 18'd1);
        end else if (((dataflow_in_loop_TOP_LOOP76_U0_ap_ready == 1'b1) & (loop_dataflow_input_count == bound_minus_1) & (ap_start == 1'b1))) begin
            loop_dataflow_input_count <= 18'd0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        loop_dataflow_output_count <= 18'd0;
    end else begin
        if ((~(loop_dataflow_output_count == bound_minus_1) & (dataflow_in_loop_TOP_LOOP76_U0_ap_continue == 1'b1) & (dataflow_in_loop_TOP_LOOP76_U0_ap_done == 1'b1))) begin
            loop_dataflow_output_count <= (loop_dataflow_output_count + 18'd1);
        end else if (((dataflow_in_loop_TOP_LOOP76_U0_ap_continue == 1'b1) & (dataflow_in_loop_TOP_LOOP76_U0_ap_done == 1'b1) & (loop_dataflow_output_count == bound_minus_1))) begin
            loop_dataflow_output_count <= 18'd0;
        end
    end
end

always @ (*) begin
    if (((dataflow_in_loop_TOP_LOOP76_U0_ap_done == 1'b1) & (loop_dataflow_output_count == bound_minus_1))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = 1'b0;
    end
end

always @ (*) begin
    if (((dataflow_in_loop_TOP_LOOP76_U0_ap_idle == 1'b1) & (loop_dataflow_output_count == 18'd0) & (ap_start == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((dataflow_in_loop_TOP_LOOP76_U0_ap_ready == 1'b1) & (loop_dataflow_input_count == bound_minus_1) & (ap_start == 1'b1))) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((~(loop_dataflow_output_count == bound_minus_1) | (ap_continue == 1'b1))) begin
        dataflow_in_loop_TOP_LOOP76_U0_ap_continue = 1'b1;
    end else begin
        dataflow_in_loop_TOP_LOOP76_U0_ap_continue = 1'b0;
    end
end

assign adjustments_address0 = dataflow_in_loop_TOP_LOOP76_U0_adjustments_address0;

assign adjustments_address1 = 10'd0;

assign adjustments_ce0 = dataflow_in_loop_TOP_LOOP76_U0_adjustments_ce0;

assign adjustments_ce1 = 1'b0;

assign adjustments_d0 = 48'd0;

assign adjustments_d1 = 48'd0;

assign adjustments_we0 = 1'b0;

assign adjustments_we1 = 1'b0;

assign ap_sync_continue = ap_continue;

assign ap_sync_done = dataflow_in_loop_TOP_LOOP76_U0_ap_done;

assign ap_sync_ready = dataflow_in_loop_TOP_LOOP76_U0_ap_ready;

assign bound_minus_1 = (18'd196000 - 18'd1);

assign dataflow_in_loop_TOP_LOOP76_U0_ap_start = ap_start;

assign dataflow_in_loop_TOP_LOOP76_U0_in_data_full_n = in_data_empty_n;

assign dataflow_in_loop_TOP_LOOP76_U0_in_data_write = 1'b0;

assign dataflow_in_loop_TOP_LOOP76_U0_start_full_n = 1'b1;

assign dataflow_in_loop_TOP_LOOP76_U0_start_write = 1'b0;

assign filter_data_address0 = dataflow_in_loop_TOP_LOOP76_U0_filter_data_address0;

assign filter_data_address1 = 17'd0;

assign filter_data_ce0 = dataflow_in_loop_TOP_LOOP76_U0_filter_data_ce0;

assign filter_data_ce1 = 1'b0;

assign filter_data_d0 = 16'd0;

assign filter_data_d1 = 16'd0;

assign filter_data_we0 = 1'b0;

assign filter_data_we1 = 1'b0;

assign in_data_address0 = dataflow_in_loop_TOP_LOOP76_U0_in_data_address0;

assign in_data_address1 = 13'd0;

assign in_data_ce0 = dataflow_in_loop_TOP_LOOP76_U0_in_data_ce0;

assign in_data_ce1 = 1'b0;

assign in_data_d0 = 64'd0;

assign in_data_d1 = 64'd0;

assign in_data_read = dataflow_in_loop_TOP_LOOP76_U0_in_data_write;

assign in_data_we0 = 1'b0;

assign in_data_we1 = 1'b0;

assign out_data_address0 = 16'd0;

assign out_data_address1 = dataflow_in_loop_TOP_LOOP76_U0_out_data_address1;

assign out_data_ce0 = 1'b0;

assign out_data_ce1 = dataflow_in_loop_TOP_LOOP76_U0_out_data_ce1;

assign out_data_d0 = 64'd0;

assign out_data_d1 = dataflow_in_loop_TOP_LOOP76_U0_out_data_d1;

assign out_data_we0 = 1'b0;

assign out_data_we1 = dataflow_in_loop_TOP_LOOP76_U0_out_data_we1;

assign out_data_write = dataflow_in_loop_TOP_LOOP76_U0_out_data_write;

endmodule //td_fused_top_tdf12_13
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf12_accum_1 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        accum_in_0_address0,
        accum_in_0_ce0,
        accum_in_0_q0,
        accum_in_0_address1,
        accum_in_0_ce1,
        accum_in_0_q1,
        accum_out_address0,
        accum_out_ce0,
        accum_out_we0,
        accum_out_d0,
        accum_out_address1,
        accum_out_ce1,
        accum_out_we1,
        accum_out_d1
);

parameter    ap_ST_fsm_state1 = 8'd1;
parameter    ap_ST_fsm_pp0_stage0 = 8'd2;
parameter    ap_ST_fsm_pp0_stage1 = 8'd4;
parameter    ap_ST_fsm_pp0_stage2 = 8'd8;
parameter    ap_ST_fsm_pp0_stage3 = 8'd16;
parameter    ap_ST_fsm_state12 = 8'd32;
parameter    ap_ST_fsm_state13 = 8'd64;
parameter    ap_ST_fsm_state14 = 8'd128;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [6:0] accum_in_0_address0;
output   accum_in_0_ce0;
input  [15:0] accum_in_0_q0;
output  [6:0] accum_in_0_address1;
output   accum_in_0_ce1;
input  [15:0] accum_in_0_q1;
output  [2:0] accum_out_address0;
output   accum_out_ce0;
output   accum_out_we0;
output  [15:0] accum_out_d0;
output  [2:0] accum_out_address1;
output   accum_out_ce1;
output   accum_out_we1;
output  [15:0] accum_out_d1;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg[6:0] accum_in_0_address0;
reg accum_in_0_ce0;
reg[6:0] accum_in_0_address1;
reg accum_in_0_ce1;
reg accum_out_ce0;
reg accum_out_we0;
reg accum_out_ce1;
reg accum_out_we1;

reg    ap_done_reg;
  reg   [7:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg   [7:0] x_reg_170;
reg   [15:0] psum_7_08_reg_182;
reg   [15:0] psum_6_07_reg_194;
reg   [15:0] psum_5_06_reg_206;
reg   [15:0] psum_4_05_reg_218;
reg   [15:0] psum_3_04_reg_230;
reg   [15:0] psum_2_03_reg_242;
reg   [15:0] psum_1_02_reg_254;
reg   [15:0] psum_0_01_reg_266;
wire   [0:0] tmp_fu_323_p3;
reg   [0:0] tmp_reg_494;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state6_pp0_stage0_iter1;
wire    ap_block_state10_pp0_stage0_iter2;
wire    ap_block_pp0_stage0_11001;
reg   [0:0] tmp_reg_494_pp0_iter1_reg;
reg   [0:0] tmp_reg_494_pp0_iter2_reg;
wire   [6:0] trunc_ln25_fu_336_p1;
reg   [6:0] trunc_ln25_reg_498;
reg   [15:0] accum_in_0_load_reg_518;
wire    ap_CS_fsm_pp0_stage1;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_state3_pp0_stage1_iter0;
wire    ap_block_state7_pp0_stage1_iter1;
wire    ap_block_state11_pp0_stage1_iter2;
wire    ap_block_pp0_stage1_11001;
reg   [15:0] accum_in_0_load_58_reg_523;
reg   [15:0] accum_in_0_load_59_reg_538;
wire    ap_CS_fsm_pp0_stage2;
wire    ap_block_state4_pp0_stage2_iter0;
wire    ap_block_state8_pp0_stage2_iter1;
wire    ap_block_pp0_stage2_11001;
reg   [15:0] accum_in_0_load_60_reg_543;
wire   [7:0] add_ln25_fu_391_p2;
reg   [7:0] add_ln25_reg_558;
wire    ap_CS_fsm_pp0_stage3;
wire    ap_block_state5_pp0_stage3_iter0;
wire    ap_block_state9_pp0_stage3_iter1;
wire    ap_block_pp0_stage3_11001;
reg   [15:0] accum_in_0_load_61_reg_563;
reg   [15:0] accum_in_0_load_62_reg_568;
reg   [15:0] accum_in_0_load_63_reg_583;
reg    ap_enable_reg_pp0_iter1;
reg   [15:0] accum_in_0_load_64_reg_588;
wire   [15:0] grp_fu_307_p2;
wire   [15:0] grp_fu_312_p2;
reg    ap_enable_reg_pp0_iter2;
wire   [3:0] add_ln33_fu_434_p2;
wire    ap_CS_fsm_state13;
wire   [0:0] tmp_48_fu_417_p3;
reg    ap_block_state1;
wire    ap_block_pp0_stage2_subdone;
reg    ap_condition_pp0_exit_iter0_state4;
wire    ap_block_pp0_stage3_subdone;
wire    ap_block_pp0_stage1_subdone;
reg   [7:0] ap_phi_mux_x_phi_fu_174_p4;
wire    ap_block_pp0_stage0;
wire   [15:0] ap_phi_mux_psum_7_08_phi_fu_186_p4;
wire    ap_block_pp0_stage1;
wire   [15:0] ap_phi_mux_psum_6_07_phi_fu_198_p4;
wire   [15:0] ap_phi_mux_psum_5_06_phi_fu_210_p4;
wire   [15:0] ap_phi_mux_psum_4_05_phi_fu_222_p4;
wire   [15:0] ap_phi_mux_psum_3_04_phi_fu_234_p4;
wire    ap_block_pp0_stage3;
wire   [15:0] ap_phi_mux_psum_2_03_phi_fu_246_p4;
wire    ap_block_pp0_stage2;
reg   [3:0] q_reg_278;
wire    ap_CS_fsm_state12;
reg   [15:0] ap_phi_mux_phi_ln45_phi_fu_292_p8;
wire   [2:0] trunc_ln33_fu_430_p1;
wire   [63:0] zext_ln25_fu_331_p1;
wire   [63:0] zext_ln29_fu_346_p1;
wire   [63:0] zext_ln29_19_fu_356_p1;
wire   [63:0] zext_ln29_20_fu_366_p1;
wire   [63:0] zext_ln29_21_fu_376_p1;
wire   [63:0] zext_ln29_22_fu_386_p1;
wire   [63:0] zext_ln29_23_fu_402_p1;
wire   [63:0] zext_ln29_24_fu_412_p1;
wire   [63:0] zext_ln33_fu_425_p1;
wire   [63:0] zext_ln33_4_fu_446_p1;
reg   [15:0] grp_fu_307_p0;
reg   [15:0] grp_fu_307_p1;
reg   [15:0] grp_fu_312_p0;
reg   [15:0] grp_fu_312_p1;
wire   [6:0] or_ln29_fu_340_p2;
wire   [6:0] or_ln29_19_fu_351_p2;
wire   [6:0] or_ln29_20_fu_361_p2;
wire   [6:0] or_ln29_21_fu_371_p2;
wire   [6:0] or_ln29_22_fu_381_p2;
wire   [6:0] or_ln29_23_fu_397_p2;
wire   [6:0] or_ln29_24_fu_407_p2;
wire   [2:0] or_ln33_fu_440_p2;
wire   [0:0] icmp_ln45_fu_451_p2;
wire   [0:0] icmp_ln45_7_fu_465_p2;
wire   [15:0] select_ln45_fu_457_p3;
wire   [0:0] icmp_ln45_8_fu_479_p2;
wire   [15:0] select_ln45_7_fu_471_p3;
wire    ap_CS_fsm_state14;
reg   [7:0] ap_NS_fsm;
wire    ap_block_pp0_stage0_subdone;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
reg    ap_condition_517;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 8'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
end

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U775(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(grp_fu_307_p0),
    .din1(grp_fu_307_p1),
    .dout(grp_fu_307_p2)
);

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U776(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(grp_fu_312_p0),
    .din1(grp_fu_312_p1),
    .dout(grp_fu_312_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state14)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage2_subdone) & (1'b1 == ap_condition_pp0_exit_iter0_state4) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage3_subdone) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b0)) | ((1'b0 == ap_block_pp0_stage3_subdone) & (1'b1 == ap_CS_fsm_pp0_stage3)))) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end else if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter2 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state12)) begin
        q_reg_278 <= 4'd0;
    end else if (((tmp_48_fu_417_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state13))) begin
        q_reg_278 <= add_ln33_fu_434_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (tmp_reg_494 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        x_reg_170 <= add_ln25_reg_558;
    end else if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        x_reg_170 <= 8'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage1_11001) & (tmp_reg_494 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
        accum_in_0_load_58_reg_523 <= accum_in_0_q0;
        accum_in_0_load_reg_518 <= accum_in_0_q1;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage2_11001) & (tmp_reg_494 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage2) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
        accum_in_0_load_59_reg_538 <= accum_in_0_q1;
        accum_in_0_load_60_reg_543 <= accum_in_0_q0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage3_11001) & (tmp_reg_494 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage3) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
        accum_in_0_load_61_reg_563 <= accum_in_0_q1;
        accum_in_0_load_62_reg_568 <= accum_in_0_q0;
        add_ln25_reg_558 <= add_ln25_fu_391_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (tmp_reg_494 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        accum_in_0_load_63_reg_583 <= accum_in_0_q1;
        accum_in_0_load_64_reg_588 <= accum_in_0_q0;
    end
end

always @ (posedge ap_clk) begin
    if (((tmp_reg_494_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage2_11001) & (1'b1 == ap_CS_fsm_pp0_stage2) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        psum_0_01_reg_266 <= grp_fu_307_p2;
        psum_1_02_reg_254 <= grp_fu_312_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((tmp_reg_494_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage3_11001) & (1'b1 == ap_CS_fsm_pp0_stage3) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        psum_2_03_reg_242 <= grp_fu_307_p2;
        psum_3_04_reg_230 <= grp_fu_312_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((tmp_reg_494_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        psum_4_05_reg_218 <= grp_fu_307_p2;
        psum_5_06_reg_206 <= grp_fu_312_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((tmp_reg_494_pp0_iter2_reg == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
        psum_6_07_reg_194 <= grp_fu_307_p2;
        psum_7_08_reg_182 <= grp_fu_312_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_reg_494 <= ap_phi_mux_x_phi_fu_174_p4[32'd7];
        tmp_reg_494_pp0_iter1_reg <= tmp_reg_494;
        tmp_reg_494_pp0_iter2_reg <= tmp_reg_494_pp0_iter1_reg;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (tmp_fu_323_p3 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        trunc_ln25_reg_498 <= trunc_ln25_fu_336_p1;
    end
end

always @ (*) begin
    if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
        if (((1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            accum_in_0_address0 = zext_ln29_24_fu_412_p1;
        end else if (((1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            accum_in_0_address0 = zext_ln29_22_fu_386_p1;
        end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            accum_in_0_address0 = zext_ln29_20_fu_366_p1;
        end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            accum_in_0_address0 = zext_ln29_fu_346_p1;
        end else begin
            accum_in_0_address0 = 'bx;
        end
    end else begin
        accum_in_0_address0 = 'bx;
    end
end

always @ (*) begin
    if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
        if (((1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            accum_in_0_address1 = zext_ln29_23_fu_402_p1;
        end else if (((1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            accum_in_0_address1 = zext_ln29_21_fu_376_p1;
        end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            accum_in_0_address1 = zext_ln29_19_fu_356_p1;
        end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            accum_in_0_address1 = zext_ln25_fu_331_p1;
        end else begin
            accum_in_0_address1 = 'bx;
        end
    end else begin
        accum_in_0_address1 = 'bx;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1)) | ((1'b0 == ap_block_pp0_stage3_11001) & (1'b1 == ap_CS_fsm_pp0_stage3) & (ap_enable_reg_pp0_iter0 == 1'b1)) | ((1'b0 == ap_block_pp0_stage2_11001) & (1'b1 == ap_CS_fsm_pp0_stage2) & (ap_enable_reg_pp0_iter0 == 1'b1)) | ((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1)))) begin
        accum_in_0_ce0 = 1'b1;
    end else begin
        accum_in_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1)) | ((1'b0 == ap_block_pp0_stage3_11001) & (1'b1 == ap_CS_fsm_pp0_stage3) & (ap_enable_reg_pp0_iter0 == 1'b1)) | ((1'b0 == ap_block_pp0_stage2_11001) & (1'b1 == ap_CS_fsm_pp0_stage2) & (ap_enable_reg_pp0_iter0 == 1'b1)) | ((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1)))) begin
        accum_in_0_ce1 = 1'b1;
    end else begin
        accum_in_0_ce1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state13)) begin
        accum_out_ce0 = 1'b1;
    end else begin
        accum_out_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state13)) begin
        accum_out_ce1 = 1'b1;
    end else begin
        accum_out_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((tmp_48_fu_417_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state13))) begin
        accum_out_we0 = 1'b1;
    end else begin
        accum_out_we0 = 1'b0;
    end
end

always @ (*) begin
    if (((tmp_48_fu_417_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state13))) begin
        accum_out_we1 = 1'b1;
    end else begin
        accum_out_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((tmp_reg_494 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state4 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state4 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state14)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((tmp_48_fu_417_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state13))) begin
        if ((trunc_ln33_fu_430_p1 == 3'd0)) begin
            ap_phi_mux_phi_ln45_phi_fu_292_p8 = psum_0_01_reg_266;
        end else if ((1'b1 == ap_condition_517)) begin
            ap_phi_mux_phi_ln45_phi_fu_292_p8 = psum_6_07_reg_194;
        end else if ((trunc_ln33_fu_430_p1 == 3'd4)) begin
            ap_phi_mux_phi_ln45_phi_fu_292_p8 = psum_4_05_reg_218;
        end else if ((trunc_ln33_fu_430_p1 == 3'd2)) begin
            ap_phi_mux_phi_ln45_phi_fu_292_p8 = psum_2_03_reg_242;
        end else begin
            ap_phi_mux_phi_ln45_phi_fu_292_p8 = 'bx;
        end
    end else begin
        ap_phi_mux_phi_ln45_phi_fu_292_p8 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0) & (tmp_reg_494 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_x_phi_fu_174_p4 = add_ln25_reg_558;
    end else begin
        ap_phi_mux_x_phi_fu_174_p4 = x_reg_170;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state14)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_307_p0 = ap_phi_mux_psum_6_07_phi_fu_198_p4;
    end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_307_p0 = ap_phi_mux_psum_4_05_phi_fu_222_p4;
    end else if (((1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
        grp_fu_307_p0 = ap_phi_mux_psum_2_03_phi_fu_246_p4;
    end else if (((1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
        grp_fu_307_p0 = grp_fu_307_p2;
    end else begin
        grp_fu_307_p0 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_307_p1 = accum_in_0_load_63_reg_583;
    end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_307_p1 = accum_in_0_load_61_reg_563;
    end else if (((1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
        grp_fu_307_p1 = accum_in_0_load_59_reg_538;
    end else if (((1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
        grp_fu_307_p1 = accum_in_0_load_reg_518;
    end else begin
        grp_fu_307_p1 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_312_p0 = ap_phi_mux_psum_7_08_phi_fu_186_p4;
    end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_312_p0 = ap_phi_mux_psum_5_06_phi_fu_210_p4;
    end else if (((1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
        grp_fu_312_p0 = ap_phi_mux_psum_3_04_phi_fu_234_p4;
    end else if (((1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
        grp_fu_312_p0 = grp_fu_312_p2;
    end else begin
        grp_fu_312_p0 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_312_p1 = accum_in_0_load_64_reg_588;
    end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_312_p1 = accum_in_0_load_62_reg_568;
    end else if (((1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
        grp_fu_312_p1 = accum_in_0_load_60_reg_543;
    end else if (((1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
        grp_fu_312_p1 = accum_in_0_load_58_reg_523;
    end else begin
        grp_fu_312_p1 = 'bx;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_pp0_stage1 : begin
            if ((~((1'b0 == ap_block_pp0_stage1_subdone) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b0)) & (1'b0 == ap_block_pp0_stage1_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage2;
            end else if (((1'b0 == ap_block_pp0_stage1_subdone) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
                ap_NS_fsm = ap_ST_fsm_state12;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end
        end
        ap_ST_fsm_pp0_stage2 : begin
            if ((~((1'b0 == ap_block_pp0_stage2_subdone) & (tmp_reg_494 == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1)) & (1'b0 == ap_block_pp0_stage2_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage3;
            end else if (((1'b0 == ap_block_pp0_stage2_subdone) & (tmp_reg_494 == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
                ap_NS_fsm = ap_ST_fsm_state12;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage2;
            end
        end
        ap_ST_fsm_pp0_stage3 : begin
            if ((1'b0 == ap_block_pp0_stage3_subdone)) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage3;
            end
        end
        ap_ST_fsm_state12 : begin
            ap_NS_fsm = ap_ST_fsm_state13;
        end
        ap_ST_fsm_state13 : begin
            if (((tmp_48_fu_417_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state13))) begin
                ap_NS_fsm = ap_ST_fsm_state13;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state14;
            end
        end
        ap_ST_fsm_state14 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign accum_out_address0 = zext_ln33_4_fu_446_p1;

assign accum_out_address1 = zext_ln33_fu_425_p1;

assign accum_out_d0 = ((icmp_ln45_8_fu_479_p2[0:0] == 1'b1) ? psum_5_06_reg_206 : select_ln45_7_fu_471_p3);

assign accum_out_d1 = ap_phi_mux_phi_ln45_phi_fu_292_p8;

assign add_ln25_fu_391_p2 = (x_reg_170 + 8'd8);

assign add_ln33_fu_434_p2 = (q_reg_278 + 4'd2);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_pp0_stage1 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_pp0_stage2 = ap_CS_fsm[32'd3];

assign ap_CS_fsm_pp0_stage3 = ap_CS_fsm[32'd4];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state12 = ap_CS_fsm[32'd5];

assign ap_CS_fsm_state13 = ap_CS_fsm[32'd6];

assign ap_CS_fsm_state14 = ap_CS_fsm[32'd7];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1_subdone = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage2 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage2_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage2_subdone = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage3 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage3_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage3_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((ap_done_reg == 1'b1) | (ap_start == 1'b0));
end

assign ap_block_state10_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state11_pp0_stage1_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage1_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage2_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage3_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage1_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage2_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state9_pp0_stage3_iter1 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_condition_517 = (~(trunc_ln33_fu_430_p1 == 3'd0) & ~(trunc_ln33_fu_430_p1 == 3'd4) & ~(trunc_ln33_fu_430_p1 == 3'd2));
end

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign ap_phi_mux_psum_2_03_phi_fu_246_p4 = grp_fu_307_p2;

assign ap_phi_mux_psum_3_04_phi_fu_234_p4 = grp_fu_312_p2;

assign ap_phi_mux_psum_4_05_phi_fu_222_p4 = grp_fu_307_p2;

assign ap_phi_mux_psum_5_06_phi_fu_210_p4 = grp_fu_312_p2;

assign ap_phi_mux_psum_6_07_phi_fu_198_p4 = grp_fu_307_p2;

assign ap_phi_mux_psum_7_08_phi_fu_186_p4 = grp_fu_312_p2;

assign icmp_ln45_7_fu_465_p2 = ((or_ln33_fu_440_p2 == 3'd3) ? 1'b1 : 1'b0);

assign icmp_ln45_8_fu_479_p2 = ((or_ln33_fu_440_p2 == 3'd5) ? 1'b1 : 1'b0);

assign icmp_ln45_fu_451_p2 = ((or_ln33_fu_440_p2 == 3'd1) ? 1'b1 : 1'b0);

assign or_ln29_19_fu_351_p2 = (trunc_ln25_reg_498 | 7'd2);

assign or_ln29_20_fu_361_p2 = (trunc_ln25_reg_498 | 7'd3);

assign or_ln29_21_fu_371_p2 = (trunc_ln25_reg_498 | 7'd4);

assign or_ln29_22_fu_381_p2 = (trunc_ln25_reg_498 | 7'd5);

assign or_ln29_23_fu_397_p2 = (trunc_ln25_reg_498 | 7'd6);

assign or_ln29_24_fu_407_p2 = (trunc_ln25_reg_498 | 7'd7);

assign or_ln29_fu_340_p2 = (trunc_ln25_fu_336_p1 | 7'd1);

assign or_ln33_fu_440_p2 = (trunc_ln33_fu_430_p1 | 3'd1);

assign select_ln45_7_fu_471_p3 = ((icmp_ln45_7_fu_465_p2[0:0] == 1'b1) ? psum_3_04_reg_230 : select_ln45_fu_457_p3);

assign select_ln45_fu_457_p3 = ((icmp_ln45_fu_451_p2[0:0] == 1'b1) ? psum_1_02_reg_254 : psum_7_08_reg_182);

assign tmp_48_fu_417_p3 = q_reg_278[32'd3];

assign tmp_fu_323_p3 = ap_phi_mux_x_phi_fu_174_p4[32'd7];

assign trunc_ln25_fu_336_p1 = ap_phi_mux_x_phi_fu_174_p4[6:0];

assign trunc_ln33_fu_430_p1 = q_reg_278[2:0];

assign zext_ln25_fu_331_p1 = ap_phi_mux_x_phi_fu_174_p4;

assign zext_ln29_19_fu_356_p1 = or_ln29_19_fu_351_p2;

assign zext_ln29_20_fu_366_p1 = or_ln29_20_fu_361_p2;

assign zext_ln29_21_fu_376_p1 = or_ln29_21_fu_371_p2;

assign zext_ln29_22_fu_386_p1 = or_ln29_22_fu_381_p2;

assign zext_ln29_23_fu_402_p1 = or_ln29_23_fu_397_p2;

assign zext_ln29_24_fu_412_p1 = or_ln29_24_fu_407_p2;

assign zext_ln29_fu_346_p1 = or_ln29_fu_340_p2;

assign zext_ln33_4_fu_446_p1 = or_ln33_fu_440_p2;

assign zext_ln33_fu_425_p1 = q_reg_278;

endmodule //td_fused_top_tdf12_accum_1
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf12_accum_2 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        accum_in_20,
        accum_in_20_ap_vld,
        accum_in_address0,
        accum_in_ce0,
        accum_in_q0
);

parameter    ap_ST_fsm_state1 = 7'd1;
parameter    ap_ST_fsm_state2 = 7'd2;
parameter    ap_ST_fsm_state3 = 7'd4;
parameter    ap_ST_fsm_state4 = 7'd8;
parameter    ap_ST_fsm_state5 = 7'd16;
parameter    ap_ST_fsm_state6 = 7'd32;
parameter    ap_ST_fsm_state7 = 7'd64;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [15:0] accum_in_20;
output   accum_in_20_ap_vld;
output  [2:0] accum_in_address0;
output   accum_in_ce0;
input  [15:0] accum_in_q0;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg[15:0] accum_in_20;
reg accum_in_20_ap_vld;
reg accum_in_ce0;

reg    ap_done_reg;
  reg   [6:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
wire   [3:0] add_ln57_fu_74_p2;
reg   [3:0] add_ln57_reg_91;
wire    ap_CS_fsm_state2;
wire   [0:0] icmp_ln57_fu_85_p2;
wire    ap_CS_fsm_state3;
wire   [15:0] grp_fu_68_p2;
wire    ap_CS_fsm_state7;
reg   [3:0] i_1_1_reg_44;
reg    ap_block_state1;
reg   [15:0] sum_01_reg_55;
wire   [63:0] zext_ln57_fu_80_p1;
reg   [15:0] accum_in_20_preg;
reg   [6:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 7'd1;
#0 accum_in_20_preg = 16'd0;
end

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U779(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(sum_01_reg_55),
    .din1(accum_in_q0),
    .dout(grp_fu_68_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        accum_in_20_preg <= 16'd0;
    end else begin
        if (((icmp_ln57_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
            accum_in_20_preg <= sum_01_reg_55;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if (((icmp_ln57_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        i_1_1_reg_44 <= 4'd0;
    end else if ((1'b1 == ap_CS_fsm_state7)) begin
        i_1_1_reg_44 <= add_ln57_reg_91;
    end
end

always @ (posedge ap_clk) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        sum_01_reg_55 <= 16'd0;
    end else if ((1'b1 == ap_CS_fsm_state7)) begin
        sum_01_reg_55 <= grp_fu_68_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        add_ln57_reg_91 <= add_ln57_fu_74_p2;
    end
end

always @ (*) begin
    if (((icmp_ln57_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        accum_in_20 = sum_01_reg_55;
    end else begin
        accum_in_20 = accum_in_20_preg;
    end
end

always @ (*) begin
    if (((icmp_ln57_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        accum_in_20_ap_vld = 1'b1;
    end else begin
        accum_in_20_ap_vld = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        accum_in_ce0 = 1'b1;
    end else begin
        accum_in_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln57_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln57_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_state2 : begin
            if (((icmp_ln57_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end
        end
        ap_ST_fsm_state3 : begin
            ap_NS_fsm = ap_ST_fsm_state4;
        end
        ap_ST_fsm_state4 : begin
            ap_NS_fsm = ap_ST_fsm_state5;
        end
        ap_ST_fsm_state5 : begin
            ap_NS_fsm = ap_ST_fsm_state6;
        end
        ap_ST_fsm_state6 : begin
            ap_NS_fsm = ap_ST_fsm_state7;
        end
        ap_ST_fsm_state7 : begin
            ap_NS_fsm = ap_ST_fsm_state2;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign accum_in_address0 = zext_ln57_fu_80_p1;

assign add_ln57_fu_74_p2 = (i_1_1_reg_44 + 4'd1);

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state7 = ap_CS_fsm[32'd6];

always @ (*) begin
    ap_block_state1 = ((ap_done_reg == 1'b1) | (ap_start == 1'b0));
end

assign icmp_ln57_fu_85_p2 = ((i_1_1_reg_44 == 4'd8) ? 1'b1 : 1'b0);

assign zext_ln57_fu_80_p1 = i_1_1_reg_44;

endmodule //td_fused_top_tdf12_accum_2
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_tdf12_adjustments_ram (addr0, ce0, q0, addr1, ce1, d1, we1,  clk);

parameter DWIDTH = 48;
parameter AWIDTH = 10;
parameter MEM_SIZE = 1000;

input[AWIDTH-1:0] addr0;
input ce0;
output wire[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
input clk;

 reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];
wire [AWIDTH-1:0] addr0_t0; 
reg [AWIDTH-1:0] addr0_t1; 
reg [DWIDTH-1:0] q0_t0;
reg [DWIDTH-1:0] q0_t1;
wire [AWIDTH-1:0] addr1_t0; 
reg [AWIDTH-1:0] addr1_t1; 
wire [DWIDTH-1:0] d1_t0; 
wire we1_t0; 
reg [DWIDTH-1:0] d1_t1; 
reg we1_t1; 


assign addr0_t0 = addr0;
assign q0 = q0_t1;
assign addr1_t0 = addr1;
assign d1_t0 = d1;
assign we1_t0 = we1;

always @(posedge clk)  
begin
    if (ce0) 
    begin
        addr0_t1 <= addr0_t0; 
        q0_t1 <= q0_t0;
    end
    if (ce1) 
    begin
        addr1_t1 <= addr1_t0; 
        d1_t1 <= d1_t0;
        we1_t1 <= we1_t0;
    end
end


always @(posedge clk)  
begin 
    if (ce0) begin
        q0_t0 <= ram[addr0_t1];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1_t1) 
            ram[addr1_t1] <= d1_t1; 
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_tdf12_adjustments(
    reset,
    clk,
    address0,
    ce0,
    q0,
    address1,
    ce1,
    we1,
    d1);

parameter DataWidth = 32'd48;
parameter AddressRange = 32'd1000;
parameter AddressWidth = 32'd10;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;



td_fused_top_tdf12_adjustments_ram td_fused_top_tdf12_adjustments_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 )
);

endmodule

// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf12_adjust (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        sums_read,
        adjustments_address0,
        adjustments_ce0,
        adjustments_q0,
        indices_23_dout,
        indices_23_empty_n,
        indices_23_read,
        ap_return
);

parameter    ap_ST_fsm_state1 = 17'd1;
parameter    ap_ST_fsm_state2 = 17'd2;
parameter    ap_ST_fsm_state3 = 17'd4;
parameter    ap_ST_fsm_state4 = 17'd8;
parameter    ap_ST_fsm_state5 = 17'd16;
parameter    ap_ST_fsm_state6 = 17'd32;
parameter    ap_ST_fsm_state7 = 17'd64;
parameter    ap_ST_fsm_state8 = 17'd128;
parameter    ap_ST_fsm_state9 = 17'd256;
parameter    ap_ST_fsm_state10 = 17'd512;
parameter    ap_ST_fsm_state11 = 17'd1024;
parameter    ap_ST_fsm_state12 = 17'd2048;
parameter    ap_ST_fsm_state13 = 17'd4096;
parameter    ap_ST_fsm_state14 = 17'd8192;
parameter    ap_ST_fsm_state15 = 17'd16384;
parameter    ap_ST_fsm_state16 = 17'd32768;
parameter    ap_ST_fsm_state17 = 17'd65536;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
input  [15:0] sums_read;
output  [9:0] adjustments_address0;
output   adjustments_ce0;
input  [47:0] adjustments_q0;
input  [9:0] indices_23_dout;
input   indices_23_empty_n;
output   indices_23_read;
output  [15:0] ap_return;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg adjustments_ce0;
reg indices_23_read;

reg    ap_done_reg;
  reg   [16:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    indices_23_blk_n;
wire    ap_CS_fsm_state4;
reg   [15:0] tmp_82_i_i_reg_167;
reg   [15:0] tmp_83_i_i_reg_172;
wire   [15:0] grp_fu_81_p2;
reg   [15:0] sub_i_i_i_reg_177;
wire    ap_CS_fsm_state8;
wire    ap_CS_fsm_state9;
wire   [15:0] grp_fu_86_p2;
reg   [15:0] mul_i_i_i_reg_187;
wire    ap_CS_fsm_state12;
wire    ap_CS_fsm_state13;
wire   [63:0] zext_ln220_fu_90_p1;
reg    ap_block_state1;
wire    ap_CS_fsm_state2;
wire    ap_CS_fsm_state3;
wire   [15:0] grp_fu_77_p1;
wire   [15:0] grp_fu_81_p1;
wire   [15:0] grp_fu_86_p1;
wire   [15:0] trunc_ln220_fu_95_p1;
wire   [15:0] grp_fu_77_p2;
wire    ap_CS_fsm_state17;
wire   [15:0] bitcast_ln648_fu_132_p1;
wire   [0:0] tmp_fu_136_p3;
reg   [16:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 17'd1;
end

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U783(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(mul_i_i_i_reg_187),
    .din1(grp_fu_77_p1),
    .dout(grp_fu_77_p2)
);

td_fused_top_hsub_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hsub_16ns_16ns_16_5_full_dsp_1_U784(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(sums_read),
    .din1(grp_fu_81_p1),
    .dout(grp_fu_81_p2)
);

td_fused_top_hmul_16ns_16ns_16_4_max_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hmul_16ns_16ns_16_4_max_dsp_1_U785(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(sub_i_i_i_reg_177),
    .din1(grp_fu_86_p1),
    .dout(grp_fu_86_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state17)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state12)) begin
        mul_i_i_i_reg_187 <= grp_fu_86_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state8)) begin
        sub_i_i_i_reg_177 <= grp_fu_81_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        tmp_82_i_i_reg_167 <= {{adjustments_q0[31:16]}};
        tmp_83_i_i_reg_172 <= {{adjustments_q0[47:32]}};
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state2) | (~((indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1)))) begin
        adjustments_ce0 = 1'b1;
    end else begin
        adjustments_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state17)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state17)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_23_blk_n = indices_23_empty_n;
    end else begin
        indices_23_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_23_read = 1'b1;
    end else begin
        indices_23_read = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_state2 : begin
            ap_NS_fsm = ap_ST_fsm_state3;
        end
        ap_ST_fsm_state3 : begin
            ap_NS_fsm = ap_ST_fsm_state4;
        end
        ap_ST_fsm_state4 : begin
            ap_NS_fsm = ap_ST_fsm_state5;
        end
        ap_ST_fsm_state5 : begin
            ap_NS_fsm = ap_ST_fsm_state6;
        end
        ap_ST_fsm_state6 : begin
            ap_NS_fsm = ap_ST_fsm_state7;
        end
        ap_ST_fsm_state7 : begin
            ap_NS_fsm = ap_ST_fsm_state8;
        end
        ap_ST_fsm_state8 : begin
            ap_NS_fsm = ap_ST_fsm_state9;
        end
        ap_ST_fsm_state9 : begin
            ap_NS_fsm = ap_ST_fsm_state10;
        end
        ap_ST_fsm_state10 : begin
            ap_NS_fsm = ap_ST_fsm_state11;
        end
        ap_ST_fsm_state11 : begin
            ap_NS_fsm = ap_ST_fsm_state12;
        end
        ap_ST_fsm_state12 : begin
            ap_NS_fsm = ap_ST_fsm_state13;
        end
        ap_ST_fsm_state13 : begin
            ap_NS_fsm = ap_ST_fsm_state14;
        end
        ap_ST_fsm_state14 : begin
            ap_NS_fsm = ap_ST_fsm_state15;
        end
        ap_ST_fsm_state15 : begin
            ap_NS_fsm = ap_ST_fsm_state16;
        end
        ap_ST_fsm_state16 : begin
            ap_NS_fsm = ap_ST_fsm_state17;
        end
        ap_ST_fsm_state17 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign adjustments_address0 = zext_ln220_fu_90_p1;

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state12 = ap_CS_fsm[32'd11];

assign ap_CS_fsm_state13 = ap_CS_fsm[32'd12];

assign ap_CS_fsm_state17 = ap_CS_fsm[32'd16];

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

assign ap_CS_fsm_state8 = ap_CS_fsm[32'd7];

assign ap_CS_fsm_state9 = ap_CS_fsm[32'd8];

always @ (*) begin
    ap_block_state1 = ((indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0));
end

assign ap_return = ((tmp_fu_136_p3[0:0] == 1'b1) ? 16'd0 : grp_fu_77_p2);

assign bitcast_ln648_fu_132_p1 = grp_fu_77_p2;

assign grp_fu_77_p1 = tmp_83_i_i_reg_172;

assign grp_fu_81_p1 = trunc_ln220_fu_95_p1;

assign grp_fu_86_p1 = tmp_82_i_i_reg_167;

assign tmp_fu_136_p3 = bitcast_ln648_fu_132_p1[32'd15];

assign trunc_ln220_fu_95_p1 = adjustments_q0[15:0];

assign zext_ln220_fu_90_p1 = indices_23_dout;

endmodule //td_fused_top_tdf12_adjust
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf12_dot_product (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        ifmap_vec_0_0_address0,
        ifmap_vec_0_0_ce0,
        ifmap_vec_0_0_q0,
        weight_vecs_0_0_0_address0,
        weight_vecs_0_0_0_ce0,
        weight_vecs_0_0_0_q0,
        products_0_address0,
        products_0_ce0,
        products_0_we0,
        products_0_d0
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state9 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [6:0] ifmap_vec_0_0_address0;
output   ifmap_vec_0_0_ce0;
input  [15:0] ifmap_vec_0_0_q0;
output  [6:0] weight_vecs_0_0_0_address0;
output   weight_vecs_0_0_0_ce0;
input  [15:0] weight_vecs_0_0_0_q0;
output  [6:0] products_0_address0;
output   products_0_ce0;
output   products_0_we0;
output  [15:0] products_0_d0;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg ifmap_vec_0_0_ce0;
reg weight_vecs_0_0_0_ce0;
reg products_0_ce0;
reg products_0_we0;

reg    ap_done_reg;
  reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg   [7:0] ic_0_0_reg_69;
wire   [7:0] add_ln149_fu_84_p2;
wire    ap_CS_fsm_pp0_stage0;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
wire    ap_block_state4_pp0_stage0_iter2;
wire    ap_block_state5_pp0_stage0_iter3;
wire    ap_block_state6_pp0_stage0_iter4;
wire    ap_block_state7_pp0_stage0_iter5;
wire    ap_block_state8_pp0_stage0_iter6;
wire    ap_block_pp0_stage0_11001;
wire   [0:0] icmp_ln149_fu_90_p2;
reg   [0:0] icmp_ln149_reg_107;
reg   [0:0] icmp_ln149_reg_107_pp0_iter1_reg;
reg   [0:0] icmp_ln149_reg_107_pp0_iter2_reg;
reg   [0:0] icmp_ln149_reg_107_pp0_iter3_reg;
reg   [0:0] icmp_ln149_reg_107_pp0_iter4_reg;
reg   [0:0] icmp_ln149_reg_107_pp0_iter5_reg;
wire   [63:0] idxprom17_0_0_fu_96_p1;
reg   [63:0] idxprom17_0_0_reg_111;
reg   [63:0] idxprom17_0_0_reg_111_pp0_iter1_reg;
reg   [63:0] idxprom17_0_0_reg_111_pp0_iter2_reg;
reg   [63:0] idxprom17_0_0_reg_111_pp0_iter3_reg;
reg   [63:0] idxprom17_0_0_reg_111_pp0_iter4_reg;
reg   [63:0] idxprom17_0_0_reg_111_pp0_iter5_reg;
reg   [15:0] ifmap_vec_0_0_load_reg_126;
reg   [15:0] weight_vecs_0_0_0_load_reg_131;
wire   [15:0] grp_fu_80_p2;
reg   [15:0] mul_reg_136;
reg    ap_block_state1;
wire    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_exit_iter0_state2;
reg    ap_enable_reg_pp0_iter1;
reg    ap_enable_reg_pp0_iter2;
reg    ap_enable_reg_pp0_iter3;
reg    ap_enable_reg_pp0_iter4;
reg    ap_enable_reg_pp0_iter5;
reg    ap_enable_reg_pp0_iter6;
wire    ap_block_pp0_stage0;
wire    ap_CS_fsm_state9;
reg   [2:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
#0 ap_enable_reg_pp0_iter4 = 1'b0;
#0 ap_enable_reg_pp0_iter5 = 1'b0;
#0 ap_enable_reg_pp0_iter6 = 1'b0;
end

td_fused_top_hmul_16ns_16ns_16_4_max_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hmul_16ns_16ns_16_4_max_dsp_1_U771(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(ifmap_vec_0_0_load_reg_126),
    .din1(weight_vecs_0_0_0_load_reg_131),
    .dout(grp_fu_80_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b1 == ap_condition_pp0_exit_iter0_state2))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            if ((1'b1 == ap_condition_pp0_exit_iter0_state2)) begin
                ap_enable_reg_pp0_iter1 <= (1'b1 ^ ap_condition_pp0_exit_iter0_state2);
            end else if ((1'b1 == 1'b1)) begin
                ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
            end
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter4 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter5 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter5 <= ap_enable_reg_pp0_iter4;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter6 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter6 <= ap_enable_reg_pp0_iter5;
        end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter6 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln149_fu_90_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ic_0_0_reg_69 <= add_ln149_fu_84_p2;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ic_0_0_reg_69 <= 8'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln149_reg_107 <= icmp_ln149_fu_90_p2;
        icmp_ln149_reg_107_pp0_iter1_reg <= icmp_ln149_reg_107;
        idxprom17_0_0_reg_111_pp0_iter1_reg[7 : 0] <= idxprom17_0_0_reg_111[7 : 0];
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        icmp_ln149_reg_107_pp0_iter2_reg <= icmp_ln149_reg_107_pp0_iter1_reg;
        icmp_ln149_reg_107_pp0_iter3_reg <= icmp_ln149_reg_107_pp0_iter2_reg;
        icmp_ln149_reg_107_pp0_iter4_reg <= icmp_ln149_reg_107_pp0_iter3_reg;
        icmp_ln149_reg_107_pp0_iter5_reg <= icmp_ln149_reg_107_pp0_iter4_reg;
        idxprom17_0_0_reg_111_pp0_iter2_reg[7 : 0] <= idxprom17_0_0_reg_111_pp0_iter1_reg[7 : 0];
        idxprom17_0_0_reg_111_pp0_iter3_reg[7 : 0] <= idxprom17_0_0_reg_111_pp0_iter2_reg[7 : 0];
        idxprom17_0_0_reg_111_pp0_iter4_reg[7 : 0] <= idxprom17_0_0_reg_111_pp0_iter3_reg[7 : 0];
        idxprom17_0_0_reg_111_pp0_iter5_reg[7 : 0] <= idxprom17_0_0_reg_111_pp0_iter4_reg[7 : 0];
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln149_fu_90_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        idxprom17_0_0_reg_111[7 : 0] <= idxprom17_0_0_fu_96_p1[7 : 0];
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln149_reg_107 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ifmap_vec_0_0_load_reg_126 <= ifmap_vec_0_0_q0;
        weight_vecs_0_0_0_load_reg_131 <= weight_vecs_0_0_0_q0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln149_reg_107_pp0_iter4_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        mul_reg_136 <= grp_fu_80_p2;
    end
end

always @ (*) begin
    if ((icmp_ln149_fu_90_p2 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state2 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state2 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state9)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state9)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ifmap_vec_0_0_ce0 = 1'b1;
    end else begin
        ifmap_vec_0_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter6 == 1'b1))) begin
        products_0_ce0 = 1'b1;
    end else begin
        products_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln149_reg_107_pp0_iter5_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter6 == 1'b1))) begin
        products_0_we0 = 1'b1;
    end else begin
        products_0_we0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        weight_vecs_0_0_0_ce0 = 1'b1;
    end else begin
        weight_vecs_0_0_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((~((icmp_ln149_fu_90_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0)) & ~((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter6 == 1'b1) & (ap_enable_reg_pp0_iter5 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if ((((icmp_ln149_fu_90_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0)) | ((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter6 == 1'b1) & (ap_enable_reg_pp0_iter5 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_state9;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state9 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln149_fu_84_p2 = (ic_0_0_reg_69 + 8'd1);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state9 = ap_CS_fsm[32'd2];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (ap_done_reg == 1'b1));
end

assign ap_block_state2_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter4 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage0_iter5 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage0_iter6 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign icmp_ln149_fu_90_p2 = ((ic_0_0_reg_69 == 8'd128) ? 1'b1 : 1'b0);

assign idxprom17_0_0_fu_96_p1 = ic_0_0_reg_69;

assign ifmap_vec_0_0_address0 = idxprom17_0_0_fu_96_p1;

assign products_0_address0 = idxprom17_0_0_reg_111_pp0_iter5_reg;

assign products_0_d0 = mul_reg_136;

assign weight_vecs_0_0_0_address0 = idxprom17_0_0_fu_96_p1;

always @ (posedge ap_clk) begin
    idxprom17_0_0_reg_111[63:8] <= 56'b00000000000000000000000000000000000000000000000000000000;
    idxprom17_0_0_reg_111_pp0_iter1_reg[63:8] <= 56'b00000000000000000000000000000000000000000000000000000000;
    idxprom17_0_0_reg_111_pp0_iter2_reg[63:8] <= 56'b00000000000000000000000000000000000000000000000000000000;
    idxprom17_0_0_reg_111_pp0_iter3_reg[63:8] <= 56'b00000000000000000000000000000000000000000000000000000000;
    idxprom17_0_0_reg_111_pp0_iter4_reg[63:8] <= 56'b00000000000000000000000000000000000000000000000000000000;
    idxprom17_0_0_reg_111_pp0_iter5_reg[63:8] <= 56'b00000000000000000000000000000000000000000000000000000000;
end

endmodule //td_fused_top_tdf12_dot_product
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_tdf12_filters_ram (addr0, ce0, q0, addr1, ce1, d1, we1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 17;
parameter MEM_SIZE = 128000;

input[AWIDTH-1:0] addr0;
input ce0;
output wire[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
input clk;

 reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];
wire [AWIDTH-1:0] addr0_t0; 
reg [AWIDTH-1:0] addr0_t1; 
reg [DWIDTH-1:0] q0_t0;
reg [DWIDTH-1:0] q0_t1;
wire [AWIDTH-1:0] addr1_t0; 
reg [AWIDTH-1:0] addr1_t1; 
wire [DWIDTH-1:0] d1_t0; 
wire we1_t0; 
reg [DWIDTH-1:0] d1_t1; 
reg we1_t1; 


assign addr0_t0 = addr0;
assign q0 = q0_t1;
assign addr1_t0 = addr1;
assign d1_t0 = d1;
assign we1_t0 = we1;

always @(posedge clk)  
begin
    if (ce0) 
    begin
        addr0_t1 <= addr0_t0; 
        q0_t1 <= q0_t0;
    end
    if (ce1) 
    begin
        addr1_t1 <= addr1_t0; 
        d1_t1 <= d1_t0;
        we1_t1 <= we1_t0;
    end
end


always @(posedge clk)  
begin 
    if (ce0) begin
        q0_t0 <= ram[addr0_t1];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1_t1) 
            ram[addr1_t1] <= d1_t1; 
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_tdf12_filters(
    reset,
    clk,
    address0,
    ce0,
    q0,
    address1,
    ce1,
    we1,
    d1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd128000;
parameter AddressWidth = 32'd17;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;



td_fused_top_tdf12_filters_ram td_fused_top_tdf12_filters_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 )
);

endmodule

// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf12_get_next_ijk (
        ap_clk,
        ap_rst,
        ap_start,
        start_full_n,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        start_out,
        start_write,
        indices_0_din,
        indices_0_full_n,
        indices_0_write,
        indices_1_din,
        indices_1_full_n,
        indices_1_write,
        indices_2_out_din,
        indices_2_out_full_n,
        indices_2_out_write,
        indices_2_out1_din,
        indices_2_out1_full_n,
        indices_2_out1_write
);

parameter    ap_ST_fsm_state1 = 1'd1;

input   ap_clk;
input   ap_rst;
input   ap_start;
input   start_full_n;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output   start_out;
output   start_write;
output  [15:0] indices_0_din;
input   indices_0_full_n;
output   indices_0_write;
output  [15:0] indices_1_din;
input   indices_1_full_n;
output   indices_1_write;
output  [9:0] indices_2_out_din;
input   indices_2_out_full_n;
output   indices_2_out_write;
output  [9:0] indices_2_out1_din;
input   indices_2_out1_full_n;
output   indices_2_out1_write;

reg ap_done;
reg ap_idle;
reg start_write;
reg indices_0_write;
reg indices_1_write;
reg indices_2_out_write;
reg indices_2_out1_write;

reg    real_start;
reg    start_once_reg;
reg    ap_done_reg;
  reg   [0:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    internal_ap_ready;
reg   [15:0] i_5;
reg   [15:0] j_5;
reg   [15:0] k_5;
reg    indices_0_blk_n;
reg    indices_1_blk_n;
reg    indices_2_out_blk_n;
reg    indices_2_out1_blk_n;
reg   [0:0] ap_phi_mux_j_9_flag_0_i_phi_fu_77_p6;
reg    ap_block_state1;
wire   [0:0] icmp_ln78_fu_141_p2;
wire   [0:0] icmp_ln81_fu_154_p2;
reg   [15:0] ap_phi_mux_j_9_new_0_i_phi_fu_91_p6;
wire   [15:0] add_ln80_fu_147_p2;
reg   [15:0] ap_phi_mux_k_9_new_0_i_phi_fu_104_p6;
wire   [15:0] add_ln77_fu_134_p2;
wire   [15:0] select_ln84_fu_172_p3;
wire   [9:0] trunc_ln76_fu_128_p1;
wire   [15:0] add_ln83_fu_160_p2;
wire   [0:0] icmp_ln84_fu_166_p2;
reg   [0:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 start_once_reg = 1'b0;
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 1'd1;
#0 i_5 = 16'd0;
#0 j_5 = 16'd0;
#0 k_5 = 16'd0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((~((real_start == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        start_once_reg <= 1'b0;
    end else begin
        if (((real_start == 1'b1) & (internal_ap_ready == 1'b0))) begin
            start_once_reg <= 1'b1;
        end else if ((internal_ap_ready == 1'b1)) begin
            start_once_reg <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((~((real_start == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (icmp_ln81_fu_154_p2 == 1'd1) & (icmp_ln78_fu_141_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1))) begin
        i_5 <= select_ln84_fu_172_p3;
    end
end

always @ (posedge ap_clk) begin
    if ((~((real_start == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (ap_phi_mux_j_9_flag_0_i_phi_fu_77_p6 == 1'd1) & (1'b1 == ap_CS_fsm_state1))) begin
        j_5 <= ap_phi_mux_j_9_new_0_i_phi_fu_91_p6;
    end
end

always @ (posedge ap_clk) begin
    if ((~((real_start == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        k_5 <= ap_phi_mux_k_9_new_0_i_phi_fu_104_p6;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((real_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln78_fu_141_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_phi_mux_j_9_flag_0_i_phi_fu_77_p6 = 1'd0;
    end else if ((((icmp_ln81_fu_154_p2 == 1'd0) & (icmp_ln78_fu_141_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1)) | ((icmp_ln81_fu_154_p2 == 1'd1) & (icmp_ln78_fu_141_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1)))) begin
        ap_phi_mux_j_9_flag_0_i_phi_fu_77_p6 = 1'd1;
    end else begin
        ap_phi_mux_j_9_flag_0_i_phi_fu_77_p6 = 'bx;
    end
end

always @ (*) begin
    if (((icmp_ln78_fu_141_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1))) begin
        if ((icmp_ln81_fu_154_p2 == 1'd0)) begin
            ap_phi_mux_j_9_new_0_i_phi_fu_91_p6 = add_ln80_fu_147_p2;
        end else if ((icmp_ln81_fu_154_p2 == 1'd1)) begin
            ap_phi_mux_j_9_new_0_i_phi_fu_91_p6 = 16'd0;
        end else begin
            ap_phi_mux_j_9_new_0_i_phi_fu_91_p6 = 'bx;
        end
    end else begin
        ap_phi_mux_j_9_new_0_i_phi_fu_91_p6 = 'bx;
    end
end

always @ (*) begin
    if (((icmp_ln78_fu_141_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_phi_mux_k_9_new_0_i_phi_fu_104_p6 = add_ln77_fu_134_p2;
    end else if ((((icmp_ln81_fu_154_p2 == 1'd0) & (icmp_ln78_fu_141_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1)) | ((icmp_ln81_fu_154_p2 == 1'd1) & (icmp_ln78_fu_141_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1)))) begin
        ap_phi_mux_k_9_new_0_i_phi_fu_104_p6 = 16'd0;
    end else begin
        ap_phi_mux_k_9_new_0_i_phi_fu_104_p6 = 'bx;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_0_blk_n = indices_0_full_n;
    end else begin
        indices_0_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_0_write = 1'b1;
    end else begin
        indices_0_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_1_blk_n = indices_1_full_n;
    end else begin
        indices_1_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_1_write = 1'b1;
    end else begin
        indices_1_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_2_out1_blk_n = indices_2_out1_full_n;
    end else begin
        indices_2_out1_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_2_out1_write = 1'b1;
    end else begin
        indices_2_out1_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_2_out_blk_n = indices_2_out_full_n;
    end else begin
        indices_2_out_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_2_out_write = 1'b1;
    end else begin
        indices_2_out_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        internal_ap_ready = 1'b1;
    end else begin
        internal_ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((start_full_n == 1'b0) & (start_once_reg == 1'b0))) begin
        real_start = 1'b0;
    end else begin
        real_start = ap_start;
    end
end

always @ (*) begin
    if (((real_start == 1'b1) & (start_once_reg == 1'b0))) begin
        start_write = 1'b1;
    end else begin
        start_write = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln77_fu_134_p2 = (k_5 + 16'd1);

assign add_ln80_fu_147_p2 = (j_5 + 16'd1);

assign add_ln83_fu_160_p2 = (i_5 + 16'd1);

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

always @ (*) begin
    ap_block_state1 = ((real_start == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1));
end

assign ap_ready = internal_ap_ready;

assign icmp_ln78_fu_141_p2 = ((add_ln77_fu_134_p2 == 16'd1000) ? 1'b1 : 1'b0);

assign icmp_ln81_fu_154_p2 = ((add_ln80_fu_147_p2 == 16'd14) ? 1'b1 : 1'b0);

assign icmp_ln84_fu_166_p2 = ((add_ln83_fu_160_p2 == 16'd14) ? 1'b1 : 1'b0);

assign indices_0_din = i_5;

assign indices_1_din = j_5;

assign indices_2_out1_din = trunc_ln76_fu_128_p1;

assign indices_2_out_din = trunc_ln76_fu_128_p1;

assign select_ln84_fu_172_p3 = ((icmp_ln84_fu_166_p2[0:0] == 1'b1) ? 16'd0 : add_ln83_fu_160_p2);

assign start_out = real_start;

assign trunc_ln76_fu_128_p1 = k_5[9:0];

endmodule //td_fused_top_tdf12_get_next_ijk
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf12_readFilters78 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        filter_data_address0,
        filter_data_ce0,
        filter_data_q0,
        indices_23_dout,
        indices_23_empty_n,
        indices_23_read,
        weight_vecs_0_0_0_address0,
        weight_vecs_0_0_0_ce0,
        weight_vecs_0_0_0_we0,
        weight_vecs_0_0_0_d0
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state6 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [16:0] filter_data_address0;
output   filter_data_ce0;
input  [15:0] filter_data_q0;
input  [9:0] indices_23_dout;
input   indices_23_empty_n;
output   indices_23_read;
output  [6:0] weight_vecs_0_0_0_address0;
output   weight_vecs_0_0_0_ce0;
output   weight_vecs_0_0_0_we0;
output  [15:0] weight_vecs_0_0_0_d0;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg filter_data_ce0;
reg indices_23_read;
reg weight_vecs_0_0_0_ce0;
reg weight_vecs_0_0_0_we0;

reg    ap_done_reg;
  reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    indices_23_blk_n;
reg   [7:0] kk_0_0_i_i_reg_93;
reg   [7:0] kk_0_0_i_i_reg_93_pp0_iter1_reg;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
wire    ap_block_state4_pp0_stage0_iter2;
wire    ap_block_state5_pp0_stage0_iter3;
wire    ap_block_pp0_stage0_11001;
reg   [7:0] kk_0_0_i_i_reg_93_pp0_iter2_reg;
wire   [16:0] tmp_fu_105_p3;
reg   [16:0] tmp_reg_144;
wire   [7:0] add_ln49_fu_113_p2;
reg   [7:0] add_ln49_reg_149;
reg    ap_enable_reg_pp0_iter0;
wire   [0:0] icmp_ln49_fu_119_p2;
reg   [0:0] icmp_ln49_reg_154;
reg   [0:0] icmp_ln49_reg_154_pp0_iter1_reg;
reg   [0:0] icmp_ln49_reg_154_pp0_iter2_reg;
reg    ap_block_state1;
wire    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_exit_iter0_state2;
reg    ap_enable_reg_pp0_iter1;
reg    ap_enable_reg_pp0_iter2;
reg    ap_enable_reg_pp0_iter3;
reg   [7:0] ap_phi_mux_kk_0_0_i_i_phi_fu_97_p4;
wire    ap_block_pp0_stage0;
wire   [63:0] zext_ln55_59_fu_134_p1;
wire   [63:0] idxprom16_0_0_i_i_fu_139_p1;
wire   [16:0] zext_ln55_fu_125_p1;
wire   [16:0] add_ln55_fu_129_p2;
wire    ap_CS_fsm_state6;
reg   [2:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state6)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_condition_pp0_exit_iter0_state2) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            if ((1'b1 == ap_condition_pp0_exit_iter0_state2)) begin
                ap_enable_reg_pp0_iter1 <= (1'b1 ^ ap_condition_pp0_exit_iter0_state2);
            end else if ((1'b1 == 1'b1)) begin
                ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
            end
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end else if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter3 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln49_reg_154 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        kk_0_0_i_i_reg_93 <= add_ln49_reg_149;
    end else if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        kk_0_0_i_i_reg_93 <= 8'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        add_ln49_reg_149 <= add_ln49_fu_113_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln49_reg_154 <= icmp_ln49_fu_119_p2;
        icmp_ln49_reg_154_pp0_iter1_reg <= icmp_ln49_reg_154;
        kk_0_0_i_i_reg_93_pp0_iter1_reg <= kk_0_0_i_i_reg_93;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        icmp_ln49_reg_154_pp0_iter2_reg <= icmp_ln49_reg_154_pp0_iter1_reg;
        kk_0_0_i_i_reg_93_pp0_iter2_reg <= kk_0_0_i_i_reg_93_pp0_iter1_reg;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state1)) begin
        tmp_reg_144[16 : 7] <= tmp_fu_105_p3[16 : 7];
    end
end

always @ (*) begin
    if ((icmp_ln49_fu_119_p2 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state2 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state2 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state6)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln49_reg_154 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_kk_0_0_i_i_phi_fu_97_p4 = add_ln49_reg_149;
    end else begin
        ap_phi_mux_kk_0_0_i_i_phi_fu_97_p4 = kk_0_0_i_i_reg_93;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state6)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter3 == 1'b1)))) begin
        filter_data_ce0 = 1'b1;
    end else begin
        filter_data_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_23_blk_n = indices_23_empty_n;
    end else begin
        indices_23_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_23_read = 1'b1;
    end else begin
        indices_23_read = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter3 == 1'b1))) begin
        weight_vecs_0_0_0_ce0 = 1'b1;
    end else begin
        weight_vecs_0_0_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln49_reg_154_pp0_iter2_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter3 == 1'b1))) begin
        weight_vecs_0_0_0_we0 = 1'b1;
    end else begin
        weight_vecs_0_0_0_we0 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((~((icmp_ln49_fu_119_p2 == 1'd1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter1 == 1'b0)) & ~((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter3 == 1'b1) & (ap_enable_reg_pp0_iter2 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if ((((icmp_ln49_fu_119_p2 == 1'd1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter1 == 1'b0)) | ((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter3 == 1'b1) & (ap_enable_reg_pp0_iter2 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_state6;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state6 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln49_fu_113_p2 = (ap_phi_mux_kk_0_0_i_i_phi_fu_97_p4 + 8'd1);

assign add_ln55_fu_129_p2 = (tmp_reg_144 + zext_ln55_fu_125_p1);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state6 = ap_CS_fsm[32'd2];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1));
end

assign ap_block_state2_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign filter_data_address0 = zext_ln55_59_fu_134_p1;

assign icmp_ln49_fu_119_p2 = ((ap_phi_mux_kk_0_0_i_i_phi_fu_97_p4 == 8'd128) ? 1'b1 : 1'b0);

assign idxprom16_0_0_i_i_fu_139_p1 = kk_0_0_i_i_reg_93_pp0_iter2_reg;

assign tmp_fu_105_p3 = {{indices_23_dout}, {7'd0}};

assign weight_vecs_0_0_0_address0 = idxprom16_0_0_i_i_fu_139_p1;

assign weight_vecs_0_0_0_d0 = filter_data_q0;

assign zext_ln55_59_fu_134_p1 = add_ln55_fu_129_p2;

assign zext_ln55_fu_125_p1 = ap_phi_mux_kk_0_0_i_i_phi_fu_97_p4;

always @ (posedge ap_clk) begin
    tmp_reg_144[6:0] <= 7'b0000000;
end

endmodule //td_fused_top_tdf12_readFilters78
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf12_readInputs (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        in_data_address0,
        in_data_ce0,
        in_data_q0,
        indices_01_dout,
        indices_01_empty_n,
        indices_01_read,
        indices_12_dout,
        indices_12_empty_n,
        indices_12_read,
        ifmap_vec_0_0_address0,
        ifmap_vec_0_0_ce0,
        ifmap_vec_0_0_we0,
        ifmap_vec_0_0_d0,
        ifmap_vec_0_0_address1,
        ifmap_vec_0_0_ce1,
        ifmap_vec_0_0_we1,
        ifmap_vec_0_0_d1,
        indices_01_out_din,
        indices_01_out_full_n,
        indices_01_out_write,
        indices_12_out_din,
        indices_12_out_full_n,
        indices_12_out_write
);

parameter    ap_ST_fsm_state1 = 5'd1;
parameter    ap_ST_fsm_state2 = 5'd2;
parameter    ap_ST_fsm_pp0_stage0 = 5'd4;
parameter    ap_ST_fsm_pp0_stage1 = 5'd8;
parameter    ap_ST_fsm_state8 = 5'd16;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [12:0] in_data_address0;
output   in_data_ce0;
input  [63:0] in_data_q0;
input  [15:0] indices_01_dout;
input   indices_01_empty_n;
output   indices_01_read;
input  [15:0] indices_12_dout;
input   indices_12_empty_n;
output   indices_12_read;
output  [6:0] ifmap_vec_0_0_address0;
output   ifmap_vec_0_0_ce0;
output   ifmap_vec_0_0_we0;
output  [15:0] ifmap_vec_0_0_d0;
output  [6:0] ifmap_vec_0_0_address1;
output   ifmap_vec_0_0_ce1;
output   ifmap_vec_0_0_we1;
output  [15:0] ifmap_vec_0_0_d1;
output  [3:0] indices_01_out_din;
input   indices_01_out_full_n;
output   indices_01_out_write;
output  [7:0] indices_12_out_din;
input   indices_12_out_full_n;
output   indices_12_out_write;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg in_data_ce0;
reg indices_01_read;
reg indices_12_read;
reg[6:0] ifmap_vec_0_0_address0;
reg ifmap_vec_0_0_ce0;
reg ifmap_vec_0_0_we0;
reg[15:0] ifmap_vec_0_0_d0;
reg[6:0] ifmap_vec_0_0_address1;
reg ifmap_vec_0_0_ce1;
reg ifmap_vec_0_0_we1;
reg[15:0] ifmap_vec_0_0_d1;
reg indices_01_out_write;
reg indices_12_out_write;

reg    ap_done_reg;
  reg   [4:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    indices_01_blk_n;
reg    indices_12_blk_n;
reg    indices_01_out_blk_n;
reg    indices_12_out_blk_n;
reg   [7:0] kk_0_i_i_reg_180;
reg   [7:0] kk_0_i_i_reg_180_pp0_iter1_reg;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_block_state3_pp0_stage0_iter0;
wire    ap_block_state5_pp0_stage0_iter1;
wire    ap_block_state7_pp0_stage0_iter2;
wire    ap_block_pp0_stage0_11001;
wire   [3:0] trunc_ln135_fu_192_p1;
reg   [3:0] trunc_ln135_reg_434;
reg   [15:0] col_coord_reg_439;
wire   [0:0] is_padding_fu_214_p2;
reg   [0:0] is_padding_reg_444;
wire   [9:0] add_ln32_fu_274_p2;
reg   [9:0] add_ln32_reg_454;
wire    ap_CS_fsm_state2;
wire   [0:0] icmp_ln25_fu_280_p2;
reg   [0:0] icmp_ln25_reg_459;
reg   [0:0] icmp_ln25_reg_459_pp0_iter1_reg;
wire   [7:0] add_ln25_fu_308_p2;
reg   [7:0] add_ln25_reg_468;
wire    ap_CS_fsm_pp0_stage1;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_state4_pp0_stage1_iter0;
wire    ap_block_state6_pp0_stage1_iter1;
wire    ap_block_pp0_stage1_11001;
wire   [6:0] empty_130_fu_314_p1;
reg   [6:0] empty_130_reg_473;
wire   [15:0] select_ln33_26_fu_386_p3;
reg   [15:0] select_ln33_26_reg_479;
wire   [15:0] select_ln33_27_fu_407_p3;
reg   [15:0] select_ln33_27_reg_484;
wire    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_exit_iter0_state3;
reg    ap_enable_reg_pp0_iter1;
wire    ap_block_pp0_stage1_subdone;
reg    ap_enable_reg_pp0_iter2;
reg   [7:0] ap_phi_mux_kk_0_i_i_phi_fu_184_p4;
wire    ap_block_pp0_stage0;
wire   [63:0] sext_ln32_fu_303_p1;
wire   [63:0] zext_ln32_fu_318_p1;
wire    ap_block_pp0_stage1;
wire   [63:0] zext_ln32_28_fu_345_p1;
wire   [63:0] zext_ln32_29_fu_419_p1;
wire   [63:0] zext_ln32_30_fu_429_p1;
reg    ap_block_state1;
wire   [15:0] select_ln33_fu_331_p3;
wire   [15:0] select_ln33_25_fu_364_p3;
wire   [0:0] cmp7_i_i_fu_202_p2;
wire   [0:0] icmp_ln24_fu_208_p2;
wire   [3:0] empty_128_fu_220_p1;
wire   [3:0] row_coord_int_fu_223_p3;
wire   [7:0] tmp_fu_236_p3;
wire   [4:0] tmp_s_fu_248_p3;
wire   [8:0] zext_ln32_31_fu_244_p1;
wire   [8:0] zext_ln32_32_fu_256_p1;
wire   [8:0] sub_ln32_fu_260_p2;
wire   [3:0] col_coord_int_fu_229_p3;
wire   [9:0] sub_ln32_cast_fu_266_p1;
wire   [9:0] zext_ln32_33_fu_270_p1;
wire   [4:0] lshr_ln_fu_286_p4;
wire   [14:0] tmp_47_fu_296_p3;
wire   [15:0] trunc_ln32_fu_323_p1;
wire   [15:0] bitcast_ln32_fu_327_p1;
wire   [6:0] or_ln25_fu_339_p2;
wire   [15:0] tmp_79_i_i_fu_350_p4;
wire   [15:0] bitcast_ln32_25_fu_360_p1;
wire   [15:0] tmp_80_i_i_fu_372_p4;
wire   [15:0] bitcast_ln32_26_fu_382_p1;
wire   [15:0] tmp_81_i_i_fu_393_p4;
wire   [15:0] bitcast_ln32_27_fu_403_p1;
wire   [6:0] or_ln25_17_fu_414_p2;
wire   [6:0] or_ln25_18_fu_424_p2;
wire    ap_CS_fsm_state8;
reg   [4:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 5'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b1 == ap_condition_pp0_exit_iter0_state3))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1)) | ((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b0)))) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            ap_enable_reg_pp0_iter2 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln25_reg_459 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        kk_0_i_i_reg_180 <= add_ln25_reg_468;
    end else if ((1'b1 == ap_CS_fsm_state2)) begin
        kk_0_i_i_reg_180 <= 8'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln25_reg_459 == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
        add_ln25_reg_468 <= add_ln25_fu_308_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        add_ln32_reg_454 <= add_ln32_fu_274_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state1)) begin
        col_coord_reg_439 <= indices_12_dout;
        is_padding_reg_444 <= is_padding_fu_214_p2;
        trunc_ln135_reg_434 <= trunc_ln135_fu_192_p1;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln25_reg_459_pp0_iter1_reg == 1'd0))) begin
        empty_130_reg_473 <= empty_130_fu_314_p1;
        select_ln33_26_reg_479 <= select_ln33_26_fu_386_p3;
        select_ln33_27_reg_484 <= select_ln33_27_fu_407_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln25_reg_459 <= icmp_ln25_fu_280_p2;
        icmp_ln25_reg_459_pp0_iter1_reg <= icmp_ln25_reg_459;
        kk_0_i_i_reg_180_pp0_iter1_reg <= kk_0_i_i_reg_180;
    end
end

always @ (*) begin
    if ((icmp_ln25_fu_280_p2 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state3 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state3 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state8)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln25_reg_459 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_kk_0_i_i_phi_fu_184_p4 = add_ln25_reg_468;
    end else begin
        ap_phi_mux_kk_0_i_i_phi_fu_184_p4 = kk_0_i_i_reg_180;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state8)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        ifmap_vec_0_0_address0 = zext_ln32_30_fu_429_p1;
    end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ifmap_vec_0_0_address0 = zext_ln32_28_fu_345_p1;
    end else begin
        ifmap_vec_0_0_address0 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        ifmap_vec_0_0_address1 = zext_ln32_29_fu_419_p1;
    end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ifmap_vec_0_0_address1 = zext_ln32_fu_318_p1;
    end else begin
        ifmap_vec_0_0_address1 = 'bx;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1)) | ((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1)))) begin
        ifmap_vec_0_0_ce0 = 1'b1;
    end else begin
        ifmap_vec_0_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1)) | ((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1)))) begin
        ifmap_vec_0_0_ce1 = 1'b1;
    end else begin
        ifmap_vec_0_0_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        ifmap_vec_0_0_d0 = select_ln33_27_reg_484;
    end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ifmap_vec_0_0_d0 = select_ln33_25_fu_364_p3;
    end else begin
        ifmap_vec_0_0_d0 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        ifmap_vec_0_0_d1 = select_ln33_26_reg_479;
    end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ifmap_vec_0_0_d1 = select_ln33_fu_331_p3;
    end else begin
        ifmap_vec_0_0_d1 = 'bx;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1) & (icmp_ln25_reg_459_pp0_iter1_reg == 1'd0)) | ((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln25_reg_459_pp0_iter1_reg == 1'd0)))) begin
        ifmap_vec_0_0_we0 = 1'b1;
    end else begin
        ifmap_vec_0_0_we0 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1) & (icmp_ln25_reg_459_pp0_iter1_reg == 1'd0)) | ((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln25_reg_459_pp0_iter1_reg == 1'd0)))) begin
        ifmap_vec_0_0_we1 = 1'b1;
    end else begin
        ifmap_vec_0_0_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1)) | ((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1)) | ((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1)) | ((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1)))) begin
        in_data_ce0 = 1'b1;
    end else begin
        in_data_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_01_blk_n = indices_01_empty_n;
    end else begin
        indices_01_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_01_out_blk_n = indices_01_out_full_n;
    end else begin
        indices_01_out_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((indices_12_out_full_n == 1'b0) | (indices_01_out_full_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_01_out_write = 1'b1;
    end else begin
        indices_01_out_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((indices_12_out_full_n == 1'b0) | (indices_01_out_full_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_01_read = 1'b1;
    end else begin
        indices_01_read = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_12_blk_n = indices_12_empty_n;
    end else begin
        indices_12_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_12_out_blk_n = indices_12_out_full_n;
    end else begin
        indices_12_out_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((indices_12_out_full_n == 1'b0) | (indices_01_out_full_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_12_out_write = 1'b1;
    end else begin
        indices_12_out_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((indices_12_out_full_n == 1'b0) | (indices_01_out_full_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_12_read = 1'b1;
    end else begin
        indices_12_read = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((indices_12_out_full_n == 1'b0) | (indices_01_out_full_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_state2 : begin
            ap_NS_fsm = ap_ST_fsm_pp0_stage0;
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((~((icmp_ln25_fu_280_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1)) & ~((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0)) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end else if ((((icmp_ln25_fu_280_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1)) | ((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_state8;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_pp0_stage1 : begin
            if ((1'b0 == ap_block_pp0_stage1_subdone)) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end
        end
        ap_ST_fsm_state8 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln25_fu_308_p2 = (kk_0_i_i_reg_180 + 8'd4);

assign add_ln32_fu_274_p2 = ((sub_ln32_cast_fu_266_p1) + (zext_ln32_33_fu_270_p1));

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_pp0_stage1 = ap_CS_fsm[32'd3];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state8 = ap_CS_fsm[32'd4];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((indices_12_out_full_n == 1'b0) | (indices_01_out_full_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0));
end

assign ap_block_state3_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage1_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage1_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign bitcast_ln32_25_fu_360_p1 = tmp_79_i_i_fu_350_p4;

assign bitcast_ln32_26_fu_382_p1 = tmp_80_i_i_fu_372_p4;

assign bitcast_ln32_27_fu_403_p1 = tmp_81_i_i_fu_393_p4;

assign bitcast_ln32_fu_327_p1 = trunc_ln32_fu_323_p1;

assign cmp7_i_i_fu_202_p2 = ((indices_01_dout > 16'd13) ? 1'b1 : 1'b0);

assign col_coord_int_fu_229_p3 = ((is_padding_reg_444[0:0] == 1'b1) ? 4'd0 : empty_128_fu_220_p1);

assign empty_128_fu_220_p1 = col_coord_reg_439[3:0];

assign empty_130_fu_314_p1 = kk_0_i_i_reg_180_pp0_iter1_reg[6:0];

assign icmp_ln24_fu_208_p2 = ((indices_12_dout > 16'd13) ? 1'b1 : 1'b0);

assign icmp_ln25_fu_280_p2 = ((ap_phi_mux_kk_0_i_i_phi_fu_184_p4 == 8'd128) ? 1'b1 : 1'b0);

assign in_data_address0 = sext_ln32_fu_303_p1;

assign indices_01_out_din = indices_01_dout[3:0];

assign indices_12_out_din = indices_12_dout[7:0];

assign is_padding_fu_214_p2 = (icmp_ln24_fu_208_p2 | cmp7_i_i_fu_202_p2);

assign lshr_ln_fu_286_p4 = {{ap_phi_mux_kk_0_i_i_phi_fu_184_p4[6:2]}};

assign or_ln25_17_fu_414_p2 = (empty_130_reg_473 | 7'd2);

assign or_ln25_18_fu_424_p2 = (empty_130_reg_473 | 7'd3);

assign or_ln25_fu_339_p2 = (empty_130_fu_314_p1 | 7'd1);

assign row_coord_int_fu_223_p3 = ((is_padding_reg_444[0:0] == 1'b1) ? 4'd0 : trunc_ln135_reg_434);

assign select_ln33_25_fu_364_p3 = ((is_padding_reg_444[0:0] == 1'b1) ? 16'd0 : bitcast_ln32_25_fu_360_p1);

assign select_ln33_26_fu_386_p3 = ((is_padding_reg_444[0:0] == 1'b1) ? 16'd0 : bitcast_ln32_26_fu_382_p1);

assign select_ln33_27_fu_407_p3 = ((is_padding_reg_444[0:0] == 1'b1) ? 16'd0 : bitcast_ln32_27_fu_403_p1);

assign select_ln33_fu_331_p3 = ((is_padding_reg_444[0:0] == 1'b1) ? 16'd0 : bitcast_ln32_fu_327_p1);

assign sext_ln32_fu_303_p1 = (tmp_47_fu_296_p3);

assign sub_ln32_cast_fu_266_p1 = (sub_ln32_fu_260_p2);

assign sub_ln32_fu_260_p2 = (zext_ln32_31_fu_244_p1 - zext_ln32_32_fu_256_p1);

assign tmp_47_fu_296_p3 = {{add_ln32_reg_454}, {lshr_ln_fu_286_p4}};

assign tmp_79_i_i_fu_350_p4 = {{in_data_q0[31:16]}};

assign tmp_80_i_i_fu_372_p4 = {{in_data_q0[47:32]}};

assign tmp_81_i_i_fu_393_p4 = {{in_data_q0[63:48]}};

assign tmp_fu_236_p3 = {{row_coord_int_fu_223_p3}, {4'd0}};

assign tmp_s_fu_248_p3 = {{row_coord_int_fu_223_p3}, {1'd0}};

assign trunc_ln135_fu_192_p1 = indices_01_dout[3:0];

assign trunc_ln32_fu_323_p1 = in_data_q0[15:0];

assign zext_ln32_28_fu_345_p1 = or_ln25_fu_339_p2;

assign zext_ln32_29_fu_419_p1 = or_ln25_17_fu_414_p2;

assign zext_ln32_30_fu_429_p1 = or_ln25_18_fu_424_p2;

assign zext_ln32_31_fu_244_p1 = tmp_fu_236_p3;

assign zext_ln32_32_fu_256_p1 = tmp_s_fu_248_p3;

assign zext_ln32_33_fu_270_p1 = col_coord_int_fu_229_p3;

assign zext_ln32_fu_318_p1 = kk_0_i_i_reg_180_pp0_iter1_reg;

endmodule //td_fused_top_tdf12_readInputs
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf12_writeOutputs_unaligned (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        indices_01_dout,
        indices_01_empty_n,
        indices_01_read,
        indices_12_dout,
        indices_12_empty_n,
        indices_12_read,
        p_read,
        out_data_address1,
        out_data_ce1,
        out_data_we1,
        out_data_d1
);

parameter    ap_ST_fsm_state1 = 4'd1;
parameter    ap_ST_fsm_state2 = 4'd2;
parameter    ap_ST_fsm_state3 = 4'd4;
parameter    ap_ST_fsm_state4 = 4'd8;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
input  [3:0] indices_01_dout;
input   indices_01_empty_n;
output   indices_01_read;
input  [7:0] indices_12_dout;
input   indices_12_empty_n;
output   indices_12_read;
input  [15:0] p_read;
output  [15:0] out_data_address1;
output   out_data_ce1;
output   out_data_we1;
output  [63:0] out_data_d1;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg indices_01_read;
reg indices_12_read;
reg out_data_ce1;
reg out_data_we1;

reg    ap_done_reg;
  reg   [3:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg   [15:0] outputCount_2;
reg   [15:0] outputChanIdx_2;
reg   [15:0] outputRow_7_0;
reg   [15:0] outputRow_7_1;
reg   [15:0] outputRow_7_2;
reg   [15:0] outputRow_7_3;
reg    indices_01_blk_n;
reg    indices_12_blk_n;
wire   [9:0] add_ln94_fu_157_p2;
reg   [9:0] add_ln94_reg_315;
wire   [15:0] mul_ln89_fu_166_p2;
reg   [15:0] mul_ln89_reg_320;
wire    ap_CS_fsm_state2;
wire   [15:0] add_ln87_fu_204_p2;
wire    ap_CS_fsm_state3;
wire   [0:0] icmp_ln88_fu_210_p2;
reg   [0:0] icmp_ln88_reg_333;
reg   [15:0] ap_phi_mux_empty_phi_fu_112_p4;
reg   [15:0] empty_reg_109;
wire    ap_CS_fsm_state4;
wire   [63:0] zext_ln94_22_fu_237_p1;
wire   [15:0] select_ln97_fu_295_p3;
wire   [1:0] trunc_ln86_fu_176_p1;
reg   [15:0] ap_sig_allocacmp_outputRow_7_0_load;
reg   [15:0] ap_sig_allocacmp_outputRow_7_1_load;
reg   [15:0] ap_sig_allocacmp_outputRow_7_2_load;
reg   [15:0] ap_sig_allocacmp_outputRow_7_3_load;
reg    ap_block_state1;
wire   [7:0] tmp_fu_119_p3;
wire   [4:0] tmp_s_fu_131_p3;
wire   [8:0] zext_ln94_fu_127_p1;
wire   [8:0] zext_ln94_19_fu_139_p1;
wire   [8:0] sub_ln94_fu_143_p2;
wire   [9:0] sub_ln94_cast_fu_149_p1;
wire   [9:0] zext_ln94_20_fu_153_p1;
wire   [8:0] mul_ln89_fu_166_p1;
wire   [8:0] trunc_ln94_fu_224_p1;
wire   [15:0] zext_ln94_21_fu_228_p1;
wire   [15:0] add_ln94_8_fu_232_p2;
wire   [15:0] bitcast_ln94_24_fu_266_p1;
wire   [15:0] bitcast_ln94_23_fu_258_p1;
wire   [15:0] bitcast_ln94_22_fu_250_p1;
wire   [15:0] bitcast_ln94_fu_242_p1;
wire   [15:0] add_ln96_fu_283_p2;
wire   [0:0] icmp_ln97_fu_289_p2;
reg   [3:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 4'd1;
#0 outputCount_2 = 16'd0;
#0 outputChanIdx_2 = 16'd0;
#0 outputRow_7_0 = 16'd0;
#0 outputRow_7_1 = 16'd0;
#0 outputRow_7_2 = 16'd0;
#0 outputRow_7_3 = 16'd0;
end

td_fused_top_mul_10s_9ns_16_1_1 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 10 ),
    .din1_WIDTH( 9 ),
    .dout_WIDTH( 16 ))
mul_10s_9ns_16_1_1_U789(
    .din0(add_ln94_reg_315),
    .din1(mul_ln89_fu_166_p1),
    .dout(mul_ln89_fu_166_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state4)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln88_reg_333 == 1'd1) & (1'b1 == ap_CS_fsm_state4))) begin
        empty_reg_109 <= 16'd0;
    end else if (((icmp_ln88_fu_210_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state3))) begin
        empty_reg_109 <= add_ln87_fu_204_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state1)) begin
        add_ln94_reg_315 <= add_ln94_fu_157_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state3)) begin
        icmp_ln88_reg_333 <= icmp_ln88_fu_210_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        mul_ln89_reg_320 <= mul_ln89_fu_166_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln88_fu_210_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state3))) begin
        outputChanIdx_2 <= select_ln97_fu_295_p3;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        outputCount_2 <= ap_phi_mux_empty_phi_fu_112_p4;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln86_fu_176_p1 == 2'd0) & (1'b1 == ap_CS_fsm_state3))) begin
        outputRow_7_0 <= p_read;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln86_fu_176_p1 == 2'd1) & (1'b1 == ap_CS_fsm_state3))) begin
        outputRow_7_1 <= p_read;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln86_fu_176_p1 == 2'd2) & (1'b1 == ap_CS_fsm_state3))) begin
        outputRow_7_2 <= p_read;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln86_fu_176_p1 == 2'd3) & (1'b1 == ap_CS_fsm_state3))) begin
        outputRow_7_3 <= p_read;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln88_reg_333 == 1'd1) & (1'b1 == ap_CS_fsm_state4))) begin
        ap_phi_mux_empty_phi_fu_112_p4 = 16'd0;
    end else begin
        ap_phi_mux_empty_phi_fu_112_p4 = empty_reg_109;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((trunc_ln86_fu_176_p1 == 2'd0) & (1'b1 == ap_CS_fsm_state3))) begin
        ap_sig_allocacmp_outputRow_7_0_load = p_read;
    end else begin
        ap_sig_allocacmp_outputRow_7_0_load = outputRow_7_0;
    end
end

always @ (*) begin
    if (((trunc_ln86_fu_176_p1 == 2'd1) & (1'b1 == ap_CS_fsm_state3))) begin
        ap_sig_allocacmp_outputRow_7_1_load = p_read;
    end else begin
        ap_sig_allocacmp_outputRow_7_1_load = outputRow_7_1;
    end
end

always @ (*) begin
    if (((trunc_ln86_fu_176_p1 == 2'd2) & (1'b1 == ap_CS_fsm_state3))) begin
        ap_sig_allocacmp_outputRow_7_2_load = p_read;
    end else begin
        ap_sig_allocacmp_outputRow_7_2_load = outputRow_7_2;
    end
end

always @ (*) begin
    if (((trunc_ln86_fu_176_p1 == 2'd3) & (1'b1 == ap_CS_fsm_state3))) begin
        ap_sig_allocacmp_outputRow_7_3_load = p_read;
    end else begin
        ap_sig_allocacmp_outputRow_7_3_load = outputRow_7_3;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_01_blk_n = indices_01_empty_n;
    end else begin
        indices_01_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_01_read = 1'b1;
    end else begin
        indices_01_read = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_12_blk_n = indices_12_empty_n;
    end else begin
        indices_12_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_12_read = 1'b1;
    end else begin
        indices_12_read = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state3))) begin
        out_data_ce1 = 1'b1;
    end else begin
        out_data_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln88_fu_210_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state3))) begin
        out_data_we1 = 1'b1;
    end else begin
        out_data_we1 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_start == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_state2 : begin
            ap_NS_fsm = ap_ST_fsm_state3;
        end
        ap_ST_fsm_state3 : begin
            ap_NS_fsm = ap_ST_fsm_state4;
        end
        ap_ST_fsm_state4 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln87_fu_204_p2 = (outputCount_2 + 16'd1);

assign add_ln94_8_fu_232_p2 = (mul_ln89_reg_320 + zext_ln94_21_fu_228_p1);

assign add_ln94_fu_157_p2 = ((sub_ln94_cast_fu_149_p1) + (zext_ln94_20_fu_153_p1));

assign add_ln96_fu_283_p2 = (outputChanIdx_2 + 16'd1);

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1));
end

assign bitcast_ln94_22_fu_250_p1 = ap_sig_allocacmp_outputRow_7_1_load;

assign bitcast_ln94_23_fu_258_p1 = ap_sig_allocacmp_outputRow_7_2_load;

assign bitcast_ln94_24_fu_266_p1 = ap_sig_allocacmp_outputRow_7_3_load;

assign bitcast_ln94_fu_242_p1 = ap_sig_allocacmp_outputRow_7_0_load;

assign icmp_ln88_fu_210_p2 = ((add_ln87_fu_204_p2 == 16'd4) ? 1'b1 : 1'b0);

assign icmp_ln97_fu_289_p2 = ((add_ln96_fu_283_p2 == 16'd250) ? 1'b1 : 1'b0);

assign mul_ln89_fu_166_p1 = 16'd250;

assign out_data_address1 = zext_ln94_22_fu_237_p1;

assign out_data_d1 = {{{{bitcast_ln94_24_fu_266_p1}, {bitcast_ln94_23_fu_258_p1}}, {bitcast_ln94_22_fu_250_p1}}, {bitcast_ln94_fu_242_p1}};

assign select_ln97_fu_295_p3 = ((icmp_ln97_fu_289_p2[0:0] == 1'b1) ? 16'd0 : add_ln96_fu_283_p2);

assign sub_ln94_cast_fu_149_p1 = (sub_ln94_fu_143_p2);

assign sub_ln94_fu_143_p2 = (zext_ln94_fu_127_p1 - zext_ln94_19_fu_139_p1);

assign tmp_fu_119_p3 = {{indices_01_dout}, {4'd0}};

assign tmp_s_fu_131_p3 = {{indices_01_dout}, {1'd0}};

assign trunc_ln86_fu_176_p1 = outputCount_2[1:0];

assign trunc_ln94_fu_224_p1 = outputChanIdx_2[8:0];

assign zext_ln94_19_fu_139_p1 = tmp_s_fu_131_p3;

assign zext_ln94_20_fu_153_p1 = indices_12_dout;

assign zext_ln94_21_fu_228_p1 = trunc_ln94_fu_224_p1;

assign zext_ln94_22_fu_237_p1 = add_ln94_8_fu_232_p2;

assign zext_ln94_fu_127_p1 = tmp_fu_119_p3;

endmodule //td_fused_top_tdf12_writeOutputs_unaligned
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf1_accum_1 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        accum_in_0_address0,
        accum_in_0_ce0,
        accum_in_0_q0,
        accum_in_0_address1,
        accum_in_0_ce1,
        accum_in_0_q1,
        accum_out_address0,
        accum_out_ce0,
        accum_out_we0,
        accum_out_d0
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state9 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [4:0] accum_in_0_address0;
output   accum_in_0_ce0;
input  [15:0] accum_in_0_q0;
output  [4:0] accum_in_0_address1;
output   accum_in_0_ce1;
input  [15:0] accum_in_0_q1;
output  [3:0] accum_out_address0;
output   accum_out_ce0;
output   accum_out_we0;
output  [15:0] accum_out_d0;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg accum_in_0_ce0;
reg accum_in_0_ce1;
reg accum_out_ce0;
reg accum_out_we0;

reg    ap_done_reg;
  reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg   [3:0] out_idx_reg_76;
reg   [3:0] out_idx_reg_76_pp0_iter1_reg;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
wire    ap_block_state4_pp0_stage0_iter2;
wire    ap_block_state5_pp0_stage0_iter3;
wire    ap_block_state6_pp0_stage0_iter4;
wire    ap_block_state7_pp0_stage0_iter5;
wire    ap_block_state8_pp0_stage0_iter6;
wire    ap_block_pp0_stage0_11001;
reg   [3:0] out_idx_reg_76_pp0_iter2_reg;
reg   [3:0] out_idx_reg_76_pp0_iter3_reg;
reg   [3:0] out_idx_reg_76_pp0_iter4_reg;
reg   [3:0] out_idx_reg_76_pp0_iter5_reg;
wire   [3:0] add_ln59_fu_94_p2;
reg   [3:0] add_ln59_reg_147;
reg    ap_enable_reg_pp0_iter0;
wire   [0:0] icmp_ln45_fu_100_p2;
reg   [0:0] icmp_ln45_reg_152;
reg   [0:0] icmp_ln45_reg_152_pp0_iter1_reg;
reg   [0:0] icmp_ln45_reg_152_pp0_iter2_reg;
reg   [0:0] icmp_ln45_reg_152_pp0_iter3_reg;
reg   [0:0] icmp_ln45_reg_152_pp0_iter4_reg;
reg   [0:0] icmp_ln45_reg_152_pp0_iter5_reg;
wire   [4:0] i_1_1_fu_106_p3;
reg   [4:0] i_1_1_reg_156;
wire   [0:0] icmp_ln55_fu_120_p2;
reg   [0:0] icmp_ln55_reg_161;
wire   [15:0] select_ln55_fu_135_p3;
reg   [15:0] select_ln55_reg_176;
reg    ap_enable_reg_pp0_iter2;
reg    ap_block_state1;
wire    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_exit_iter0_state2;
reg    ap_enable_reg_pp0_iter1;
reg    ap_enable_reg_pp0_iter3;
reg    ap_enable_reg_pp0_iter4;
reg    ap_enable_reg_pp0_iter5;
reg    ap_enable_reg_pp0_iter6;
reg   [3:0] ap_phi_mux_out_idx_phi_fu_80_p4;
wire    ap_block_pp0_stage0;
wire   [63:0] zext_ln55_1_fu_126_p1;
wire   [63:0] zext_ln55_fu_131_p1;
wire   [63:0] zext_ln45_fu_142_p1;
wire   [15:0] grp_fu_88_p2;
wire   [4:0] or_ln55_fu_114_p2;
wire    ap_CS_fsm_state9;
reg   [2:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
#0 ap_enable_reg_pp0_iter4 = 1'b0;
#0 ap_enable_reg_pp0_iter5 = 1'b0;
#0 ap_enable_reg_pp0_iter6 = 1'b0;
end

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U25(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(select_ln55_reg_176),
    .din1(accum_in_0_q0),
    .dout(grp_fu_88_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b1 == ap_condition_pp0_exit_iter0_state2))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            if ((1'b1 == ap_condition_pp0_exit_iter0_state2)) begin
                ap_enable_reg_pp0_iter1 <= (1'b1 ^ ap_condition_pp0_exit_iter0_state2);
            end else if ((1'b1 == 1'b1)) begin
                ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
            end
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter4 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter5 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter5 <= ap_enable_reg_pp0_iter4;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter6 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter6 <= ap_enable_reg_pp0_iter5;
        end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter6 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        out_idx_reg_76 <= 4'd0;
    end else if (((icmp_ln45_reg_152 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        out_idx_reg_76 <= add_ln59_reg_147;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        add_ln59_reg_147 <= add_ln59_fu_94_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln45_fu_100_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        i_1_1_reg_156[4 : 1] <= i_1_1_fu_106_p3[4 : 1];
        icmp_ln55_reg_161 <= icmp_ln55_fu_120_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln45_reg_152 <= icmp_ln45_fu_100_p2;
        icmp_ln45_reg_152_pp0_iter1_reg <= icmp_ln45_reg_152;
        out_idx_reg_76_pp0_iter1_reg <= out_idx_reg_76;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        icmp_ln45_reg_152_pp0_iter2_reg <= icmp_ln45_reg_152_pp0_iter1_reg;
        icmp_ln45_reg_152_pp0_iter3_reg <= icmp_ln45_reg_152_pp0_iter2_reg;
        icmp_ln45_reg_152_pp0_iter4_reg <= icmp_ln45_reg_152_pp0_iter3_reg;
        icmp_ln45_reg_152_pp0_iter5_reg <= icmp_ln45_reg_152_pp0_iter4_reg;
        out_idx_reg_76_pp0_iter2_reg <= out_idx_reg_76_pp0_iter1_reg;
        out_idx_reg_76_pp0_iter3_reg <= out_idx_reg_76_pp0_iter2_reg;
        out_idx_reg_76_pp0_iter4_reg <= out_idx_reg_76_pp0_iter3_reg;
        out_idx_reg_76_pp0_iter5_reg <= out_idx_reg_76_pp0_iter4_reg;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln45_reg_152 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        select_ln55_reg_176 <= select_ln55_fu_135_p3;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        accum_in_0_ce0 = 1'b1;
    end else begin
        accum_in_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        accum_in_0_ce1 = 1'b1;
    end else begin
        accum_in_0_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter6 == 1'b1))) begin
        accum_out_ce0 = 1'b1;
    end else begin
        accum_out_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln45_reg_152_pp0_iter5_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter6 == 1'b1))) begin
        accum_out_we0 = 1'b1;
    end else begin
        accum_out_we0 = 1'b0;
    end
end

always @ (*) begin
    if ((icmp_ln45_fu_100_p2 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state2 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state2 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state9)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln45_reg_152 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_out_idx_phi_fu_80_p4 = add_ln59_reg_147;
    end else begin
        ap_phi_mux_out_idx_phi_fu_80_p4 = out_idx_reg_76;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state9)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((~((icmp_ln45_fu_100_p2 == 1'd1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter1 == 1'b0)) & ~((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter6 == 1'b1) & (ap_enable_reg_pp0_iter5 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if ((((icmp_ln45_fu_100_p2 == 1'd1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter1 == 1'b0)) | ((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter6 == 1'b1) & (ap_enable_reg_pp0_iter5 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_state9;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state9 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign accum_in_0_address0 = zext_ln55_fu_131_p1;

assign accum_in_0_address1 = zext_ln55_1_fu_126_p1;

assign accum_out_address0 = zext_ln45_fu_142_p1;

assign accum_out_d0 = grp_fu_88_p2;

assign add_ln59_fu_94_p2 = (ap_phi_mux_out_idx_phi_fu_80_p4 + 4'd1);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state9 = ap_CS_fsm[32'd2];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (ap_done_reg == 1'b1));
end

assign ap_block_state2_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter4 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage0_iter5 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage0_iter6 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign i_1_1_fu_106_p3 = {{ap_phi_mux_out_idx_phi_fu_80_p4}, {1'd0}};

assign icmp_ln45_fu_100_p2 = ((ap_phi_mux_out_idx_phi_fu_80_p4 == 4'd14) ? 1'b1 : 1'b0);

assign icmp_ln55_fu_120_p2 = ((or_ln55_fu_114_p2 < 5'd27) ? 1'b1 : 1'b0);

assign or_ln55_fu_114_p2 = (i_1_1_fu_106_p3 | 5'd1);

assign select_ln55_fu_135_p3 = ((icmp_ln55_reg_161[0:0] == 1'b1) ? accum_in_0_q1 : 16'd0);

assign zext_ln45_fu_142_p1 = out_idx_reg_76_pp0_iter5_reg;

assign zext_ln55_1_fu_126_p1 = or_ln55_fu_114_p2;

assign zext_ln55_fu_131_p1 = i_1_1_reg_156;

always @ (posedge ap_clk) begin
    i_1_1_reg_156[0] <= 1'b0;
end

endmodule //td_fused_top_tdf1_accum_1
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf1_accum_2 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        accum_in_address0,
        accum_in_ce0,
        accum_in_q0,
        accum_in_address1,
        accum_in_ce1,
        accum_in_q1,
        accum_out_address0,
        accum_out_ce0,
        accum_out_we0,
        accum_out_d0
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state8 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [3:0] accum_in_address0;
output   accum_in_ce0;
input  [15:0] accum_in_q0;
output  [3:0] accum_in_address1;
output   accum_in_ce1;
input  [15:0] accum_in_q1;
output  [2:0] accum_out_address0;
output   accum_out_ce0;
output   accum_out_we0;
output  [15:0] accum_out_d0;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg accum_in_ce0;
reg accum_in_ce1;
reg accum_out_ce0;
reg accum_out_we0;

reg    ap_done_reg;
  reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg   [2:0] out_idx_reg_72;
reg   [2:0] out_idx_reg_72_pp0_iter1_reg;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
wire    ap_block_state4_pp0_stage0_iter2;
wire    ap_block_state5_pp0_stage0_iter3;
wire    ap_block_state6_pp0_stage0_iter4;
wire    ap_block_state7_pp0_stage0_iter5;
wire    ap_block_pp0_stage0_11001;
reg   [2:0] out_idx_reg_72_pp0_iter2_reg;
reg   [2:0] out_idx_reg_72_pp0_iter3_reg;
reg   [2:0] out_idx_reg_72_pp0_iter4_reg;
wire   [2:0] add_ln89_fu_91_p2;
reg   [2:0] add_ln89_reg_132;
reg    ap_enable_reg_pp0_iter0;
wire   [0:0] icmp_ln75_fu_97_p2;
reg   [0:0] icmp_ln75_reg_137;
reg   [0:0] icmp_ln75_reg_137_pp0_iter1_reg;
reg   [0:0] icmp_ln75_reg_137_pp0_iter2_reg;
reg   [0:0] icmp_ln75_reg_137_pp0_iter3_reg;
reg   [0:0] icmp_ln75_reg_137_pp0_iter4_reg;
reg    ap_enable_reg_pp0_iter1;
reg    ap_block_state1;
wire    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_exit_iter0_state2;
reg    ap_enable_reg_pp0_iter2;
reg    ap_enable_reg_pp0_iter3;
reg    ap_enable_reg_pp0_iter4;
reg    ap_enable_reg_pp0_iter5;
reg   [2:0] ap_phi_mux_out_idx_phi_fu_76_p4;
wire    ap_block_pp0_stage0;
wire   [63:0] zext_ln85_fu_111_p1;
wire   [63:0] zext_ln85_1_fu_122_p1;
wire   [63:0] zext_ln75_fu_127_p1;
wire   [15:0] grp_fu_84_p2;
wire   [3:0] i_1_1_fu_103_p3;
wire   [3:0] or_ln85_fu_116_p2;
wire    ap_CS_fsm_state8;
reg   [2:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
#0 ap_enable_reg_pp0_iter4 = 1'b0;
#0 ap_enable_reg_pp0_iter5 = 1'b0;
end

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U29(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(accum_in_q0),
    .din1(accum_in_q1),
    .dout(grp_fu_84_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b1 == ap_condition_pp0_exit_iter0_state2))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            if ((1'b1 == ap_condition_pp0_exit_iter0_state2)) begin
                ap_enable_reg_pp0_iter1 <= (1'b1 ^ ap_condition_pp0_exit_iter0_state2);
            end else if ((1'b1 == 1'b1)) begin
                ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
            end
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter4 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter5 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter5 <= ap_enable_reg_pp0_iter4;
        end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter5 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        out_idx_reg_72 <= 3'd0;
    end else if (((ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln75_reg_137 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        out_idx_reg_72 <= add_ln89_reg_132;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        add_ln89_reg_132 <= add_ln89_fu_91_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln75_reg_137 <= icmp_ln75_fu_97_p2;
        icmp_ln75_reg_137_pp0_iter1_reg <= icmp_ln75_reg_137;
        out_idx_reg_72_pp0_iter1_reg <= out_idx_reg_72;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        icmp_ln75_reg_137_pp0_iter2_reg <= icmp_ln75_reg_137_pp0_iter1_reg;
        icmp_ln75_reg_137_pp0_iter3_reg <= icmp_ln75_reg_137_pp0_iter2_reg;
        icmp_ln75_reg_137_pp0_iter4_reg <= icmp_ln75_reg_137_pp0_iter3_reg;
        out_idx_reg_72_pp0_iter2_reg <= out_idx_reg_72_pp0_iter1_reg;
        out_idx_reg_72_pp0_iter3_reg <= out_idx_reg_72_pp0_iter2_reg;
        out_idx_reg_72_pp0_iter4_reg <= out_idx_reg_72_pp0_iter3_reg;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        accum_in_ce0 = 1'b1;
    end else begin
        accum_in_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        accum_in_ce1 = 1'b1;
    end else begin
        accum_in_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter5 == 1'b1))) begin
        accum_out_ce0 = 1'b1;
    end else begin
        accum_out_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln75_reg_137_pp0_iter4_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter5 == 1'b1))) begin
        accum_out_we0 = 1'b1;
    end else begin
        accum_out_we0 = 1'b0;
    end
end

always @ (*) begin
    if ((icmp_ln75_fu_97_p2 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state2 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state2 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state8)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln75_reg_137 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_phi_mux_out_idx_phi_fu_76_p4 = add_ln89_reg_132;
    end else begin
        ap_phi_mux_out_idx_phi_fu_76_p4 = out_idx_reg_72;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state8)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((~((ap_enable_reg_pp0_iter1 == 1'b0) & (icmp_ln75_fu_97_p2 == 1'd1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone)) & ~((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter5 == 1'b1) & (ap_enable_reg_pp0_iter4 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if ((((ap_enable_reg_pp0_iter1 == 1'b0) & (icmp_ln75_fu_97_p2 == 1'd1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone)) | ((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter5 == 1'b1) & (ap_enable_reg_pp0_iter4 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_state8;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state8 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign accum_in_address0 = zext_ln85_1_fu_122_p1;

assign accum_in_address1 = zext_ln85_fu_111_p1;

assign accum_out_address0 = zext_ln75_fu_127_p1;

assign accum_out_d0 = grp_fu_84_p2;

assign add_ln89_fu_91_p2 = (ap_phi_mux_out_idx_phi_fu_76_p4 + 3'd1);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state8 = ap_CS_fsm[32'd2];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (ap_done_reg == 1'b1));
end

assign ap_block_state2_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter4 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage0_iter5 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign i_1_1_fu_103_p3 = {{ap_phi_mux_out_idx_phi_fu_76_p4}, {1'd0}};

assign icmp_ln75_fu_97_p2 = ((ap_phi_mux_out_idx_phi_fu_76_p4 == 3'd7) ? 1'b1 : 1'b0);

assign or_ln85_fu_116_p2 = (i_1_1_fu_103_p3 | 4'd1);

assign zext_ln75_fu_127_p1 = out_idx_reg_72_pp0_iter4_reg;

assign zext_ln85_1_fu_122_p1 = or_ln85_fu_116_p2;

assign zext_ln85_fu_111_p1 = i_1_1_fu_103_p3;

endmodule //td_fused_top_tdf1_accum_2
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf1_accum_3 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        accum_in_18,
        accum_in_18_ap_vld,
        accum_in_address0,
        accum_in_ce0,
        accum_in_q0
);

parameter    ap_ST_fsm_state1 = 7'd1;
parameter    ap_ST_fsm_state2 = 7'd2;
parameter    ap_ST_fsm_state3 = 7'd4;
parameter    ap_ST_fsm_state4 = 7'd8;
parameter    ap_ST_fsm_state5 = 7'd16;
parameter    ap_ST_fsm_state6 = 7'd32;
parameter    ap_ST_fsm_state7 = 7'd64;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [15:0] accum_in_18;
output   accum_in_18_ap_vld;
output  [2:0] accum_in_address0;
output   accum_in_ce0;
input  [15:0] accum_in_q0;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg[15:0] accum_in_18;
reg accum_in_18_ap_vld;
reg accum_in_ce0;

reg    ap_done_reg;
  reg   [6:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
wire   [2:0] add_ln102_fu_74_p2;
reg   [2:0] add_ln102_reg_91;
wire    ap_CS_fsm_state2;
wire   [0:0] icmp_ln102_fu_85_p2;
wire    ap_CS_fsm_state3;
wire   [15:0] grp_fu_68_p2;
wire    ap_CS_fsm_state7;
reg   [2:0] i_1_1_reg_44;
reg    ap_block_state1;
reg   [15:0] sum_01_reg_55;
wire   [63:0] zext_ln102_fu_80_p1;
reg   [15:0] accum_in_18_preg;
reg   [6:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 7'd1;
#0 accum_in_18_preg = 16'd0;
end

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U32(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(sum_01_reg_55),
    .din1(accum_in_q0),
    .dout(grp_fu_68_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        accum_in_18_preg <= 16'd0;
    end else begin
        if (((icmp_ln102_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
            accum_in_18_preg <= sum_01_reg_55;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if (((icmp_ln102_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        i_1_1_reg_44 <= 3'd0;
    end else if ((1'b1 == ap_CS_fsm_state7)) begin
        i_1_1_reg_44 <= add_ln102_reg_91;
    end
end

always @ (posedge ap_clk) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        sum_01_reg_55 <= 16'd0;
    end else if ((1'b1 == ap_CS_fsm_state7)) begin
        sum_01_reg_55 <= grp_fu_68_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        add_ln102_reg_91 <= add_ln102_fu_74_p2;
    end
end

always @ (*) begin
    if (((icmp_ln102_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        accum_in_18 = sum_01_reg_55;
    end else begin
        accum_in_18 = accum_in_18_preg;
    end
end

always @ (*) begin
    if (((icmp_ln102_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        accum_in_18_ap_vld = 1'b1;
    end else begin
        accum_in_18_ap_vld = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        accum_in_ce0 = 1'b1;
    end else begin
        accum_in_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln102_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln102_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_state2 : begin
            if (((icmp_ln102_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end
        end
        ap_ST_fsm_state3 : begin
            ap_NS_fsm = ap_ST_fsm_state4;
        end
        ap_ST_fsm_state4 : begin
            ap_NS_fsm = ap_ST_fsm_state5;
        end
        ap_ST_fsm_state5 : begin
            ap_NS_fsm = ap_ST_fsm_state6;
        end
        ap_ST_fsm_state6 : begin
            ap_NS_fsm = ap_ST_fsm_state7;
        end
        ap_ST_fsm_state7 : begin
            ap_NS_fsm = ap_ST_fsm_state2;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign accum_in_address0 = zext_ln102_fu_80_p1;

assign add_ln102_fu_74_p2 = (i_1_1_reg_44 + 3'd1);

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state7 = ap_CS_fsm[32'd6];

always @ (*) begin
    ap_block_state1 = ((ap_done_reg == 1'b1) | (ap_start == 1'b0));
end

assign icmp_ln102_fu_85_p2 = ((i_1_1_reg_44 == 3'd7) ? 1'b1 : 1'b0);

assign zext_ln102_fu_80_p1 = i_1_1_reg_44;

endmodule //td_fused_top_tdf1_accum_3
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_tdf1_adjustments_ram (addr0, ce0, q0, addr1, ce1, d1, we1,  clk);

parameter DWIDTH = 48;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
output wire[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
input clk;

 reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];
wire [AWIDTH-1:0] addr0_t0; 
reg [AWIDTH-1:0] addr0_t1; 
reg [DWIDTH-1:0] q0_t0;
reg [DWIDTH-1:0] q0_t1;
wire [AWIDTH-1:0] addr1_t0; 
reg [AWIDTH-1:0] addr1_t1; 
wire [DWIDTH-1:0] d1_t0; 
wire we1_t0; 
reg [DWIDTH-1:0] d1_t1; 
reg we1_t1; 


assign addr0_t0 = addr0;
assign q0 = q0_t1;
assign addr1_t0 = addr1;
assign d1_t0 = d1;
assign we1_t0 = we1;

always @(posedge clk)  
begin
    if (ce0) 
    begin
        addr0_t1 <= addr0_t0; 
        q0_t1 <= q0_t0;
    end
    if (ce1) 
    begin
        addr1_t1 <= addr1_t0; 
        d1_t1 <= d1_t0;
        we1_t1 <= we1_t0;
    end
end


always @(posedge clk)  
begin 
    if (ce0) begin
        q0_t0 <= ram[addr0_t1];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1_t1) 
            ram[addr1_t1] <= d1_t1; 
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_tdf1_adjustments(
    reset,
    clk,
    address0,
    ce0,
    q0,
    address1,
    ce1,
    we1,
    d1);

parameter DataWidth = 32'd48;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;



td_fused_top_tdf1_adjustments_ram td_fused_top_tdf1_adjustments_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 )
);

endmodule

// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf1_adjust (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        sums_read,
        adjustments_address0,
        adjustments_ce0,
        adjustments_q0,
        input_indices_23_dout,
        input_indices_23_empty_n,
        input_indices_23_read,
        ap_return
);

parameter    ap_ST_fsm_state1 = 17'd1;
parameter    ap_ST_fsm_state2 = 17'd2;
parameter    ap_ST_fsm_state3 = 17'd4;
parameter    ap_ST_fsm_state4 = 17'd8;
parameter    ap_ST_fsm_state5 = 17'd16;
parameter    ap_ST_fsm_state6 = 17'd32;
parameter    ap_ST_fsm_state7 = 17'd64;
parameter    ap_ST_fsm_state8 = 17'd128;
parameter    ap_ST_fsm_state9 = 17'd256;
parameter    ap_ST_fsm_state10 = 17'd512;
parameter    ap_ST_fsm_state11 = 17'd1024;
parameter    ap_ST_fsm_state12 = 17'd2048;
parameter    ap_ST_fsm_state13 = 17'd4096;
parameter    ap_ST_fsm_state14 = 17'd8192;
parameter    ap_ST_fsm_state15 = 17'd16384;
parameter    ap_ST_fsm_state16 = 17'd32768;
parameter    ap_ST_fsm_state17 = 17'd65536;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
input  [15:0] sums_read;
output  [3:0] adjustments_address0;
output   adjustments_ce0;
input  [47:0] adjustments_q0;
input  [3:0] input_indices_23_dout;
input   input_indices_23_empty_n;
output   input_indices_23_read;
output  [15:0] ap_return;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg adjustments_ce0;
reg input_indices_23_read;

reg    ap_done_reg;
  reg   [16:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    input_indices_23_blk_n;
wire    ap_CS_fsm_state4;
reg   [15:0] tmp_74_i_i_reg_167;
reg   [15:0] tmp_75_i_i_reg_172;
wire   [15:0] grp_fu_81_p2;
reg   [15:0] sub_i_i_i_reg_177;
wire    ap_CS_fsm_state8;
wire    ap_CS_fsm_state9;
wire   [15:0] grp_fu_86_p2;
reg   [15:0] mul_i_i_i_reg_187;
wire    ap_CS_fsm_state12;
wire    ap_CS_fsm_state13;
wire   [63:0] zext_ln220_fu_90_p1;
reg    ap_block_state1;
wire    ap_CS_fsm_state2;
wire    ap_CS_fsm_state3;
wire   [15:0] grp_fu_77_p1;
wire   [15:0] grp_fu_81_p1;
wire   [15:0] grp_fu_86_p1;
wire   [15:0] trunc_ln220_fu_95_p1;
wire   [15:0] grp_fu_77_p2;
wire    ap_CS_fsm_state17;
wire   [15:0] bitcast_ln648_fu_132_p1;
wire   [0:0] tmp_fu_136_p3;
reg   [16:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 17'd1;
end

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U36(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(mul_i_i_i_reg_187),
    .din1(grp_fu_77_p1),
    .dout(grp_fu_77_p2)
);

td_fused_top_hsub_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hsub_16ns_16ns_16_5_full_dsp_1_U37(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(sums_read),
    .din1(grp_fu_81_p1),
    .dout(grp_fu_81_p2)
);

td_fused_top_hmul_16ns_16ns_16_4_max_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hmul_16ns_16ns_16_4_max_dsp_1_U38(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(sub_i_i_i_reg_177),
    .din1(grp_fu_86_p1),
    .dout(grp_fu_86_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state17)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state12)) begin
        mul_i_i_i_reg_187 <= grp_fu_86_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state8)) begin
        sub_i_i_i_reg_177 <= grp_fu_81_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        tmp_74_i_i_reg_167 <= {{adjustments_q0[31:16]}};
        tmp_75_i_i_reg_172 <= {{adjustments_q0[47:32]}};
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state2) | (~((input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1)))) begin
        adjustments_ce0 = 1'b1;
    end else begin
        adjustments_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state17)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state17)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        input_indices_23_blk_n = input_indices_23_empty_n;
    end else begin
        input_indices_23_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        input_indices_23_read = 1'b1;
    end else begin
        input_indices_23_read = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_state2 : begin
            ap_NS_fsm = ap_ST_fsm_state3;
        end
        ap_ST_fsm_state3 : begin
            ap_NS_fsm = ap_ST_fsm_state4;
        end
        ap_ST_fsm_state4 : begin
            ap_NS_fsm = ap_ST_fsm_state5;
        end
        ap_ST_fsm_state5 : begin
            ap_NS_fsm = ap_ST_fsm_state6;
        end
        ap_ST_fsm_state6 : begin
            ap_NS_fsm = ap_ST_fsm_state7;
        end
        ap_ST_fsm_state7 : begin
            ap_NS_fsm = ap_ST_fsm_state8;
        end
        ap_ST_fsm_state8 : begin
            ap_NS_fsm = ap_ST_fsm_state9;
        end
        ap_ST_fsm_state9 : begin
            ap_NS_fsm = ap_ST_fsm_state10;
        end
        ap_ST_fsm_state10 : begin
            ap_NS_fsm = ap_ST_fsm_state11;
        end
        ap_ST_fsm_state11 : begin
            ap_NS_fsm = ap_ST_fsm_state12;
        end
        ap_ST_fsm_state12 : begin
            ap_NS_fsm = ap_ST_fsm_state13;
        end
        ap_ST_fsm_state13 : begin
            ap_NS_fsm = ap_ST_fsm_state14;
        end
        ap_ST_fsm_state14 : begin
            ap_NS_fsm = ap_ST_fsm_state15;
        end
        ap_ST_fsm_state15 : begin
            ap_NS_fsm = ap_ST_fsm_state16;
        end
        ap_ST_fsm_state16 : begin
            ap_NS_fsm = ap_ST_fsm_state17;
        end
        ap_ST_fsm_state17 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign adjustments_address0 = zext_ln220_fu_90_p1;

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state12 = ap_CS_fsm[32'd11];

assign ap_CS_fsm_state13 = ap_CS_fsm[32'd12];

assign ap_CS_fsm_state17 = ap_CS_fsm[32'd16];

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

assign ap_CS_fsm_state8 = ap_CS_fsm[32'd7];

assign ap_CS_fsm_state9 = ap_CS_fsm[32'd8];

always @ (*) begin
    ap_block_state1 = ((input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0));
end

assign ap_return = ((tmp_fu_136_p3[0:0] == 1'b1) ? 16'd0 : grp_fu_77_p2);

assign bitcast_ln648_fu_132_p1 = grp_fu_77_p2;

assign grp_fu_77_p1 = tmp_75_i_i_reg_172;

assign grp_fu_81_p1 = trunc_ln220_fu_95_p1;

assign grp_fu_86_p1 = tmp_74_i_i_reg_167;

assign tmp_fu_136_p3 = bitcast_ln648_fu_132_p1[32'd15];

assign trunc_ln220_fu_95_p1 = adjustments_q0[15:0];

assign zext_ln220_fu_90_p1 = input_indices_23_dout;

endmodule //td_fused_top_tdf1_adjust
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf1_dot_product (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        ifmap_vec_address0,
        ifmap_vec_ce0,
        ifmap_vec_q0,
        weight_vecs_0_address0,
        weight_vecs_0_ce0,
        weight_vecs_0_q0,
        products_0_address0,
        products_0_ce0,
        products_0_we0,
        products_0_d0
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state8 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [4:0] ifmap_vec_address0;
output   ifmap_vec_ce0;
input  [15:0] ifmap_vec_q0;
output  [4:0] weight_vecs_0_address0;
output   weight_vecs_0_ce0;
input  [15:0] weight_vecs_0_q0;
output  [4:0] products_0_address0;
output   products_0_ce0;
output   products_0_we0;
output  [15:0] products_0_d0;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg ifmap_vec_ce0;
reg weight_vecs_0_ce0;
reg products_0_ce0;
reg products_0_we0;

reg    ap_done_reg;
  reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg   [4:0] indvar_flatten21_reg_93;
reg   [1:0] ii_reg_104;
reg   [3:0] indvar_flatten_reg_116;
reg   [1:0] jj_reg_127;
reg   [1:0] ic_reg_138;
wire   [4:0] add_ln147_6_fu_156_p2;
wire    ap_CS_fsm_pp0_stage0;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
wire    ap_block_state4_pp0_stage0_iter2;
wire    ap_block_state5_pp0_stage0_iter3;
wire    ap_block_state6_pp0_stage0_iter4;
wire    ap_block_state7_pp0_stage0_iter5;
wire    ap_block_pp0_stage0_11001;
wire   [0:0] icmp_ln147_fu_162_p2;
reg   [0:0] icmp_ln147_reg_466;
reg   [0:0] icmp_ln147_reg_466_pp0_iter1_reg;
reg   [0:0] icmp_ln147_reg_466_pp0_iter2_reg;
reg   [0:0] icmp_ln147_reg_466_pp0_iter3_reg;
reg   [0:0] icmp_ln147_reg_466_pp0_iter4_reg;
wire   [1:0] add_ln147_fu_168_p2;
reg   [1:0] add_ln147_reg_470;
wire   [0:0] icmp_ln148_fu_174_p2;
reg   [0:0] icmp_ln148_reg_476;
wire   [1:0] select_ln147_17_fu_180_p3;
reg   [1:0] select_ln147_17_reg_485;
wire   [3:0] select_ln148_18_fu_194_p3;
wire   [1:0] select_ln148_16_fu_359_p3;
reg   [1:0] select_ln148_16_reg_497;
reg    ap_enable_reg_pp0_iter1;
wire   [4:0] p_fu_445_p2;
reg   [4:0] p_reg_512;
reg   [4:0] p_reg_512_pp0_iter2_reg;
reg   [4:0] p_reg_512_pp0_iter3_reg;
reg   [4:0] p_reg_512_pp0_iter4_reg;
wire   [1:0] add_ln149_fu_451_p2;
reg    ap_block_state1;
wire    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_flush_enable;
reg    ap_enable_reg_pp0_iter2;
reg    ap_condition_pp0_exit_iter1_state3;
reg    ap_enable_reg_pp0_iter3;
reg    ap_enable_reg_pp0_iter4;
reg    ap_enable_reg_pp0_iter5;
reg   [1:0] ap_phi_mux_ii_phi_fu_108_p4;
wire    ap_block_pp0_stage0;
reg   [1:0] ap_phi_mux_jj_phi_fu_131_p4;
wire   [63:0] p_cast27_fu_439_p1;
wire   [63:0] idxprom30_fu_457_p1;
wire   [15:0] grp_fu_149_p2;
wire   [3:0] add_ln148_6_fu_188_p2;
wire   [3:0] shl_ln_fu_206_p3;
wire   [4:0] zext_ln150_7_fu_214_p1;
wire   [4:0] zext_ln150_fu_202_p1;
wire   [4:0] sub_ln150_fu_218_p2;
wire   [4:0] zext_ln150_8_fu_224_p1;
wire   [4:0] add_ln150_fu_228_p2;
wire   [4:0] shl_ln150_fu_234_p2;
wire   [3:0] tmp_s_fu_256_p3;
wire   [4:0] tmp_145_cast_fu_263_p1;
wire   [4:0] select_ln147_22_cast_fu_253_p1;
wire   [4:0] empty_122_fu_267_p2;
wire   [3:0] shl_ln150_mid1_fu_280_p3;
wire   [4:0] zext_ln150_13_fu_287_p1;
wire   [4:0] zext_ln150_12_fu_277_p1;
wire   [4:0] sub_ln150_6_fu_291_p2;
wire   [4:0] shl_ln150_1_fu_304_p2;
wire   [4:0] sub_ln150_7_fu_310_p2;
wire   [4:0] sub_ln150_1_fu_240_p2;
wire   [0:0] icmp_ln149_fu_328_p2;
wire   [0:0] xor_ln147_fu_323_p2;
wire   [1:0] select_ln147_fu_246_p3;
wire   [0:0] and_ln147_fu_334_p2;
wire   [0:0] or_ln148_fu_346_p2;
wire   [1:0] add_ln148_fu_340_p2;
wire   [5:0] sext_ln150_fu_273_p1;
wire   [5:0] select_ln148_21_cast_fu_367_p1;
wire   [5:0] empty_123_fu_371_p2;
wire   [2:0] empty_125_fu_381_p1;
wire   [4:0] p_shl_cast_fu_385_p3;
wire   [4:0] empty_124_fu_377_p1;
wire   [4:0] select_ln147_18_fu_297_p3;
wire   [4:0] zext_ln150_14_fu_399_p1;
wire   [4:0] add_ln150_6_fu_403_p2;
wire   [4:0] shl_ln150_2_fu_409_p2;
wire   [4:0] sub_ln150_8_fu_415_p2;
wire   [4:0] select_ln147_19_fu_316_p3;
wire   [1:0] select_ln148_fu_351_p3;
wire   [4:0] empty_126_fu_393_p2;
wire   [4:0] select_ln148_cast_fu_429_p1;
wire   [4:0] empty_127_fu_433_p2;
wire   [4:0] select_ln148_17_fu_421_p3;
wire    ap_CS_fsm_state8;
reg   [2:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
#0 ap_enable_reg_pp0_iter4 = 1'b0;
#0 ap_enable_reg_pp0_iter5 = 1'b0;
end

td_fused_top_hmul_16ns_16ns_16_4_max_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hmul_16ns_16ns_16_4_max_dsp_1_U20(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(ifmap_vec_q0),
    .din1(weight_vecs_0_q0),
    .dout(grp_fu_149_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if ((1'b1 == ap_condition_pp0_flush_enable)) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            if ((1'b1 == ap_condition_pp0_exit_iter1_state3)) begin
                ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter0;
            end else if ((1'b1 == 1'b1)) begin
                ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
            end
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter4 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter5 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter5 <= ap_enable_reg_pp0_iter4;
        end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter5 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln147_reg_466 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ic_reg_138 <= add_ln149_fu_451_p2;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ic_reg_138 <= 2'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln147_reg_466 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ii_reg_104 <= select_ln147_17_reg_485;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ii_reg_104 <= 2'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_fu_162_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        indvar_flatten21_reg_93 <= add_ln147_6_fu_156_p2;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indvar_flatten21_reg_93 <= 5'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_fu_162_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        indvar_flatten_reg_116 <= select_ln148_18_fu_194_p3;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indvar_flatten_reg_116 <= 4'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_reg_466_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        jj_reg_127 <= select_ln148_16_reg_497;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        jj_reg_127 <= 2'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_fu_162_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        add_ln147_reg_470 <= add_ln147_fu_168_p2;
        icmp_ln148_reg_476 <= icmp_ln148_fu_174_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln147_reg_466 <= icmp_ln147_fu_162_p2;
        icmp_ln147_reg_466_pp0_iter1_reg <= icmp_ln147_reg_466;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        icmp_ln147_reg_466_pp0_iter2_reg <= icmp_ln147_reg_466_pp0_iter1_reg;
        icmp_ln147_reg_466_pp0_iter3_reg <= icmp_ln147_reg_466_pp0_iter2_reg;
        icmp_ln147_reg_466_pp0_iter4_reg <= icmp_ln147_reg_466_pp0_iter3_reg;
        p_reg_512_pp0_iter2_reg <= p_reg_512;
        p_reg_512_pp0_iter3_reg <= p_reg_512_pp0_iter2_reg;
        p_reg_512_pp0_iter4_reg <= p_reg_512_pp0_iter3_reg;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_reg_466 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        p_reg_512 <= p_fu_445_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_fu_162_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        select_ln147_17_reg_485 <= select_ln147_17_fu_180_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln147_reg_466 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        select_ln148_16_reg_497 <= select_ln148_16_fu_359_p3;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_condition_pp0_exit_iter1_state3 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter1_state3 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln147_fu_162_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_condition_pp0_flush_enable = 1'b1;
    end else begin
        ap_condition_pp0_flush_enable = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state8)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln147_reg_466 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_phi_mux_ii_phi_fu_108_p4 = select_ln147_17_reg_485;
    end else begin
        ap_phi_mux_ii_phi_fu_108_p4 = ii_reg_104;
    end
end

always @ (*) begin
    if (((icmp_ln147_reg_466_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        ap_phi_mux_jj_phi_fu_131_p4 = select_ln148_16_reg_497;
    end else begin
        ap_phi_mux_jj_phi_fu_131_p4 = jj_reg_127;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state8)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ifmap_vec_ce0 = 1'b1;
    end else begin
        ifmap_vec_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter5 == 1'b1))) begin
        products_0_ce0 = 1'b1;
    end else begin
        products_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln147_reg_466_pp0_iter4_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter5 == 1'b1))) begin
        products_0_we0 = 1'b1;
    end else begin
        products_0_we0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        weight_vecs_0_ce0 = 1'b1;
    end else begin
        weight_vecs_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((~((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b0)) & ~((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter5 == 1'b1) & (ap_enable_reg_pp0_iter4 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if ((((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b0)) | ((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter5 == 1'b1) & (ap_enable_reg_pp0_iter4 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_state8;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state8 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln147_6_fu_156_p2 = (indvar_flatten21_reg_93 + 5'd1);

assign add_ln147_fu_168_p2 = (ap_phi_mux_ii_phi_fu_108_p4 + 2'd1);

assign add_ln148_6_fu_188_p2 = (indvar_flatten_reg_116 + 4'd1);

assign add_ln148_fu_340_p2 = (select_ln147_fu_246_p3 + 2'd1);

assign add_ln149_fu_451_p2 = (select_ln148_fu_351_p3 + 2'd1);

assign add_ln150_6_fu_403_p2 = (select_ln147_18_fu_297_p3 + zext_ln150_14_fu_399_p1);

assign add_ln150_fu_228_p2 = (sub_ln150_fu_218_p2 + zext_ln150_8_fu_224_p1);

assign and_ln147_fu_334_p2 = (xor_ln147_fu_323_p2 & icmp_ln149_fu_328_p2);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state8 = ap_CS_fsm[32'd2];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (ap_done_reg == 1'b1));
end

assign ap_block_state2_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter4 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage0_iter5 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign empty_122_fu_267_p2 = (tmp_145_cast_fu_263_p1 - select_ln147_22_cast_fu_253_p1);

assign empty_123_fu_371_p2 = ((sext_ln150_fu_273_p1) + (select_ln148_21_cast_fu_367_p1));

assign empty_124_fu_377_p1 = empty_123_fu_371_p2[4:0];

assign empty_125_fu_381_p1 = empty_123_fu_371_p2[2:0];

assign empty_126_fu_393_p2 = (p_shl_cast_fu_385_p3 - empty_124_fu_377_p1);

assign empty_127_fu_433_p2 = (empty_126_fu_393_p2 + select_ln148_cast_fu_429_p1);

assign icmp_ln147_fu_162_p2 = ((indvar_flatten21_reg_93 == 5'd27) ? 1'b1 : 1'b0);

assign icmp_ln148_fu_174_p2 = ((indvar_flatten_reg_116 == 4'd9) ? 1'b1 : 1'b0);

assign icmp_ln149_fu_328_p2 = ((ic_reg_138 == 2'd3) ? 1'b1 : 1'b0);

assign idxprom30_fu_457_p1 = p_reg_512_pp0_iter4_reg;

assign ifmap_vec_address0 = p_cast27_fu_439_p1;

assign or_ln148_fu_346_p2 = (icmp_ln148_reg_476 | and_ln147_fu_334_p2);

assign p_cast27_fu_439_p1 = empty_127_fu_433_p2;

assign p_fu_445_p2 = (select_ln148_17_fu_421_p3 + select_ln148_cast_fu_429_p1);

assign p_shl_cast_fu_385_p3 = {{empty_125_fu_381_p1}, {2'd0}};

assign products_0_address0 = idxprom30_fu_457_p1;

assign products_0_d0 = grp_fu_149_p2;

assign select_ln147_17_fu_180_p3 = ((icmp_ln148_fu_174_p2[0:0] == 1'b1) ? add_ln147_fu_168_p2 : ap_phi_mux_ii_phi_fu_108_p4);

assign select_ln147_18_fu_297_p3 = ((icmp_ln148_reg_476[0:0] == 1'b1) ? sub_ln150_6_fu_291_p2 : sub_ln150_fu_218_p2);

assign select_ln147_19_fu_316_p3 = ((icmp_ln148_reg_476[0:0] == 1'b1) ? sub_ln150_7_fu_310_p2 : sub_ln150_1_fu_240_p2);

assign select_ln147_22_cast_fu_253_p1 = select_ln147_17_reg_485;

assign select_ln147_fu_246_p3 = ((icmp_ln148_reg_476[0:0] == 1'b1) ? 2'd0 : ap_phi_mux_jj_phi_fu_131_p4);

assign select_ln148_16_fu_359_p3 = ((and_ln147_fu_334_p2[0:0] == 1'b1) ? add_ln148_fu_340_p2 : select_ln147_fu_246_p3);

assign select_ln148_17_fu_421_p3 = ((and_ln147_fu_334_p2[0:0] == 1'b1) ? sub_ln150_8_fu_415_p2 : select_ln147_19_fu_316_p3);

assign select_ln148_18_fu_194_p3 = ((icmp_ln148_fu_174_p2[0:0] == 1'b1) ? 4'd1 : add_ln148_6_fu_188_p2);

assign select_ln148_21_cast_fu_367_p1 = select_ln148_16_fu_359_p3;

assign select_ln148_cast_fu_429_p1 = select_ln148_fu_351_p3;

assign select_ln148_fu_351_p3 = ((or_ln148_fu_346_p2[0:0] == 1'b1) ? 2'd0 : ic_reg_138);

assign sext_ln150_fu_273_p1 = (empty_122_fu_267_p2);

assign shl_ln150_1_fu_304_p2 = sub_ln150_6_fu_291_p2 << 5'd2;

assign shl_ln150_2_fu_409_p2 = add_ln150_6_fu_403_p2 << 5'd2;

assign shl_ln150_fu_234_p2 = add_ln150_fu_228_p2 << 5'd2;

assign shl_ln150_mid1_fu_280_p3 = {{add_ln147_reg_470}, {2'd0}};

assign shl_ln_fu_206_p3 = {{ii_reg_104}, {2'd0}};

assign sub_ln150_1_fu_240_p2 = (shl_ln150_fu_234_p2 - add_ln150_fu_228_p2);

assign sub_ln150_6_fu_291_p2 = (zext_ln150_13_fu_287_p1 - zext_ln150_12_fu_277_p1);

assign sub_ln150_7_fu_310_p2 = (shl_ln150_1_fu_304_p2 - sub_ln150_6_fu_291_p2);

assign sub_ln150_8_fu_415_p2 = (shl_ln150_2_fu_409_p2 - add_ln150_6_fu_403_p2);

assign sub_ln150_fu_218_p2 = (zext_ln150_7_fu_214_p1 - zext_ln150_fu_202_p1);

assign tmp_145_cast_fu_263_p1 = tmp_s_fu_256_p3;

assign tmp_s_fu_256_p3 = {{select_ln147_17_reg_485}, {2'd0}};

assign weight_vecs_0_address0 = p_cast27_fu_439_p1;

assign xor_ln147_fu_323_p2 = (icmp_ln148_reg_476 ^ 1'd1);

assign zext_ln150_12_fu_277_p1 = add_ln147_reg_470;

assign zext_ln150_13_fu_287_p1 = shl_ln150_mid1_fu_280_p3;

assign zext_ln150_14_fu_399_p1 = add_ln148_fu_340_p2;

assign zext_ln150_7_fu_214_p1 = shl_ln_fu_206_p3;

assign zext_ln150_8_fu_224_p1 = ap_phi_mux_jj_phi_fu_131_p4;

assign zext_ln150_fu_202_p1 = ii_reg_104;

endmodule //td_fused_top_tdf1_dot_product
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_tdf1_filters_ram (addr0, ce0, q0, addr1, ce1, d1, we1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 9;
parameter MEM_SIZE = 432;

input[AWIDTH-1:0] addr0;
input ce0;
output wire[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
input clk;

 reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];
wire [AWIDTH-1:0] addr0_t0; 
reg [AWIDTH-1:0] addr0_t1; 
reg [DWIDTH-1:0] q0_t0;
reg [DWIDTH-1:0] q0_t1;
wire [AWIDTH-1:0] addr1_t0; 
reg [AWIDTH-1:0] addr1_t1; 
wire [DWIDTH-1:0] d1_t0; 
wire we1_t0; 
reg [DWIDTH-1:0] d1_t1; 
reg we1_t1; 


assign addr0_t0 = addr0;
assign q0 = q0_t1;
assign addr1_t0 = addr1;
assign d1_t0 = d1;
assign we1_t0 = we1;

always @(posedge clk)  
begin
    if (ce0) 
    begin
        addr0_t1 <= addr0_t0; 
        q0_t1 <= q0_t0;
    end
    if (ce1) 
    begin
        addr1_t1 <= addr1_t0; 
        d1_t1 <= d1_t0;
        we1_t1 <= we1_t0;
    end
end


always @(posedge clk)  
begin 
    if (ce0) begin
        q0_t0 <= ram[addr0_t1];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1_t1) 
            ram[addr1_t1] <= d1_t1; 
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_tdf1_filters(
    reset,
    clk,
    address0,
    ce0,
    q0,
    address1,
    ce1,
    we1,
    d1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd432;
parameter AddressWidth = 32'd9;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;



td_fused_top_tdf1_filters_ram td_fused_top_tdf1_filters_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 )
);

endmodule

// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf1_get_next_ijk (
        ap_clk,
        ap_rst,
        ap_start,
        start_full_n,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        start_out,
        start_write,
        input_indices_2_out_din,
        input_indices_2_out_full_n,
        input_indices_2_out_write,
        input_indices_2_out1_din,
        input_indices_2_out1_full_n,
        input_indices_2_out1_write,
        output_indices_0_din,
        output_indices_0_full_n,
        output_indices_0_write,
        output_indices_1_din,
        output_indices_1_full_n,
        output_indices_1_write,
        resetMaximum_din,
        resetMaximum_full_n,
        resetMaximum_write,
        storeOutput_din,
        storeOutput_full_n,
        storeOutput_write,
        ap_return_0,
        ap_return_1
);

parameter    ap_ST_fsm_state1 = 1'd1;

input   ap_clk;
input   ap_rst;
input   ap_start;
input   start_full_n;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output   start_out;
output   start_write;
output  [3:0] input_indices_2_out_din;
input   input_indices_2_out_full_n;
output   input_indices_2_out_write;
output  [3:0] input_indices_2_out1_din;
input   input_indices_2_out1_full_n;
output   input_indices_2_out1_write;
output  [6:0] output_indices_0_din;
input   output_indices_0_full_n;
output   output_indices_0_write;
output  [13:0] output_indices_1_din;
input   output_indices_1_full_n;
output   output_indices_1_write;
output   resetMaximum_din;
input   resetMaximum_full_n;
output   resetMaximum_write;
output   storeOutput_din;
input   storeOutput_full_n;
output   storeOutput_write;
output  [15:0] ap_return_0;
output  [15:0] ap_return_1;

reg ap_done;
reg ap_idle;
reg start_write;
reg input_indices_2_out_write;
reg input_indices_2_out1_write;
reg output_indices_0_write;
reg output_indices_1_write;
reg resetMaximum_write;
reg storeOutput_write;

reg    real_start;
reg    start_once_reg;
reg    ap_done_reg;
  reg   [0:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    internal_ap_ready;
reg   [1:0] i_p_3;
reg   [1:0] j_p_3;
reg   [15:0] i_7;
reg   [15:0] j_7;
reg   [15:0] k_7;
reg   [15:0] i_out_3;
reg   [15:0] j_out_3;
reg    input_indices_2_out_blk_n;
reg    input_indices_2_out1_blk_n;
reg    output_indices_0_blk_n;
reg    output_indices_1_blk_n;
reg    resetMaximum_blk_n;
reg    storeOutput_blk_n;
wire   [1:0] select_ln163_fu_338_p3;
reg    ap_block_state1;
wire   [0:0] or_ln163_fu_312_p2;
wire   [1:0] select_ln163_1_fu_346_p3;
wire   [15:0] select_ln168_fu_278_p3;
wire   [0:0] and_ln163_1_fu_306_p2;
wire   [15:0] select_ln163_2_fu_360_p3;
wire   [0:0] and_ln153_fu_354_p2;
wire   [15:0] select_ln163_3_fu_388_p3;
wire   [0:0] and_ln156_fu_294_p2;
wire   [15:0] select_ln168_1_fu_286_p3;
wire   [15:0] select_ln163_4_fu_396_p3;
wire   [3:0] trunc_ln149_fu_182_p1;
wire   [1:0] or_ln145_fu_126_p2;
wire   [0:0] icmp_ln146_fu_139_p2;
wire   [0:0] icmp_ln146_1_fu_145_p2;
wire   [15:0] zext_ln147_fu_114_p1;
wire   [15:0] zext_ln148_fu_122_p1;
wire   [1:0] add_ln152_fu_206_p2;
wire   [1:0] add_ln155_fu_218_p2;
wire   [15:0] add_ln158_fu_230_p2;
wire   [15:0] add_ln162_fu_248_p2;
wire   [15:0] add_ln167_fu_266_p2;
wire   [0:0] icmp_ln168_fu_272_p2;
wire   [15:0] add_ln166_fu_260_p2;
wire   [0:0] icmp_ln153_fu_212_p2;
wire   [0:0] icmp_ln156_fu_224_p2;
wire   [0:0] icmp_ln159_fu_236_p2;
wire   [0:0] icmp_ln163_fu_254_p2;
wire   [0:0] and_ln163_fu_300_p2;
wire   [0:0] xor_ln156_fu_318_p2;
wire   [0:0] and_ln156_1_fu_324_p2;
wire   [1:0] select_ln156_fu_330_p3;
wire   [15:0] add_ln161_fu_242_p2;
wire   [0:0] xor_ln159_fu_368_p2;
wire   [0:0] and_ln159_fu_374_p2;
wire   [15:0] select_ln159_fu_380_p3;
wire   [15:0] add_ln147_fu_162_p2;
wire   [15:0] add_ln148_fu_172_p2;
reg   [0:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 start_once_reg = 1'b0;
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 1'd1;
#0 i_p_3 = 2'd0;
#0 j_p_3 = 2'd0;
#0 i_7 = 16'd0;
#0 j_7 = 16'd0;
#0 k_7 = 16'd0;
#0 i_out_3 = 16'd0;
#0 j_out_3 = 16'd0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        start_once_reg <= 1'b0;
    end else begin
        if (((real_start == 1'b1) & (internal_ap_ready == 1'b0))) begin
            start_once_reg <= 1'b1;
        end else if ((internal_ap_ready == 1'b1)) begin
            start_once_reg <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1) & (1'd1 == and_ln163_1_fu_306_p2))) begin
        i_7 <= select_ln168_fu_278_p3;
        i_out_3 <= select_ln168_1_fu_286_p3;
    end
end

always @ (posedge ap_clk) begin
    if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (or_ln163_fu_312_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1))) begin
        i_p_3 <= select_ln163_fu_338_p3;
    end
end

always @ (posedge ap_clk) begin
    if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1) & (1'd1 == and_ln153_fu_354_p2))) begin
        j_7 <= select_ln163_2_fu_360_p3;
        j_out_3 <= select_ln163_4_fu_396_p3;
    end
end

always @ (posedge ap_clk) begin
    if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        j_p_3 <= select_ln163_1_fu_346_p3;
    end
end

always @ (posedge ap_clk) begin
    if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1) & (1'd1 == and_ln156_fu_294_p2))) begin
        k_7 <= select_ln163_3_fu_388_p3;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((real_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        input_indices_2_out1_blk_n = input_indices_2_out1_full_n;
    end else begin
        input_indices_2_out1_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        input_indices_2_out1_write = 1'b1;
    end else begin
        input_indices_2_out1_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        input_indices_2_out_blk_n = input_indices_2_out_full_n;
    end else begin
        input_indices_2_out_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        input_indices_2_out_write = 1'b1;
    end else begin
        input_indices_2_out_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        internal_ap_ready = 1'b1;
    end else begin
        internal_ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        output_indices_0_blk_n = output_indices_0_full_n;
    end else begin
        output_indices_0_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        output_indices_0_write = 1'b1;
    end else begin
        output_indices_0_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        output_indices_1_blk_n = output_indices_1_full_n;
    end else begin
        output_indices_1_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        output_indices_1_write = 1'b1;
    end else begin
        output_indices_1_write = 1'b0;
    end
end

always @ (*) begin
    if (((start_full_n == 1'b0) & (start_once_reg == 1'b0))) begin
        real_start = 1'b0;
    end else begin
        real_start = ap_start;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        resetMaximum_blk_n = resetMaximum_full_n;
    end else begin
        resetMaximum_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        resetMaximum_write = 1'b1;
    end else begin
        resetMaximum_write = 1'b0;
    end
end

always @ (*) begin
    if (((real_start == 1'b1) & (start_once_reg == 1'b0))) begin
        start_write = 1'b1;
    end else begin
        start_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        storeOutput_blk_n = storeOutput_full_n;
    end else begin
        storeOutput_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        storeOutput_write = 1'b1;
    end else begin
        storeOutput_write = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln147_fu_162_p2 = (i_7 + zext_ln147_fu_114_p1);

assign add_ln148_fu_172_p2 = (j_7 + zext_ln148_fu_122_p1);

assign add_ln152_fu_206_p2 = (j_p_3 + 2'd1);

assign add_ln155_fu_218_p2 = (i_p_3 + 2'd1);

assign add_ln158_fu_230_p2 = (k_7 + 16'd1);

assign add_ln161_fu_242_p2 = (j_7 + 16'd2);

assign add_ln162_fu_248_p2 = (j_out_3 + 16'd1);

assign add_ln166_fu_260_p2 = (i_7 + 16'd2);

assign add_ln167_fu_266_p2 = (i_out_3 + 16'd1);

assign and_ln153_fu_354_p2 = (icmp_ln159_fu_236_p2 & and_ln156_fu_294_p2);

assign and_ln156_1_fu_324_p2 = (xor_ln156_fu_318_p2 & icmp_ln153_fu_212_p2);

assign and_ln156_fu_294_p2 = (icmp_ln156_fu_224_p2 & icmp_ln153_fu_212_p2);

assign and_ln159_fu_374_p2 = (xor_ln159_fu_368_p2 & and_ln156_fu_294_p2);

assign and_ln163_1_fu_306_p2 = (and_ln163_fu_300_p2 & and_ln156_fu_294_p2);

assign and_ln163_fu_300_p2 = (icmp_ln163_fu_254_p2 & icmp_ln159_fu_236_p2);

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

always @ (*) begin
    ap_block_state1 = ((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1));
end

assign ap_ready = internal_ap_ready;

assign ap_return_0 = add_ln147_fu_162_p2;

assign ap_return_1 = add_ln148_fu_172_p2;

assign icmp_ln146_1_fu_145_p2 = ((j_p_3 == 2'd1) ? 1'b1 : 1'b0);

assign icmp_ln146_fu_139_p2 = ((i_p_3 == 2'd1) ? 1'b1 : 1'b0);

assign icmp_ln153_fu_212_p2 = ((add_ln152_fu_206_p2 == 2'd2) ? 1'b1 : 1'b0);

assign icmp_ln156_fu_224_p2 = ((add_ln155_fu_218_p2 == 2'd2) ? 1'b1 : 1'b0);

assign icmp_ln159_fu_236_p2 = ((add_ln158_fu_230_p2 == 16'd16) ? 1'b1 : 1'b0);

assign icmp_ln163_fu_254_p2 = ((add_ln162_fu_248_p2 == 16'd112) ? 1'b1 : 1'b0);

assign icmp_ln168_fu_272_p2 = ((add_ln167_fu_266_p2 == 16'd112) ? 1'b1 : 1'b0);

assign input_indices_2_out1_din = trunc_ln149_fu_182_p1;

assign input_indices_2_out_din = trunc_ln149_fu_182_p1;

assign or_ln145_fu_126_p2 = (j_p_3 | i_p_3);

assign or_ln163_fu_312_p2 = (icmp_ln153_fu_212_p2 | and_ln163_1_fu_306_p2);

assign output_indices_0_din = i_out_3[6:0];

assign output_indices_1_din = j_out_3[13:0];

assign resetMaximum_din = ((or_ln145_fu_126_p2 == 2'd0) ? 1'b1 : 1'b0);

assign select_ln156_fu_330_p3 = ((and_ln156_1_fu_324_p2[0:0] == 1'b1) ? add_ln155_fu_218_p2 : 2'd0);

assign select_ln159_fu_380_p3 = ((and_ln159_fu_374_p2[0:0] == 1'b1) ? add_ln158_fu_230_p2 : 16'd0);

assign select_ln163_1_fu_346_p3 = ((or_ln163_fu_312_p2[0:0] == 1'b1) ? 2'd0 : add_ln152_fu_206_p2);

assign select_ln163_2_fu_360_p3 = ((and_ln163_1_fu_306_p2[0:0] == 1'b1) ? 16'd0 : add_ln161_fu_242_p2);

assign select_ln163_3_fu_388_p3 = ((and_ln163_1_fu_306_p2[0:0] == 1'b1) ? 16'd0 : select_ln159_fu_380_p3);

assign select_ln163_4_fu_396_p3 = ((and_ln163_1_fu_306_p2[0:0] == 1'b1) ? 16'd0 : add_ln162_fu_248_p2);

assign select_ln163_fu_338_p3 = ((and_ln163_1_fu_306_p2[0:0] == 1'b1) ? 2'd0 : select_ln156_fu_330_p3);

assign select_ln168_1_fu_286_p3 = ((icmp_ln168_fu_272_p2[0:0] == 1'b1) ? 16'd0 : add_ln167_fu_266_p2);

assign select_ln168_fu_278_p3 = ((icmp_ln168_fu_272_p2[0:0] == 1'b1) ? 16'd0 : add_ln166_fu_260_p2);

assign start_out = real_start;

assign storeOutput_din = (icmp_ln146_fu_139_p2 & icmp_ln146_1_fu_145_p2);

assign trunc_ln149_fu_182_p1 = k_7[3:0];

assign xor_ln156_fu_318_p2 = (icmp_ln156_fu_224_p2 ^ 1'd1);

assign xor_ln159_fu_368_p2 = (icmp_ln159_fu_236_p2 ^ 1'd1);

assign zext_ln147_fu_114_p1 = i_p_3;

assign zext_ln148_fu_122_p1 = j_p_3;

endmodule //td_fused_top_tdf1_get_next_ijk
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf1_poolOutputs (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        output_indices_04_dout,
        output_indices_04_empty_n,
        output_indices_04_read,
        output_indices_15_dout,
        output_indices_15_empty_n,
        output_indices_15_read,
        resetMaximum6_dout,
        resetMaximum6_empty_n,
        resetMaximum6_read,
        storeOutput7_dout,
        storeOutput7_empty_n,
        storeOutput7_read,
        p_read,
        out_data_address1,
        out_data_ce1,
        out_data_we1,
        out_data_d1
);

parameter    ap_ST_fsm_state1 = 4'd1;
parameter    ap_ST_fsm_state2 = 4'd2;
parameter    ap_ST_fsm_state3 = 4'd4;
parameter    ap_ST_fsm_state4 = 4'd8;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
input  [6:0] output_indices_04_dout;
input   output_indices_04_empty_n;
output   output_indices_04_read;
input  [13:0] output_indices_15_dout;
input   output_indices_15_empty_n;
output   output_indices_15_read;
input  [0:0] resetMaximum6_dout;
input   resetMaximum6_empty_n;
output   resetMaximum6_read;
input  [0:0] storeOutput7_dout;
input   storeOutput7_empty_n;
output   storeOutput7_read;
input  [15:0] p_read;
output  [15:0] out_data_address1;
output   out_data_ce1;
output   out_data_we1;
output  [63:0] out_data_d1;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg output_indices_04_read;
reg output_indices_15_read;
reg resetMaximum6_read;
reg storeOutput7_read;

reg    ap_done_reg;
  reg   [3:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg   [15:0] max_vals_3_0;
reg    output_indices_04_blk_n;
wire    ap_CS_fsm_state2;
reg    output_indices_15_blk_n;
reg    resetMaximum6_blk_n;
reg    storeOutput7_blk_n;
reg   [6:0] output_indices_04_read_reg_147;
reg   [13:0] output_indices_15_read_reg_152;
wire   [0:0] storeOutput7_read_read_fu_82_p2;
reg   [0:0] storeOutput7_read_reg_157;
wire    grp_tdf1_writeOutputs_unaligned_fu_88_ap_start;
wire    grp_tdf1_writeOutputs_unaligned_fu_88_ap_done;
wire    grp_tdf1_writeOutputs_unaligned_fu_88_ap_idle;
wire    grp_tdf1_writeOutputs_unaligned_fu_88_ap_ready;
wire   [15:0] grp_tdf1_writeOutputs_unaligned_fu_88_out_data_address1;
wire    grp_tdf1_writeOutputs_unaligned_fu_88_out_data_ce1;
wire    grp_tdf1_writeOutputs_unaligned_fu_88_out_data_we1;
wire   [63:0] grp_tdf1_writeOutputs_unaligned_fu_88_out_data_d1;
reg    grp_tdf1_writeOutputs_unaligned_fu_88_ap_start_reg;
wire    ap_CS_fsm_state3;
wire    ap_CS_fsm_state4;
reg    ap_block_state4_on_subcall_done;
wire   [15:0] select_ln24_fu_126_p3;
reg    ap_block_state2;
reg    ap_block_state1;
wire   [0:0] grp_fu_110_p2;
wire   [0:0] or_ln24_fu_120_p2;
reg    grp_fu_110_ce;
reg   [3:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 4'd1;
#0 max_vals_3_0 = 16'd0;
#0 grp_tdf1_writeOutputs_unaligned_fu_88_ap_start_reg = 1'b0;
end

td_fused_top_tdf1_writeOutputs_unaligned grp_tdf1_writeOutputs_unaligned_fu_88(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(grp_tdf1_writeOutputs_unaligned_fu_88_ap_start),
    .ap_done(grp_tdf1_writeOutputs_unaligned_fu_88_ap_done),
    .ap_idle(grp_tdf1_writeOutputs_unaligned_fu_88_ap_idle),
    .ap_ready(grp_tdf1_writeOutputs_unaligned_fu_88_ap_ready),
    .i(output_indices_04_read_reg_147),
    .j(output_indices_15_read_reg_152),
    .out_data_address1(grp_tdf1_writeOutputs_unaligned_fu_88_out_data_address1),
    .out_data_ce1(grp_tdf1_writeOutputs_unaligned_fu_88_out_data_ce1),
    .out_data_we1(grp_tdf1_writeOutputs_unaligned_fu_88_out_data_we1),
    .out_data_d1(grp_tdf1_writeOutputs_unaligned_fu_88_out_data_d1),
    .max_vals_3_0(max_vals_3_0)
);

td_fused_top_hcmp_16ns_16ns_1_2_no_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 1 ))
hcmp_16ns_16ns_1_2_no_dsp_1_U47(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(grp_fu_110_ce),
    .din0(max_vals_3_0),
    .din1(p_read),
    .opcode(5'd4),
    .dout(grp_fu_110_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_state4) & (1'b0 == ap_block_state4_on_subcall_done))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        grp_tdf1_writeOutputs_unaligned_fu_88_ap_start_reg <= 1'b0;
    end else begin
        if ((1'b1 == ap_CS_fsm_state3)) begin
            grp_tdf1_writeOutputs_unaligned_fu_88_ap_start_reg <= 1'b1;
        end else if ((grp_tdf1_writeOutputs_unaligned_fu_88_ap_ready == 1'b1)) begin
            grp_tdf1_writeOutputs_unaligned_fu_88_ap_start_reg <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((~((storeOutput7_empty_n == 1'b0) | (resetMaximum6_empty_n == 1'b0) | (output_indices_15_empty_n == 1'b0) | (output_indices_04_empty_n == 1'b0)) & (1'b1 == ap_CS_fsm_state2))) begin
        max_vals_3_0 <= select_ln24_fu_126_p3;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        output_indices_04_read_reg_147 <= output_indices_04_dout;
        output_indices_15_read_reg_152 <= output_indices_15_dout;
        storeOutput7_read_reg_157 <= storeOutput7_dout;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state4) & (1'b0 == ap_block_state4_on_subcall_done))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state4) & (1'b0 == ap_block_state4_on_subcall_done))) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1)) | (~((storeOutput7_empty_n == 1'b0) | (resetMaximum6_empty_n == 1'b0) | (output_indices_15_empty_n == 1'b0) | (output_indices_04_empty_n == 1'b0)) & (1'b1 == ap_CS_fsm_state2)))) begin
        grp_fu_110_ce = 1'b1;
    end else begin
        grp_fu_110_ce = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        output_indices_04_blk_n = output_indices_04_empty_n;
    end else begin
        output_indices_04_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((storeOutput7_empty_n == 1'b0) | (resetMaximum6_empty_n == 1'b0) | (output_indices_15_empty_n == 1'b0) | (output_indices_04_empty_n == 1'b0)) & (1'b1 == ap_CS_fsm_state2))) begin
        output_indices_04_read = 1'b1;
    end else begin
        output_indices_04_read = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        output_indices_15_blk_n = output_indices_15_empty_n;
    end else begin
        output_indices_15_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((storeOutput7_empty_n == 1'b0) | (resetMaximum6_empty_n == 1'b0) | (output_indices_15_empty_n == 1'b0) | (output_indices_04_empty_n == 1'b0)) & (1'b1 == ap_CS_fsm_state2))) begin
        output_indices_15_read = 1'b1;
    end else begin
        output_indices_15_read = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        resetMaximum6_blk_n = resetMaximum6_empty_n;
    end else begin
        resetMaximum6_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((storeOutput7_empty_n == 1'b0) | (resetMaximum6_empty_n == 1'b0) | (output_indices_15_empty_n == 1'b0) | (output_indices_04_empty_n == 1'b0)) & (1'b1 == ap_CS_fsm_state2))) begin
        resetMaximum6_read = 1'b1;
    end else begin
        resetMaximum6_read = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        storeOutput7_blk_n = storeOutput7_empty_n;
    end else begin
        storeOutput7_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((storeOutput7_empty_n == 1'b0) | (resetMaximum6_empty_n == 1'b0) | (output_indices_15_empty_n == 1'b0) | (output_indices_04_empty_n == 1'b0)) & (1'b1 == ap_CS_fsm_state2))) begin
        storeOutput7_read = 1'b1;
    end else begin
        storeOutput7_read = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_state2 : begin
            if ((~((storeOutput7_empty_n == 1'b0) | (resetMaximum6_empty_n == 1'b0) | (output_indices_15_empty_n == 1'b0) | (output_indices_04_empty_n == 1'b0)) & (storeOutput7_read_read_fu_82_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state2))) begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end else if ((~((storeOutput7_empty_n == 1'b0) | (resetMaximum6_empty_n == 1'b0) | (output_indices_15_empty_n == 1'b0) | (output_indices_04_empty_n == 1'b0)) & (storeOutput7_read_read_fu_82_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end
        end
        ap_ST_fsm_state3 : begin
            ap_NS_fsm = ap_ST_fsm_state4;
        end
        ap_ST_fsm_state4 : begin
            if (((1'b1 == ap_CS_fsm_state4) & (1'b0 == ap_block_state4_on_subcall_done))) begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (ap_done_reg == 1'b1));
end

always @ (*) begin
    ap_block_state2 = ((storeOutput7_empty_n == 1'b0) | (resetMaximum6_empty_n == 1'b0) | (output_indices_15_empty_n == 1'b0) | (output_indices_04_empty_n == 1'b0));
end

always @ (*) begin
    ap_block_state4_on_subcall_done = ((grp_tdf1_writeOutputs_unaligned_fu_88_ap_done == 1'b0) & (storeOutput7_read_reg_157 == 1'd1));
end

assign grp_tdf1_writeOutputs_unaligned_fu_88_ap_start = grp_tdf1_writeOutputs_unaligned_fu_88_ap_start_reg;

assign or_ln24_fu_120_p2 = (resetMaximum6_dout | grp_fu_110_p2);

assign out_data_address1 = grp_tdf1_writeOutputs_unaligned_fu_88_out_data_address1;

assign out_data_ce1 = grp_tdf1_writeOutputs_unaligned_fu_88_out_data_ce1;

assign out_data_d1 = grp_tdf1_writeOutputs_unaligned_fu_88_out_data_d1;

assign out_data_we1 = grp_tdf1_writeOutputs_unaligned_fu_88_out_data_we1;

assign select_ln24_fu_126_p3 = ((or_ln24_fu_120_p2[0:0] == 1'b1) ? p_read : max_vals_3_0);

assign storeOutput7_read_read_fu_82_p2 = storeOutput7_dout;

endmodule //td_fused_top_tdf1_poolOutputs
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf1_readFilters18 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        filter_data_address0,
        filter_data_ce0,
        filter_data_q0,
        input_indices_23_dout,
        input_indices_23_empty_n,
        input_indices_23_read,
        weight_vecs_0_address0,
        weight_vecs_0_ce0,
        weight_vecs_0_we0,
        weight_vecs_0_d0
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state7 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [8:0] filter_data_address0;
output   filter_data_ce0;
input  [15:0] filter_data_q0;
input  [3:0] input_indices_23_dout;
input   input_indices_23_empty_n;
output   input_indices_23_read;
output  [4:0] weight_vecs_0_address0;
output   weight_vecs_0_ce0;
output   weight_vecs_0_we0;
output  [15:0] weight_vecs_0_d0;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg filter_data_ce0;
reg input_indices_23_read;
reg weight_vecs_0_ce0;
reg weight_vecs_0_we0;

reg    ap_done_reg;
  reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    input_indices_23_blk_n;
reg   [4:0] indvar_flatten13_reg_117;
reg   [1:0] ii_reg_128;
reg   [3:0] indvar_flatten_reg_139;
reg   [1:0] jj_reg_150;
reg   [1:0] kk_reg_161;
wire   [7:0] sext_ln47_fu_194_p1;
reg   [7:0] sext_ln47_reg_448;
wire   [4:0] add_ln47_6_fu_198_p2;
wire    ap_CS_fsm_pp0_stage0;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
wire    ap_block_state4_pp0_stage0_iter2;
wire    ap_block_state5_pp0_stage0_iter3;
wire    ap_block_state6_pp0_stage0_iter4;
wire    ap_block_pp0_stage0_11001;
wire   [0:0] icmp_ln47_fu_204_p2;
reg   [0:0] icmp_ln47_reg_458;
reg   [0:0] icmp_ln47_reg_458_pp0_iter1_reg;
reg   [0:0] icmp_ln47_reg_458_pp0_iter2_reg;
reg   [0:0] icmp_ln47_reg_458_pp0_iter3_reg;
wire   [0:0] icmp_ln48_fu_216_p2;
reg   [0:0] icmp_ln48_reg_462;
wire   [1:0] select_ln47_6_fu_222_p3;
reg   [1:0] select_ln47_6_reg_469;
wire   [3:0] select_ln48_12_fu_236_p3;
wire   [1:0] select_ln48_11_fu_341_p3;
reg   [1:0] select_ln48_11_reg_482;
reg    ap_enable_reg_pp0_iter1;
wire   [4:0] add_ln55_24_fu_432_p2;
reg   [4:0] add_ln55_24_reg_492;
reg   [4:0] add_ln55_24_reg_492_pp0_iter2_reg;
reg   [4:0] add_ln55_24_reg_492_pp0_iter3_reg;
wire   [1:0] add_ln49_fu_438_p2;
reg    ap_block_state1;
wire    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_flush_enable;
reg    ap_enable_reg_pp0_iter2;
reg    ap_condition_pp0_exit_iter1_state3;
reg    ap_enable_reg_pp0_iter3;
reg    ap_enable_reg_pp0_iter4;
reg   [1:0] ap_phi_mux_ii_phi_fu_132_p4;
wire    ap_block_pp0_stage0;
reg   [1:0] ap_phi_mux_jj_phi_fu_154_p4;
wire   [63:0] zext_ln55_57_fu_427_p1;
wire   [63:0] zext_ln55_58_fu_444_p1;
wire   [5:0] tmp_fu_176_p3;
wire   [6:0] zext_ln55_49_fu_184_p1;
wire   [6:0] zext_ln55_fu_172_p1;
wire   [6:0] sub_ln55_fu_188_p2;
wire   [1:0] add_ln47_fu_210_p2;
wire   [3:0] add_ln48_6_fu_230_p2;
wire   [7:0] zext_ln55_51_fu_254_p1;
wire   [7:0] add_ln55_fu_257_p2;
wire   [9:0] tmp_46_fu_266_p3;
wire   [61:0] sext_ln55_1_fu_274_p1;
wire   [61:0] sext_ln55_fu_262_p1;
wire   [3:0] tmp_s_fu_284_p3;
wire   [4:0] zext_ln55_52_fu_291_p1;
wire   [4:0] zext_ln55_50_fu_251_p1;
wire   [4:0] sub_ln55_12_fu_295_p2;
wire   [0:0] icmp_ln49_fu_310_p2;
wire   [0:0] xor_ln47_fu_305_p2;
wire   [1:0] select_ln47_fu_244_p3;
wire   [0:0] and_ln47_fu_316_p2;
wire   [0:0] or_ln48_fu_328_p2;
wire   [1:0] add_ln48_fu_322_p2;
wire   [61:0] sub_ln55_11_fu_278_p2;
wire   [61:0] zext_ln55_54_fu_353_p1;
wire   [61:0] add_ln55_21_fu_357_p2;
wire   [6:0] trunc_ln55_1_fu_367_p1;
wire   [8:0] p_shl2_cast_fu_371_p3;
wire   [8:0] trunc_ln55_fu_363_p1;
wire   [5:0] sext_ln48_fu_301_p1;
wire   [5:0] zext_ln55_53_fu_349_p1;
wire   [5:0] add_ln55_22_fu_385_p2;
wire   [2:0] trunc_ln55_3_fu_395_p1;
wire   [4:0] p_shl1_cast_fu_399_p3;
wire   [4:0] trunc_ln55_2_fu_391_p1;
wire   [1:0] select_ln48_fu_333_p3;
wire   [8:0] sub_ln55_13_fu_379_p2;
wire   [8:0] zext_ln55_56_fu_417_p1;
wire   [8:0] add_ln55_23_fu_421_p2;
wire   [4:0] sub_ln55_14_fu_407_p2;
wire   [4:0] zext_ln55_55_fu_413_p1;
wire    ap_CS_fsm_state7;
reg   [2:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
#0 ap_enable_reg_pp0_iter4 = 1'b0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state7)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if ((1'b1 == ap_condition_pp0_flush_enable)) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((~((ap_start == 1'b0) | (input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            if ((1'b1 == ap_condition_pp0_exit_iter1_state3)) begin
                ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter0;
            end else if ((1'b1 == 1'b1)) begin
                ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
            end
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter4 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
        end else if ((~((ap_start == 1'b0) | (input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter4 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln47_reg_458 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ii_reg_128 <= select_ln47_6_reg_469;
    end else if ((~((ap_start == 1'b0) | (input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ii_reg_128 <= 2'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_fu_204_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        indvar_flatten13_reg_117 <= add_ln47_6_fu_198_p2;
    end else if ((~((ap_start == 1'b0) | (input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indvar_flatten13_reg_117 <= 5'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_fu_204_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        indvar_flatten_reg_139 <= select_ln48_12_fu_236_p3;
    end else if ((~((ap_start == 1'b0) | (input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indvar_flatten_reg_139 <= 4'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_reg_458_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        jj_reg_150 <= select_ln48_11_reg_482;
    end else if ((~((ap_start == 1'b0) | (input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        jj_reg_150 <= 2'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln47_reg_458 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        kk_reg_161 <= add_ln49_fu_438_p2;
    end else if ((~((ap_start == 1'b0) | (input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        kk_reg_161 <= 2'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_reg_458 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        add_ln55_24_reg_492 <= add_ln55_24_fu_432_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        add_ln55_24_reg_492_pp0_iter2_reg <= add_ln55_24_reg_492;
        add_ln55_24_reg_492_pp0_iter3_reg <= add_ln55_24_reg_492_pp0_iter2_reg;
        icmp_ln47_reg_458_pp0_iter2_reg <= icmp_ln47_reg_458_pp0_iter1_reg;
        icmp_ln47_reg_458_pp0_iter3_reg <= icmp_ln47_reg_458_pp0_iter2_reg;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln47_reg_458 <= icmp_ln47_fu_204_p2;
        icmp_ln47_reg_458_pp0_iter1_reg <= icmp_ln47_reg_458;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_fu_204_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln48_reg_462 <= icmp_ln48_fu_216_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_fu_204_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        select_ln47_6_reg_469 <= select_ln47_6_fu_222_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln47_reg_458 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        select_ln48_11_reg_482 <= select_ln48_11_fu_341_p3;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state1)) begin
        sext_ln47_reg_448 <= sext_ln47_fu_194_p1;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_condition_pp0_exit_iter1_state3 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter1_state3 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln47_fu_204_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_condition_pp0_flush_enable = 1'b1;
    end else begin
        ap_condition_pp0_flush_enable = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state7)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln47_reg_458 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_phi_mux_ii_phi_fu_132_p4 = select_ln47_6_reg_469;
    end else begin
        ap_phi_mux_ii_phi_fu_132_p4 = ii_reg_128;
    end
end

always @ (*) begin
    if (((icmp_ln47_reg_458_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        ap_phi_mux_jj_phi_fu_154_p4 = select_ln48_11_reg_482;
    end else begin
        ap_phi_mux_jj_phi_fu_154_p4 = jj_reg_150;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state7)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter3 == 1'b1)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter4 == 1'b1)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1)))) begin
        filter_data_ce0 = 1'b1;
    end else begin
        filter_data_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        input_indices_23_blk_n = input_indices_23_empty_n;
    end else begin
        input_indices_23_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        input_indices_23_read = 1'b1;
    end else begin
        input_indices_23_read = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter4 == 1'b1))) begin
        weight_vecs_0_ce0 = 1'b1;
    end else begin
        weight_vecs_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln47_reg_458_pp0_iter3_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter4 == 1'b1))) begin
        weight_vecs_0_we0 = 1'b1;
    end else begin
        weight_vecs_0_we0 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_start == 1'b0) | (input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((~((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b0)) & ~((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter4 == 1'b1) & (ap_enable_reg_pp0_iter3 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if ((((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b0)) | ((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter4 == 1'b1) & (ap_enable_reg_pp0_iter3 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_state7;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state7 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln47_6_fu_198_p2 = (indvar_flatten13_reg_117 + 5'd1);

assign add_ln47_fu_210_p2 = (ap_phi_mux_ii_phi_fu_132_p4 + 2'd1);

assign add_ln48_6_fu_230_p2 = (indvar_flatten_reg_139 + 4'd1);

assign add_ln48_fu_322_p2 = (select_ln47_fu_244_p3 + 2'd1);

assign add_ln49_fu_438_p2 = (select_ln48_fu_333_p3 + 2'd1);

assign add_ln55_21_fu_357_p2 = (sub_ln55_11_fu_278_p2 + zext_ln55_54_fu_353_p1);

assign add_ln55_22_fu_385_p2 = ((sext_ln48_fu_301_p1) + (zext_ln55_53_fu_349_p1));

assign add_ln55_23_fu_421_p2 = (sub_ln55_13_fu_379_p2 + zext_ln55_56_fu_417_p1);

assign add_ln55_24_fu_432_p2 = (sub_ln55_14_fu_407_p2 + zext_ln55_55_fu_413_p1);

assign add_ln55_fu_257_p2 = ((sext_ln47_reg_448) + (zext_ln55_51_fu_254_p1));

assign and_ln47_fu_316_p2 = (xor_ln47_fu_305_p2 & icmp_ln49_fu_310_p2);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state7 = ap_CS_fsm[32'd2];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1));
end

assign ap_block_state2_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter4 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign filter_data_address0 = zext_ln55_57_fu_427_p1;

assign icmp_ln47_fu_204_p2 = ((indvar_flatten13_reg_117 == 5'd27) ? 1'b1 : 1'b0);

assign icmp_ln48_fu_216_p2 = ((indvar_flatten_reg_139 == 4'd9) ? 1'b1 : 1'b0);

assign icmp_ln49_fu_310_p2 = ((kk_reg_161 == 2'd3) ? 1'b1 : 1'b0);

assign or_ln48_fu_328_p2 = (icmp_ln48_reg_462 | and_ln47_fu_316_p2);

assign p_shl1_cast_fu_399_p3 = {{trunc_ln55_3_fu_395_p1}, {2'd0}};

assign p_shl2_cast_fu_371_p3 = {{trunc_ln55_1_fu_367_p1}, {2'd0}};

assign select_ln47_6_fu_222_p3 = ((icmp_ln48_fu_216_p2[0:0] == 1'b1) ? add_ln47_fu_210_p2 : ap_phi_mux_ii_phi_fu_132_p4);

assign select_ln47_fu_244_p3 = ((icmp_ln48_reg_462[0:0] == 1'b1) ? 2'd0 : ap_phi_mux_jj_phi_fu_154_p4);

assign select_ln48_11_fu_341_p3 = ((and_ln47_fu_316_p2[0:0] == 1'b1) ? add_ln48_fu_322_p2 : select_ln47_fu_244_p3);

assign select_ln48_12_fu_236_p3 = ((icmp_ln48_fu_216_p2[0:0] == 1'b1) ? 4'd1 : add_ln48_6_fu_230_p2);

assign select_ln48_fu_333_p3 = ((or_ln48_fu_328_p2[0:0] == 1'b1) ? 2'd0 : kk_reg_161);

assign sext_ln47_fu_194_p1 = (sub_ln55_fu_188_p2);

assign sext_ln48_fu_301_p1 = (sub_ln55_12_fu_295_p2);

assign sext_ln55_1_fu_274_p1 = (tmp_46_fu_266_p3);

assign sext_ln55_fu_262_p1 = add_ln55_fu_257_p2;

assign sub_ln55_11_fu_278_p2 = ((sext_ln55_1_fu_274_p1) - (sext_ln55_fu_262_p1));

assign sub_ln55_12_fu_295_p2 = (zext_ln55_52_fu_291_p1 - zext_ln55_50_fu_251_p1);

assign sub_ln55_13_fu_379_p2 = (p_shl2_cast_fu_371_p3 - trunc_ln55_fu_363_p1);

assign sub_ln55_14_fu_407_p2 = (p_shl1_cast_fu_399_p3 - trunc_ln55_2_fu_391_p1);

assign sub_ln55_fu_188_p2 = (zext_ln55_49_fu_184_p1 - zext_ln55_fu_172_p1);

assign tmp_46_fu_266_p3 = {{add_ln55_fu_257_p2}, {2'd0}};

assign tmp_fu_176_p3 = {{input_indices_23_dout}, {2'd0}};

assign tmp_s_fu_284_p3 = {{select_ln47_6_reg_469}, {2'd0}};

assign trunc_ln55_1_fu_367_p1 = add_ln55_21_fu_357_p2[6:0];

assign trunc_ln55_2_fu_391_p1 = add_ln55_22_fu_385_p2[4:0];

assign trunc_ln55_3_fu_395_p1 = add_ln55_22_fu_385_p2[2:0];

assign trunc_ln55_fu_363_p1 = add_ln55_21_fu_357_p2[8:0];

assign weight_vecs_0_address0 = zext_ln55_58_fu_444_p1;

assign weight_vecs_0_d0 = filter_data_q0;

assign xor_ln47_fu_305_p2 = (icmp_ln48_reg_462 ^ 1'd1);

assign zext_ln55_49_fu_184_p1 = tmp_fu_176_p3;

assign zext_ln55_50_fu_251_p1 = select_ln47_6_reg_469;

assign zext_ln55_51_fu_254_p1 = select_ln47_6_reg_469;

assign zext_ln55_52_fu_291_p1 = tmp_s_fu_284_p3;

assign zext_ln55_53_fu_349_p1 = select_ln48_11_fu_341_p3;

assign zext_ln55_54_fu_353_p1 = select_ln48_11_fu_341_p3;

assign zext_ln55_55_fu_413_p1 = select_ln48_fu_333_p3;

assign zext_ln55_56_fu_417_p1 = select_ln48_fu_333_p3;

assign zext_ln55_57_fu_427_p1 = add_ln55_23_fu_421_p2;

assign zext_ln55_58_fu_444_p1 = add_ln55_24_reg_492_pp0_iter3_reg;

assign zext_ln55_fu_172_p1 = input_indices_23_dout;

endmodule //td_fused_top_tdf1_readFilters18
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf1_readInputs19 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        in_data_address0,
        in_data_ce0,
        in_data_q0,
        i_19,
        j_19,
        ifmap_vec_address0,
        ifmap_vec_ce0,
        ifmap_vec_we0,
        ifmap_vec_d0
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state7 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [15:0] in_data_address0;
output   in_data_ce0;
input  [63:0] in_data_q0;
input  [15:0] i_19;
input  [15:0] j_19;
output  [4:0] ifmap_vec_address0;
output   ifmap_vec_ce0;
output   ifmap_vec_we0;
output  [15:0] ifmap_vec_d0;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg in_data_ce0;
reg ifmap_vec_ce0;
reg ifmap_vec_we0;

reg    ap_done_reg;
  reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg   [4:0] indvar_flatten52_reg_144;
reg   [1:0] ii_reg_155;
reg   [3:0] indvar_flatten_reg_167;
reg   [1:0] jj_reg_178;
reg   [1:0] kk_reg_190;
wire   [17:0] p_cast_i_fu_219_p1;
reg   [17:0] p_cast_i_reg_910;
wire   [17:0] sext_ln22_fu_229_p1;
reg   [17:0] sext_ln22_reg_916;
wire   [7:0] p_cast_fu_233_p2;
reg   [7:0] p_cast_reg_922;
wire   [0:0] or_ln23_26_fu_253_p2;
reg   [0:0] or_ln23_26_reg_928;
wire   [15:0] p_mid140_fu_259_p2;
reg   [15:0] p_mid140_reg_933;
wire   [4:0] add_ln19_6_fu_265_p2;
wire    ap_CS_fsm_pp0_stage0;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
wire    ap_block_state4_pp0_stage0_iter2;
wire    ap_block_state5_pp0_stage0_iter3;
wire    ap_block_state6_pp0_stage0_iter4;
wire    ap_block_pp0_stage0_11001;
wire   [0:0] is_padding_fu_315_p2;
reg   [0:0] is_padding_reg_943;
reg   [0:0] is_padding_reg_943_pp0_iter1_reg;
reg   [0:0] is_padding_reg_943_pp0_iter2_reg;
reg   [0:0] is_padding_reg_943_pp0_iter3_reg;
wire   [0:0] icmp_ln19_fu_321_p2;
reg   [0:0] icmp_ln19_reg_950;
reg   [0:0] icmp_ln19_reg_950_pp0_iter1_reg;
reg   [0:0] icmp_ln19_reg_950_pp0_iter2_reg;
reg   [0:0] icmp_ln19_reg_950_pp0_iter3_reg;
wire   [1:0] add_ln19_fu_327_p2;
reg   [1:0] add_ln19_reg_954;
wire   [0:0] icmp_ln20_fu_333_p2;
reg   [0:0] icmp_ln20_reg_959;
reg   [0:0] icmp_ln20_reg_959_pp0_iter1_reg;
reg   [0:0] icmp_ln20_reg_959_pp0_iter2_reg;
reg   [0:0] icmp_ln20_reg_959_pp0_iter3_reg;
wire   [1:0] select_ln19_31_fu_347_p3;
reg   [1:0] select_ln19_31_reg_966;
reg   [1:0] select_ln19_31_reg_966_pp0_iter1_reg;
reg   [1:0] select_ln19_31_reg_966_pp0_iter2_reg;
reg   [1:0] select_ln19_31_reg_966_pp0_iter3_reg;
wire   [0:0] or_ln23_28_fu_378_p2;
reg   [0:0] or_ln23_28_reg_973;
reg   [0:0] or_ln23_28_reg_973_pp0_iter1_reg;
reg   [0:0] or_ln23_28_reg_973_pp0_iter2_reg;
reg   [0:0] or_ln23_28_reg_973_pp0_iter3_reg;
wire   [0:0] and_ln19_fu_395_p2;
reg   [0:0] and_ln19_reg_980;
reg   [0:0] and_ln19_reg_980_pp0_iter1_reg;
reg   [0:0] and_ln19_reg_980_pp0_iter2_reg;
reg   [0:0] and_ln19_reg_980_pp0_iter3_reg;
wire   [1:0] add_ln20_fu_401_p2;
reg   [1:0] add_ln20_reg_986;
wire   [1:0] select_ln20_fu_413_p3;
reg   [1:0] select_ln20_reg_991;
reg   [1:0] select_ln20_reg_991_pp0_iter1_reg;
reg   [1:0] select_ln20_reg_991_pp0_iter2_reg;
reg   [1:0] select_ln20_reg_991_pp0_iter3_reg;
wire   [1:0] select_ln20_26_fu_421_p3;
reg   [1:0] select_ln20_26_reg_997;
reg   [1:0] select_ln20_26_reg_997_pp0_iter1_reg;
reg   [1:0] select_ln20_26_reg_997_pp0_iter2_reg;
reg   [1:0] select_ln20_26_reg_997_pp0_iter3_reg;
wire   [0:0] or_ln23_30_fu_458_p2;
reg   [0:0] or_ln23_30_reg_1003;
reg   [0:0] or_ln23_30_reg_1003_pp0_iter1_reg;
reg   [0:0] or_ln23_30_reg_1003_pp0_iter2_reg;
reg   [0:0] or_ln23_30_reg_1003_pp0_iter3_reg;
wire   [1:0] add_ln25_fu_464_p2;
wire   [3:0] select_ln20_29_fu_476_p3;
wire   [5:0] tmp_15_fu_701_p3;
reg   [5:0] tmp_15_reg_1025;
wire   [5:0] empty_121_fu_708_p2;
reg   [5:0] empty_121_reg_1030;
wire   [0:0] icmp_ln32_fu_714_p2;
reg   [0:0] icmp_ln32_reg_1035;
reg    ap_block_state1;
wire    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_flush_enable;
reg    ap_enable_reg_pp0_iter1;
reg    ap_enable_reg_pp0_iter2;
reg    ap_condition_pp0_exit_iter1_state3;
reg    ap_enable_reg_pp0_iter3;
reg    ap_enable_reg_pp0_iter4;
reg   [1:0] ap_phi_mux_ii_phi_fu_159_p4;
wire    ap_block_pp0_stage0;
reg   [1:0] ap_phi_mux_jj_phi_fu_182_p4;
wire   [63:0] zext_ln32_26_fu_696_p1;
wire   [63:0] zext_ln33_25_fu_795_p1;
wire   [16:0] zext_ln19_fu_205_p1;
wire   [16:0] empty_116_fu_213_p2;
wire   [16:0] j_cast_i_fu_201_p1;
wire   [16:0] add_ln22_fu_223_p2;
wire   [7:0] empty_fu_209_p1;
wire   [0:0] tmp_fu_239_p3;
wire   [0:0] icmp_ln24_fu_247_p2;
wire   [17:0] ii_cast_i_fu_271_p1;
wire   [17:0] empty_117_fu_275_p2;
wire   [17:0] zext_ln20_fu_286_p1;
wire   [17:0] add_ln22_6_fu_290_p2;
wire   [0:0] tmp_43_fu_295_p3;
wire   [0:0] icmp_ln24_6_fu_303_p2;
wire   [0:0] or_ln23_fu_309_p2;
wire   [0:0] empty_118_fu_280_p2;
wire   [17:0] ii_cast_i_mid1_fu_355_p1;
wire   [17:0] p_mid114_fu_359_p2;
wire   [0:0] p_mid116_fu_364_p2;
wire   [0:0] icmp_ln25_fu_389_p2;
wire   [0:0] xor_ln19_fu_383_p2;
wire   [1:0] select_ln19_fu_339_p3;
wire   [0:0] or_ln20_fu_407_p2;
wire   [17:0] zext_ln20_6_fu_429_p1;
wire   [17:0] add_ln22_7_fu_433_p2;
wire   [0:0] tmp_44_fu_438_p3;
wire   [0:0] icmp_ln24_7_fu_446_p2;
wire   [0:0] or_ln23_29_fu_452_p2;
wire   [0:0] select_ln19_33_fu_370_p3;
wire   [3:0] add_ln20_6_fu_470_p2;
wire   [7:0] ii_cast_fu_484_p1;
wire   [7:0] p_cast1_i_fu_488_p2;
wire   [2:0] zext_ln22_fu_493_p1;
wire   [2:0] tmp2_fu_504_p2;
wire   [15:0] tmp2_cast_fu_510_p1;
wire   [15:0] empty_119_fu_514_p2;
wire   [7:0] row_coord_int_fu_497_p3;
wire   [12:0] tmp_9_fu_534_p3;
wire   [15:0] tmp_s_fu_526_p3;
wire   [15:0] zext_ln32_fu_542_p1;
wire   [15:0] sub_ln32_fu_546_p2;
wire   [15:0] col_coord_int_fu_519_p3;
wire   [7:0] ii_cast_mid1_fu_558_p1;
wire   [7:0] p_cast1_i_mid1_fu_561_p2;
wire   [7:0] row_coord_int_mid134_fu_573_p3;
wire   [12:0] tmp_12_fu_594_p3;
wire   [15:0] tmp_11_fu_586_p3;
wire   [15:0] zext_ln32_24_fu_602_p1;
wire   [15:0] sub_ln32_1_fu_606_p2;
wire   [15:0] col_coord_int_mid142_fu_580_p3;
wire   [15:0] add_ln32_1_fu_612_p2;
wire   [15:0] add_ln32_fu_552_p2;
wire   [7:0] select_ln19_32_fu_566_p3;
wire   [2:0] zext_ln22_6_fu_625_p1;
wire   [2:0] tmp2_mid1_fu_635_p2;
wire   [15:0] tmp2_cast_mid1_fu_641_p1;
wire   [15:0] p_mid1_fu_645_p2;
wire   [7:0] row_coord_int_mid1_fu_628_p3;
wire   [12:0] tmp_14_fu_665_p3;
wire   [15:0] tmp_13_fu_657_p3;
wire   [15:0] zext_ln32_25_fu_673_p1;
wire   [15:0] sub_ln32_2_fu_677_p2;
wire   [15:0] col_coord_int_mid1_fu_650_p3;
wire   [15:0] add_ln32_2_fu_683_p2;
wire   [15:0] select_ln19_35_fu_618_p3;
wire   [15:0] select_ln20_28_fu_689_p3;
wire   [3:0] tmp_10_fu_723_p3;
wire   [4:0] zext_ln33_22_fu_730_p1;
wire   [4:0] zext_ln33_fu_720_p1;
wire   [4:0] sub_ln33_fu_734_p2;
wire   [5:0] sub_ln33_cast_fu_740_p1;
wire   [5:0] zext_ln33_23_fu_749_p1;
wire   [5:0] add_ln33_fu_752_p2;
wire   [2:0] trunc_ln33_1_fu_762_p1;
wire   [4:0] p_shl4_cast_fu_766_p3;
wire   [4:0] trunc_ln33_fu_758_p1;
wire   [0:0] select_ln19_34_fu_744_p3;
wire   [4:0] sub_ln33_1_fu_774_p2;
wire   [4:0] zext_ln33_24_fu_786_p1;
wire   [4:0] add_ln33_6_fu_789_p2;
wire   [6:0] zext_ln32_27_fu_800_p1;
wire   [6:0] zext_ln32_28_fu_803_p1;
wire   [6:0] sub_ln32_3_fu_816_p2;
wire   [6:0] sub_ln32_4_fu_828_p2;
reg   [63:0] tmp_45_fu_806_p4;
wire   [6:0] xor_ln32_fu_822_p2;
wire   [6:0] select_ln32_fu_834_p3;
wire   [6:0] select_ln32_2_fu_848_p3;
wire   [6:0] sub_ln32_5_fu_855_p2;
wire   [63:0] select_ln32_1_fu_841_p3;
wire   [63:0] zext_ln32_29_fu_861_p1;
wire   [63:0] zext_ln32_30_fu_865_p1;
wire   [63:0] lshr_ln32_fu_869_p2;
wire   [63:0] lshr_ln32_1_fu_875_p2;
wire   [63:0] and_ln32_fu_881_p2;
wire   [15:0] trunc_ln32_fu_887_p1;
wire   [0:0] select_ln20_27_fu_780_p3;
wire   [15:0] in_data_elem_fu_891_p1;
wire    ap_CS_fsm_state7;
reg   [2:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
#0 ap_enable_reg_pp0_iter4 = 1'b0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state7)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if ((1'b1 == ap_condition_pp0_flush_enable)) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            if ((1'b1 == ap_condition_pp0_exit_iter1_state3)) begin
                ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter0;
            end else if ((1'b1 == 1'b1)) begin
                ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
            end
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter4 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
        end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter4 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln19_reg_950 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ii_reg_155 <= select_ln19_31_reg_966;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ii_reg_155 <= 2'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln19_fu_321_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        indvar_flatten52_reg_144 <= add_ln19_6_fu_265_p2;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indvar_flatten52_reg_144 <= 5'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln19_fu_321_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        indvar_flatten_reg_167 <= select_ln20_29_fu_476_p3;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indvar_flatten_reg_167 <= 4'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln19_reg_950 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        jj_reg_178 <= select_ln20_26_reg_997;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        jj_reg_178 <= 2'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln19_fu_321_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        kk_reg_190 <= add_ln25_fu_464_p2;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        kk_reg_190 <= 2'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln19_fu_321_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        add_ln19_reg_954 <= add_ln19_fu_327_p2;
        add_ln20_reg_986 <= add_ln20_fu_401_p2;
        and_ln19_reg_980 <= and_ln19_fu_395_p2;
        icmp_ln20_reg_959 <= icmp_ln20_fu_333_p2;
        or_ln23_28_reg_973 <= or_ln23_28_fu_378_p2;
        or_ln23_30_reg_1003 <= or_ln23_30_fu_458_p2;
        select_ln20_reg_991 <= select_ln20_fu_413_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        and_ln19_reg_980_pp0_iter1_reg <= and_ln19_reg_980;
        icmp_ln19_reg_950 <= icmp_ln19_fu_321_p2;
        icmp_ln19_reg_950_pp0_iter1_reg <= icmp_ln19_reg_950;
        icmp_ln20_reg_959_pp0_iter1_reg <= icmp_ln20_reg_959;
        is_padding_reg_943 <= is_padding_fu_315_p2;
        is_padding_reg_943_pp0_iter1_reg <= is_padding_reg_943;
        or_ln23_28_reg_973_pp0_iter1_reg <= or_ln23_28_reg_973;
        or_ln23_30_reg_1003_pp0_iter1_reg <= or_ln23_30_reg_1003;
        select_ln19_31_reg_966_pp0_iter1_reg <= select_ln19_31_reg_966;
        select_ln20_26_reg_997_pp0_iter1_reg <= select_ln20_26_reg_997;
        select_ln20_reg_991_pp0_iter1_reg <= select_ln20_reg_991;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        and_ln19_reg_980_pp0_iter2_reg <= and_ln19_reg_980_pp0_iter1_reg;
        and_ln19_reg_980_pp0_iter3_reg <= and_ln19_reg_980_pp0_iter2_reg;
        icmp_ln19_reg_950_pp0_iter2_reg <= icmp_ln19_reg_950_pp0_iter1_reg;
        icmp_ln19_reg_950_pp0_iter3_reg <= icmp_ln19_reg_950_pp0_iter2_reg;
        icmp_ln20_reg_959_pp0_iter2_reg <= icmp_ln20_reg_959_pp0_iter1_reg;
        icmp_ln20_reg_959_pp0_iter3_reg <= icmp_ln20_reg_959_pp0_iter2_reg;
        is_padding_reg_943_pp0_iter2_reg <= is_padding_reg_943_pp0_iter1_reg;
        is_padding_reg_943_pp0_iter3_reg <= is_padding_reg_943_pp0_iter2_reg;
        or_ln23_28_reg_973_pp0_iter2_reg <= or_ln23_28_reg_973_pp0_iter1_reg;
        or_ln23_28_reg_973_pp0_iter3_reg <= or_ln23_28_reg_973_pp0_iter2_reg;
        or_ln23_30_reg_1003_pp0_iter2_reg <= or_ln23_30_reg_1003_pp0_iter1_reg;
        or_ln23_30_reg_1003_pp0_iter3_reg <= or_ln23_30_reg_1003_pp0_iter2_reg;
        select_ln19_31_reg_966_pp0_iter2_reg <= select_ln19_31_reg_966_pp0_iter1_reg;
        select_ln19_31_reg_966_pp0_iter3_reg <= select_ln19_31_reg_966_pp0_iter2_reg;
        select_ln20_26_reg_997_pp0_iter2_reg <= select_ln20_26_reg_997_pp0_iter1_reg;
        select_ln20_26_reg_997_pp0_iter3_reg <= select_ln20_26_reg_997_pp0_iter2_reg;
        select_ln20_reg_991_pp0_iter2_reg <= select_ln20_reg_991_pp0_iter1_reg;
        select_ln20_reg_991_pp0_iter3_reg <= select_ln20_reg_991_pp0_iter2_reg;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln19_reg_950_pp0_iter2_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        empty_121_reg_1030[5 : 4] <= empty_121_fu_708_p2[5 : 4];
        icmp_ln32_reg_1035 <= icmp_ln32_fu_714_p2;
        tmp_15_reg_1025[5 : 4] <= tmp_15_fu_701_p3[5 : 4];
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state1)) begin
        or_ln23_26_reg_928 <= or_ln23_26_fu_253_p2;
        p_cast_i_reg_910 <= p_cast_i_fu_219_p1;
        p_cast_reg_922 <= p_cast_fu_233_p2;
        p_mid140_reg_933 <= p_mid140_fu_259_p2;
        sext_ln22_reg_916 <= sext_ln22_fu_229_p1;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln19_fu_321_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        select_ln19_31_reg_966 <= select_ln19_31_fu_347_p3;
        select_ln20_26_reg_997 <= select_ln20_26_fu_421_p3;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_condition_pp0_exit_iter1_state3 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter1_state3 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln19_fu_321_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_condition_pp0_flush_enable = 1'b1;
    end else begin
        ap_condition_pp0_flush_enable = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state7)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln19_reg_950 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_ii_phi_fu_159_p4 = select_ln19_31_reg_966;
    end else begin
        ap_phi_mux_ii_phi_fu_159_p4 = ii_reg_155;
    end
end

always @ (*) begin
    if (((icmp_ln19_reg_950 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_jj_phi_fu_182_p4 = select_ln20_26_reg_997;
    end else begin
        ap_phi_mux_jj_phi_fu_182_p4 = jj_reg_178;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state7)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter4 == 1'b1))) begin
        ifmap_vec_ce0 = 1'b1;
    end else begin
        ifmap_vec_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln19_reg_950_pp0_iter3_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter4 == 1'b1))) begin
        ifmap_vec_we0 = 1'b1;
    end else begin
        ifmap_vec_we0 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter3 == 1'b1)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter4 == 1'b1)))) begin
        in_data_ce0 = 1'b1;
    end else begin
        in_data_ce0 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((~((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b1)) & ~((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter4 == 1'b1) & (ap_enable_reg_pp0_iter3 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if ((((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter4 == 1'b1) & (ap_enable_reg_pp0_iter3 == 1'b0)) | ((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b1)))) begin
                ap_NS_fsm = ap_ST_fsm_state7;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state7 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln19_6_fu_265_p2 = (indvar_flatten52_reg_144 + 5'd1);

assign add_ln19_fu_327_p2 = (ap_phi_mux_ii_phi_fu_159_p4 + 2'd1);

assign add_ln20_6_fu_470_p2 = (indvar_flatten_reg_167 + 4'd1);

assign add_ln20_fu_401_p2 = (select_ln19_fu_339_p3 + 2'd1);

assign add_ln22_6_fu_290_p2 = ((sext_ln22_reg_916) + (zext_ln20_fu_286_p1));

assign add_ln22_7_fu_433_p2 = ((sext_ln22_reg_916) + (zext_ln20_6_fu_429_p1));

assign add_ln22_fu_223_p2 = ((j_cast_i_fu_201_p1) + (17'd131071));

assign add_ln25_fu_464_p2 = (select_ln20_fu_413_p3 + 2'd1);

assign add_ln32_1_fu_612_p2 = (sub_ln32_1_fu_606_p2 + col_coord_int_mid142_fu_580_p3);

assign add_ln32_2_fu_683_p2 = (sub_ln32_2_fu_677_p2 + col_coord_int_mid1_fu_650_p3);

assign add_ln32_fu_552_p2 = (sub_ln32_fu_546_p2 + col_coord_int_fu_519_p3);

assign add_ln33_6_fu_789_p2 = (sub_ln33_1_fu_774_p2 + zext_ln33_24_fu_786_p1);

assign add_ln33_fu_752_p2 = ((sub_ln33_cast_fu_740_p1) + (zext_ln33_23_fu_749_p1));

assign and_ln19_fu_395_p2 = (xor_ln19_fu_383_p2 & icmp_ln25_fu_389_p2);

assign and_ln32_fu_881_p2 = (lshr_ln32_fu_869_p2 & lshr_ln32_1_fu_875_p2);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state7 = ap_CS_fsm[32'd2];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (ap_done_reg == 1'b1));
end

assign ap_block_state2_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter4 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign col_coord_int_fu_519_p3 = ((is_padding_reg_943[0:0] == 1'b1) ? 16'd0 : empty_119_fu_514_p2);

assign col_coord_int_mid142_fu_580_p3 = ((or_ln23_28_reg_973[0:0] == 1'b1) ? 16'd0 : p_mid140_reg_933);

assign col_coord_int_mid1_fu_650_p3 = ((or_ln23_30_reg_1003[0:0] == 1'b1) ? 16'd0 : p_mid1_fu_645_p2);

assign empty_116_fu_213_p2 = ((zext_ln19_fu_205_p1) + (17'd131071));

assign empty_117_fu_275_p2 = ((p_cast_i_reg_910) + (ii_cast_i_fu_271_p1));

assign empty_118_fu_280_p2 = ((empty_117_fu_275_p2 > 18'd223) ? 1'b1 : 1'b0);

assign empty_119_fu_514_p2 = ((tmp2_cast_fu_510_p1) + (j_19));

assign empty_121_fu_708_p2 = (tmp_15_fu_701_p3 | 6'd15);

assign empty_fu_209_p1 = i_19[7:0];

assign icmp_ln19_fu_321_p2 = ((indvar_flatten52_reg_144 == 5'd27) ? 1'b1 : 1'b0);

assign icmp_ln20_fu_333_p2 = ((indvar_flatten_reg_167 == 4'd9) ? 1'b1 : 1'b0);

assign icmp_ln24_6_fu_303_p2 = (((add_ln22_6_fu_290_p2) > (18'd223)) ? 1'b1 : 1'b0);

assign icmp_ln24_7_fu_446_p2 = (((add_ln22_7_fu_433_p2) > (18'd223)) ? 1'b1 : 1'b0);

assign icmp_ln24_fu_247_p2 = (((add_ln22_fu_223_p2) > (17'd223)) ? 1'b1 : 1'b0);

assign icmp_ln25_fu_389_p2 = ((kk_reg_190 == 2'd3) ? 1'b1 : 1'b0);

assign icmp_ln32_fu_714_p2 = ((tmp_15_fu_701_p3 > empty_121_fu_708_p2) ? 1'b1 : 1'b0);

assign ifmap_vec_address0 = zext_ln33_25_fu_795_p1;

assign ifmap_vec_d0 = ((select_ln20_27_fu_780_p3[0:0] == 1'b1) ? 16'd0 : in_data_elem_fu_891_p1);

assign ii_cast_fu_484_p1 = ii_reg_155;

assign ii_cast_i_fu_271_p1 = ap_phi_mux_ii_phi_fu_159_p4;

assign ii_cast_i_mid1_fu_355_p1 = add_ln19_fu_327_p2;

assign ii_cast_mid1_fu_558_p1 = add_ln19_reg_954;

assign in_data_address0 = zext_ln32_26_fu_696_p1;

assign in_data_elem_fu_891_p1 = trunc_ln32_fu_887_p1;

assign is_padding_fu_315_p2 = (or_ln23_fu_309_p2 | empty_118_fu_280_p2);

assign j_cast_i_fu_201_p1 = j_19;

assign lshr_ln32_1_fu_875_p2 = 64'd18446744073709551615 >> zext_ln32_30_fu_865_p1;

assign lshr_ln32_fu_869_p2 = select_ln32_1_fu_841_p3 >> zext_ln32_29_fu_861_p1;

assign or_ln20_fu_407_p2 = (icmp_ln20_fu_333_p2 | and_ln19_fu_395_p2);

assign or_ln23_26_fu_253_p2 = (tmp_fu_239_p3 | icmp_ln24_fu_247_p2);

assign or_ln23_28_fu_378_p2 = (p_mid116_fu_364_p2 | or_ln23_26_reg_928);

assign or_ln23_29_fu_452_p2 = (tmp_44_fu_438_p3 | icmp_ln24_7_fu_446_p2);

assign or_ln23_30_fu_458_p2 = (select_ln19_33_fu_370_p3 | or_ln23_29_fu_452_p2);

assign or_ln23_fu_309_p2 = (tmp_43_fu_295_p3 | icmp_ln24_6_fu_303_p2);

assign p_cast1_i_fu_488_p2 = (p_cast_reg_922 + ii_cast_fu_484_p1);

assign p_cast1_i_mid1_fu_561_p2 = (p_cast_reg_922 + ii_cast_mid1_fu_558_p1);

assign p_cast_fu_233_p2 = ((empty_fu_209_p1) + (8'd255));

assign p_cast_i_fu_219_p1 = (empty_116_fu_213_p2);

assign p_mid114_fu_359_p2 = ((p_cast_i_reg_910) + (ii_cast_i_mid1_fu_355_p1));

assign p_mid116_fu_364_p2 = ((p_mid114_fu_359_p2 > 18'd223) ? 1'b1 : 1'b0);

assign p_mid140_fu_259_p2 = ((j_19) + (16'd65535));

assign p_mid1_fu_645_p2 = ((tmp2_cast_mid1_fu_641_p1) + (j_19));

assign p_shl4_cast_fu_766_p3 = {{trunc_ln33_1_fu_762_p1}, {2'd0}};

assign row_coord_int_fu_497_p3 = ((is_padding_reg_943[0:0] == 1'b1) ? 8'd0 : p_cast1_i_fu_488_p2);

assign row_coord_int_mid134_fu_573_p3 = ((or_ln23_28_reg_973[0:0] == 1'b1) ? 8'd0 : p_cast1_i_mid1_fu_561_p2);

assign row_coord_int_mid1_fu_628_p3 = ((or_ln23_30_reg_1003[0:0] == 1'b1) ? 8'd0 : select_ln19_32_fu_566_p3);

assign select_ln19_31_fu_347_p3 = ((icmp_ln20_fu_333_p2[0:0] == 1'b1) ? add_ln19_fu_327_p2 : ap_phi_mux_ii_phi_fu_159_p4);

assign select_ln19_32_fu_566_p3 = ((icmp_ln20_reg_959[0:0] == 1'b1) ? p_cast1_i_mid1_fu_561_p2 : p_cast1_i_fu_488_p2);

assign select_ln19_33_fu_370_p3 = ((icmp_ln20_fu_333_p2[0:0] == 1'b1) ? p_mid116_fu_364_p2 : empty_118_fu_280_p2);

assign select_ln19_34_fu_744_p3 = ((icmp_ln20_reg_959_pp0_iter3_reg[0:0] == 1'b1) ? or_ln23_28_reg_973_pp0_iter3_reg : is_padding_reg_943_pp0_iter3_reg);

assign select_ln19_35_fu_618_p3 = ((icmp_ln20_reg_959[0:0] == 1'b1) ? add_ln32_1_fu_612_p2 : add_ln32_fu_552_p2);

assign select_ln19_fu_339_p3 = ((icmp_ln20_fu_333_p2[0:0] == 1'b1) ? 2'd0 : ap_phi_mux_jj_phi_fu_182_p4);

assign select_ln20_26_fu_421_p3 = ((and_ln19_fu_395_p2[0:0] == 1'b1) ? add_ln20_fu_401_p2 : select_ln19_fu_339_p3);

assign select_ln20_27_fu_780_p3 = ((and_ln19_reg_980_pp0_iter3_reg[0:0] == 1'b1) ? or_ln23_30_reg_1003_pp0_iter3_reg : select_ln19_34_fu_744_p3);

assign select_ln20_28_fu_689_p3 = ((and_ln19_reg_980[0:0] == 1'b1) ? add_ln32_2_fu_683_p2 : select_ln19_35_fu_618_p3);

assign select_ln20_29_fu_476_p3 = ((icmp_ln20_fu_333_p2[0:0] == 1'b1) ? 4'd1 : add_ln20_6_fu_470_p2);

assign select_ln20_fu_413_p3 = ((or_ln20_fu_407_p2[0:0] == 1'b1) ? 2'd0 : kk_reg_190);

assign select_ln32_1_fu_841_p3 = ((icmp_ln32_reg_1035[0:0] == 1'b1) ? tmp_45_fu_806_p4 : in_data_q0);

assign select_ln32_2_fu_848_p3 = ((icmp_ln32_reg_1035[0:0] == 1'b1) ? xor_ln32_fu_822_p2 : zext_ln32_27_fu_800_p1);

assign select_ln32_fu_834_p3 = ((icmp_ln32_reg_1035[0:0] == 1'b1) ? sub_ln32_3_fu_816_p2 : sub_ln32_4_fu_828_p2);

assign sext_ln22_fu_229_p1 = add_ln22_fu_223_p2;

assign sub_ln32_1_fu_606_p2 = (tmp_11_fu_586_p3 - zext_ln32_24_fu_602_p1);

assign sub_ln32_2_fu_677_p2 = (tmp_13_fu_657_p3 - zext_ln32_25_fu_673_p1);

assign sub_ln32_3_fu_816_p2 = (zext_ln32_27_fu_800_p1 - zext_ln32_28_fu_803_p1);

assign sub_ln32_4_fu_828_p2 = (zext_ln32_28_fu_803_p1 - zext_ln32_27_fu_800_p1);

assign sub_ln32_5_fu_855_p2 = (7'd63 - select_ln32_fu_834_p3);

assign sub_ln32_fu_546_p2 = (tmp_s_fu_526_p3 - zext_ln32_fu_542_p1);

assign sub_ln33_1_fu_774_p2 = (p_shl4_cast_fu_766_p3 - trunc_ln33_fu_758_p1);

assign sub_ln33_cast_fu_740_p1 = (sub_ln33_fu_734_p2);

assign sub_ln33_fu_734_p2 = (zext_ln33_22_fu_730_p1 - zext_ln33_fu_720_p1);

assign tmp2_cast_fu_510_p1 = (tmp2_fu_504_p2);

assign tmp2_cast_mid1_fu_641_p1 = (tmp2_mid1_fu_635_p2);

assign tmp2_fu_504_p2 = ((zext_ln22_fu_493_p1) + (3'd7));

assign tmp2_mid1_fu_635_p2 = ((zext_ln22_6_fu_625_p1) + (3'd7));

assign tmp_10_fu_723_p3 = {{select_ln19_31_reg_966_pp0_iter3_reg}, {2'd0}};

assign tmp_11_fu_586_p3 = {{row_coord_int_mid134_fu_573_p3}, {8'd0}};

assign tmp_12_fu_594_p3 = {{row_coord_int_mid134_fu_573_p3}, {5'd0}};

assign tmp_13_fu_657_p3 = {{row_coord_int_mid1_fu_628_p3}, {8'd0}};

assign tmp_14_fu_665_p3 = {{row_coord_int_mid1_fu_628_p3}, {5'd0}};

assign tmp_15_fu_701_p3 = {{select_ln20_reg_991_pp0_iter2_reg}, {4'd0}};

assign tmp_43_fu_295_p3 = add_ln22_6_fu_290_p2[32'd17];

assign tmp_44_fu_438_p3 = add_ln22_7_fu_433_p2[32'd17];

integer ap_tvar_int_0;

always @ (in_data_q0) begin
    //for (ap_tvar_int_0 = 64 - 1; ap_tvar_int_0 >= 0; ap_tvar_int_0 = ap_tvar_int_0 - 1) begin
    for (ap_tvar_int_0 = 0; ap_tvar_int_0 < 64; ap_tvar_int_0 = ap_tvar_int_0 + 1) begin
        if (ap_tvar_int_0 > 63 - 0) begin
            tmp_45_fu_806_p4[ap_tvar_int_0] = 1'b0;
        end else begin
            tmp_45_fu_806_p4[ap_tvar_int_0] = in_data_q0[63 - ap_tvar_int_0];
        end
    end
end

assign tmp_9_fu_534_p3 = {{row_coord_int_fu_497_p3}, {5'd0}};

assign tmp_fu_239_p3 = add_ln22_fu_223_p2[32'd16];

assign tmp_s_fu_526_p3 = {{row_coord_int_fu_497_p3}, {8'd0}};

assign trunc_ln32_fu_887_p1 = and_ln32_fu_881_p2[15:0];

assign trunc_ln33_1_fu_762_p1 = add_ln33_fu_752_p2[2:0];

assign trunc_ln33_fu_758_p1 = add_ln33_fu_752_p2[4:0];

assign xor_ln19_fu_383_p2 = (icmp_ln20_fu_333_p2 ^ 1'd1);

assign xor_ln32_fu_822_p2 = (zext_ln32_27_fu_800_p1 ^ 7'd63);

assign zext_ln19_fu_205_p1 = i_19;

assign zext_ln20_6_fu_429_p1 = add_ln20_fu_401_p2;

assign zext_ln20_fu_286_p1 = ap_phi_mux_jj_phi_fu_182_p4;

assign zext_ln22_6_fu_625_p1 = add_ln20_reg_986;

assign zext_ln22_fu_493_p1 = jj_reg_178;

assign zext_ln32_24_fu_602_p1 = tmp_12_fu_594_p3;

assign zext_ln32_25_fu_673_p1 = tmp_14_fu_665_p3;

assign zext_ln32_26_fu_696_p1 = select_ln20_28_fu_689_p3;

assign zext_ln32_27_fu_800_p1 = tmp_15_reg_1025;

assign zext_ln32_28_fu_803_p1 = empty_121_reg_1030;

assign zext_ln32_29_fu_861_p1 = select_ln32_2_fu_848_p3;

assign zext_ln32_30_fu_865_p1 = sub_ln32_5_fu_855_p2;

assign zext_ln32_fu_542_p1 = tmp_9_fu_534_p3;

assign zext_ln33_22_fu_730_p1 = tmp_10_fu_723_p3;

assign zext_ln33_23_fu_749_p1 = select_ln20_26_reg_997_pp0_iter3_reg;

assign zext_ln33_24_fu_786_p1 = select_ln20_reg_991_pp0_iter3_reg;

assign zext_ln33_25_fu_795_p1 = add_ln33_6_fu_789_p2;

assign zext_ln33_fu_720_p1 = select_ln19_31_reg_966_pp0_iter3_reg;

always @ (posedge ap_clk) begin
    tmp_15_reg_1025[3:0] <= 4'b0000;
    empty_121_reg_1030[3:0] <= 4'b1111;
end

endmodule //td_fused_top_tdf1_readInputs19
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf1_writeOutputs_unaligned (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        i,
        j,
        out_data_address1,
        out_data_ce1,
        out_data_we1,
        out_data_d1,
        max_vals_3_0
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_state2 = 3'd2;
parameter    ap_ST_fsm_state3 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
input  [6:0] i;
input  [13:0] j;
output  [15:0] out_data_address1;
output   out_data_ce1;
output   out_data_we1;
output  [63:0] out_data_d1;
input  [15:0] max_vals_3_0;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg out_data_ce1;
reg out_data_we1;

  reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg   [15:0] outputCount_1;
reg   [15:0] outputChanIdx_1;
reg   [15:0] outputRow_8_0;
reg   [15:0] outputRow_8_1;
reg   [15:0] outputRow_8_2;
reg   [15:0] outputRow_8_3;
wire   [14:0] sub_ln94_fu_121_p2;
reg   [14:0] sub_ln94_reg_294;
wire   [15:0] add_ln87_fu_182_p2;
wire    ap_CS_fsm_state2;
wire   [0:0] icmp_ln88_fu_188_p2;
reg   [0:0] icmp_ln88_reg_307;
reg   [15:0] ap_phi_mux_empty_phi_fu_90_p4;
reg   [15:0] empty_reg_87;
wire    ap_CS_fsm_state3;
wire   [63:0] zext_ln94_18_fu_216_p1;
wire   [15:0] select_ln97_fu_274_p3;
wire   [1:0] trunc_ln86_fu_154_p1;
reg   [15:0] ap_sig_allocacmp_outputRow_8_0_load;
reg   [15:0] ap_sig_allocacmp_outputRow_8_1_load;
reg   [15:0] ap_sig_allocacmp_outputRow_8_2_load;
reg   [15:0] ap_sig_allocacmp_outputRow_8_3_load;
wire   [13:0] tmp_fu_97_p3;
wire   [10:0] tmp_s_fu_109_p3;
wire   [14:0] zext_ln94_fu_105_p1;
wire   [14:0] zext_ln94_15_fu_117_p1;
wire   [15:0] sub_ln94_cast14_fu_127_p1;
wire   [15:0] zext_ln94_16_fu_130_p1;
wire   [15:0] add_ln94_fu_134_p2;
wire   [3:0] trunc_ln94_fu_202_p1;
wire   [15:0] shl_ln89_fu_140_p2;
wire   [15:0] zext_ln94_17_fu_206_p1;
wire   [15:0] add_ln94_7_fu_210_p2;
wire   [15:0] bitcast_ln94_21_fu_245_p1;
wire   [15:0] bitcast_ln94_20_fu_237_p1;
wire   [15:0] bitcast_ln94_19_fu_229_p1;
wire   [15:0] bitcast_ln94_fu_221_p1;
wire   [15:0] add_ln96_fu_262_p2;
wire   [0:0] icmp_ln97_fu_268_p2;
reg   [2:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_CS_fsm = 3'd1;
#0 outputCount_1 = 16'd0;
#0 outputChanIdx_1 = 16'd0;
#0 outputRow_8_0 = 16'd0;
#0 outputRow_8_1 = 16'd0;
#0 outputRow_8_2 = 16'd0;
#0 outputRow_8_3 = 16'd0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln88_reg_307 == 1'd1) & (1'b1 == ap_CS_fsm_state3))) begin
        empty_reg_87 <= 16'd0;
    end else if (((icmp_ln88_fu_188_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state2))) begin
        empty_reg_87 <= add_ln87_fu_182_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        icmp_ln88_reg_307 <= icmp_ln88_fu_188_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln88_fu_188_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        outputChanIdx_1 <= select_ln97_fu_274_p3;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state3)) begin
        outputCount_1 <= ap_phi_mux_empty_phi_fu_90_p4;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln86_fu_154_p1 == 2'd0) & (1'b1 == ap_CS_fsm_state2))) begin
        outputRow_8_0 <= max_vals_3_0;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln86_fu_154_p1 == 2'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        outputRow_8_1 <= max_vals_3_0;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln86_fu_154_p1 == 2'd2) & (1'b1 == ap_CS_fsm_state2))) begin
        outputRow_8_2 <= max_vals_3_0;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln86_fu_154_p1 == 2'd3) & (1'b1 == ap_CS_fsm_state2))) begin
        outputRow_8_3 <= max_vals_3_0;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state1)) begin
        sub_ln94_reg_294[14 : 4] <= sub_ln94_fu_121_p2[14 : 4];
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state3) | ((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1)))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = 1'b0;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln88_reg_307 == 1'd1) & (1'b1 == ap_CS_fsm_state3))) begin
        ap_phi_mux_empty_phi_fu_90_p4 = 16'd0;
    end else begin
        ap_phi_mux_empty_phi_fu_90_p4 = empty_reg_87;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state3)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((trunc_ln86_fu_154_p1 == 2'd0) & (1'b1 == ap_CS_fsm_state2))) begin
        ap_sig_allocacmp_outputRow_8_0_load = max_vals_3_0;
    end else begin
        ap_sig_allocacmp_outputRow_8_0_load = outputRow_8_0;
    end
end

always @ (*) begin
    if (((trunc_ln86_fu_154_p1 == 2'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        ap_sig_allocacmp_outputRow_8_1_load = max_vals_3_0;
    end else begin
        ap_sig_allocacmp_outputRow_8_1_load = outputRow_8_1;
    end
end

always @ (*) begin
    if (((trunc_ln86_fu_154_p1 == 2'd2) & (1'b1 == ap_CS_fsm_state2))) begin
        ap_sig_allocacmp_outputRow_8_2_load = max_vals_3_0;
    end else begin
        ap_sig_allocacmp_outputRow_8_2_load = outputRow_8_2;
    end
end

always @ (*) begin
    if (((trunc_ln86_fu_154_p1 == 2'd3) & (1'b1 == ap_CS_fsm_state2))) begin
        ap_sig_allocacmp_outputRow_8_3_load = max_vals_3_0;
    end else begin
        ap_sig_allocacmp_outputRow_8_3_load = outputRow_8_3;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state2))) begin
        out_data_ce1 = 1'b1;
    end else begin
        out_data_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln88_fu_188_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        out_data_we1 = 1'b1;
    end else begin
        out_data_we1 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_state2 : begin
            ap_NS_fsm = ap_ST_fsm_state3;
        end
        ap_ST_fsm_state3 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln87_fu_182_p2 = (outputCount_1 + 16'd1);

assign add_ln94_7_fu_210_p2 = (shl_ln89_fu_140_p2 + zext_ln94_17_fu_206_p1);

assign add_ln94_fu_134_p2 = (sub_ln94_cast14_fu_127_p1 + zext_ln94_16_fu_130_p1);

assign add_ln96_fu_262_p2 = (outputChanIdx_1 + 16'd1);

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign bitcast_ln94_19_fu_229_p1 = ap_sig_allocacmp_outputRow_8_1_load;

assign bitcast_ln94_20_fu_237_p1 = ap_sig_allocacmp_outputRow_8_2_load;

assign bitcast_ln94_21_fu_245_p1 = ap_sig_allocacmp_outputRow_8_3_load;

assign bitcast_ln94_fu_221_p1 = ap_sig_allocacmp_outputRow_8_0_load;

assign icmp_ln88_fu_188_p2 = ((add_ln87_fu_182_p2 == 16'd4) ? 1'b1 : 1'b0);

assign icmp_ln97_fu_268_p2 = ((add_ln96_fu_262_p2 == 16'd4) ? 1'b1 : 1'b0);

assign out_data_address1 = zext_ln94_18_fu_216_p1;

assign out_data_d1 = {{{{bitcast_ln94_21_fu_245_p1}, {bitcast_ln94_20_fu_237_p1}}, {bitcast_ln94_19_fu_229_p1}}, {bitcast_ln94_fu_221_p1}};

assign select_ln97_fu_274_p3 = ((icmp_ln97_fu_268_p2[0:0] == 1'b1) ? 16'd0 : add_ln96_fu_262_p2);

assign shl_ln89_fu_140_p2 = add_ln94_fu_134_p2 << 16'd2;

assign sub_ln94_cast14_fu_127_p1 = sub_ln94_reg_294;

assign sub_ln94_fu_121_p2 = (zext_ln94_fu_105_p1 - zext_ln94_15_fu_117_p1);

assign tmp_fu_97_p3 = {{i}, {7'd0}};

assign tmp_s_fu_109_p3 = {{i}, {4'd0}};

assign trunc_ln86_fu_154_p1 = outputCount_1[1:0];

assign trunc_ln94_fu_202_p1 = outputChanIdx_1[3:0];

assign zext_ln94_15_fu_117_p1 = tmp_s_fu_109_p3;

assign zext_ln94_16_fu_130_p1 = j;

assign zext_ln94_17_fu_206_p1 = trunc_ln94_fu_202_p1;

assign zext_ln94_18_fu_216_p1 = add_ln94_7_fu_210_p2;

assign zext_ln94_fu_105_p1 = tmp_fu_97_p3;

always @ (posedge ap_clk) begin
    sub_ln94_reg_294[3:0] <= 4'b0000;
end

endmodule //td_fused_top_tdf1_writeOutputs_unaligned
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf2_113 (
        in_data_address0,
        in_data_ce0,
        in_data_d0,
        in_data_q0,
        in_data_we0,
        in_data_address1,
        in_data_ce1,
        in_data_d1,
        in_data_q1,
        in_data_we1,
        out_data_address0,
        out_data_ce0,
        out_data_d0,
        out_data_q0,
        out_data_we0,
        out_data_address1,
        out_data_ce1,
        out_data_d1,
        out_data_q1,
        out_data_we1,
        filter_data_address0,
        filter_data_ce0,
        filter_data_d0,
        filter_data_q0,
        filter_data_we0,
        filter_data_address1,
        filter_data_ce1,
        filter_data_d1,
        filter_data_q1,
        filter_data_we1,
        adjustments_address0,
        adjustments_ce0,
        adjustments_d0,
        adjustments_q0,
        adjustments_we0,
        adjustments_address1,
        adjustments_ce1,
        adjustments_d1,
        adjustments_q1,
        adjustments_we1,
        ap_clk,
        ap_rst,
        in_data_empty_n,
        in_data_read,
        out_data_full_n,
        out_data_write,
        ap_start,
        ap_done,
        ap_ready,
        ap_idle,
        ap_continue
);


output  [15:0] in_data_address0;
output   in_data_ce0;
output  [63:0] in_data_d0;
input  [63:0] in_data_q0;
output   in_data_we0;
output  [15:0] in_data_address1;
output   in_data_ce1;
output  [63:0] in_data_d1;
input  [63:0] in_data_q1;
output   in_data_we1;
output  [14:0] out_data_address0;
output   out_data_ce0;
output  [63:0] out_data_d0;
input  [63:0] out_data_q0;
output   out_data_we0;
output  [14:0] out_data_address1;
output   out_data_ce1;
output  [63:0] out_data_d1;
input  [63:0] out_data_q1;
output   out_data_we1;
output  [12:0] filter_data_address0;
output   filter_data_ce0;
output  [15:0] filter_data_d0;
input  [15:0] filter_data_q0;
output   filter_data_we0;
output  [12:0] filter_data_address1;
output   filter_data_ce1;
output  [15:0] filter_data_d1;
input  [15:0] filter_data_q1;
output   filter_data_we1;
output  [4:0] adjustments_address0;
output   adjustments_ce0;
output  [47:0] adjustments_d0;
input  [47:0] adjustments_q0;
output   adjustments_we0;
output  [4:0] adjustments_address1;
output   adjustments_ce1;
output  [47:0] adjustments_d1;
input  [47:0] adjustments_q1;
output   adjustments_we1;
input   ap_clk;
input   ap_rst;
input   in_data_empty_n;
output   in_data_read;
input   out_data_full_n;
output   out_data_write;
input   ap_start;
output   ap_done;
output   ap_ready;
output   ap_idle;
input   ap_continue;

reg ap_done;
reg ap_ready;
reg ap_idle;

wire   [15:0] dataflow_in_loop_TOP_LOOP38022_U0_in_data_address0;
wire    dataflow_in_loop_TOP_LOOP38022_U0_in_data_ce0;
wire   [63:0] dataflow_in_loop_TOP_LOOP38022_U0_in_data_d0;
wire    dataflow_in_loop_TOP_LOOP38022_U0_in_data_we0;
wire   [15:0] dataflow_in_loop_TOP_LOOP38022_U0_in_data_address1;
wire    dataflow_in_loop_TOP_LOOP38022_U0_in_data_ce1;
wire   [63:0] dataflow_in_loop_TOP_LOOP38022_U0_in_data_d1;
wire    dataflow_in_loop_TOP_LOOP38022_U0_in_data_we1;
wire   [12:0] dataflow_in_loop_TOP_LOOP38022_U0_filter_data_address0;
wire    dataflow_in_loop_TOP_LOOP38022_U0_filter_data_ce0;
wire   [15:0] dataflow_in_loop_TOP_LOOP38022_U0_filter_data_d0;
wire    dataflow_in_loop_TOP_LOOP38022_U0_filter_data_we0;
wire   [12:0] dataflow_in_loop_TOP_LOOP38022_U0_filter_data_address1;
wire    dataflow_in_loop_TOP_LOOP38022_U0_filter_data_ce1;
wire   [15:0] dataflow_in_loop_TOP_LOOP38022_U0_filter_data_d1;
wire    dataflow_in_loop_TOP_LOOP38022_U0_filter_data_we1;
wire   [4:0] dataflow_in_loop_TOP_LOOP38022_U0_adjustments_address0;
wire    dataflow_in_loop_TOP_LOOP38022_U0_adjustments_ce0;
wire   [47:0] dataflow_in_loop_TOP_LOOP38022_U0_adjustments_d0;
wire    dataflow_in_loop_TOP_LOOP38022_U0_adjustments_we0;
wire   [4:0] dataflow_in_loop_TOP_LOOP38022_U0_adjustments_address1;
wire    dataflow_in_loop_TOP_LOOP38022_U0_adjustments_ce1;
wire   [47:0] dataflow_in_loop_TOP_LOOP38022_U0_adjustments_d1;
wire    dataflow_in_loop_TOP_LOOP38022_U0_adjustments_we1;
wire   [14:0] dataflow_in_loop_TOP_LOOP38022_U0_out_data_address0;
wire    dataflow_in_loop_TOP_LOOP38022_U0_out_data_ce0;
wire   [63:0] dataflow_in_loop_TOP_LOOP38022_U0_out_data_d0;
wire    dataflow_in_loop_TOP_LOOP38022_U0_out_data_we0;
wire   [14:0] dataflow_in_loop_TOP_LOOP38022_U0_out_data_address1;
wire    dataflow_in_loop_TOP_LOOP38022_U0_out_data_ce1;
wire   [63:0] dataflow_in_loop_TOP_LOOP38022_U0_out_data_d1;
wire    dataflow_in_loop_TOP_LOOP38022_U0_out_data_we1;
wire    dataflow_in_loop_TOP_LOOP38022_U0_ap_start;
wire    dataflow_in_loop_TOP_LOOP38022_U0_in_data_read;
wire    dataflow_in_loop_TOP_LOOP38022_U0_out_data_write;
wire    dataflow_in_loop_TOP_LOOP38022_U0_ap_done;
wire    dataflow_in_loop_TOP_LOOP38022_U0_ap_ready;
wire    dataflow_in_loop_TOP_LOOP38022_U0_ap_idle;
reg    dataflow_in_loop_TOP_LOOP38022_U0_ap_continue;
wire    dataflow_in_loop_TOP_LOOP38022_U0_in_data_full_n;
wire    dataflow_in_loop_TOP_LOOP38022_U0_in_data_write;
wire    ap_sync_continue;
wire    ap_sync_done;
wire    ap_sync_ready;
reg   [18:0] loop_dataflow_input_count;
reg   [18:0] loop_dataflow_output_count;
wire   [18:0] bound_minus_1;
wire    dataflow_in_loop_TOP_LOOP38022_U0_start_full_n;
wire    dataflow_in_loop_TOP_LOOP38022_U0_start_write;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 loop_dataflow_input_count = 19'd0;
#0 loop_dataflow_output_count = 19'd0;
end

td_fused_top_dataflow_in_loop_TOP_LOOP38022 dataflow_in_loop_TOP_LOOP38022_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .in_data_address0(dataflow_in_loop_TOP_LOOP38022_U0_in_data_address0),
    .in_data_ce0(dataflow_in_loop_TOP_LOOP38022_U0_in_data_ce0),
    .in_data_d0(dataflow_in_loop_TOP_LOOP38022_U0_in_data_d0),
    .in_data_q0(in_data_q0),
    .in_data_we0(dataflow_in_loop_TOP_LOOP38022_U0_in_data_we0),
    .in_data_address1(dataflow_in_loop_TOP_LOOP38022_U0_in_data_address1),
    .in_data_ce1(dataflow_in_loop_TOP_LOOP38022_U0_in_data_ce1),
    .in_data_d1(dataflow_in_loop_TOP_LOOP38022_U0_in_data_d1),
    .in_data_q1(64'd0),
    .in_data_we1(dataflow_in_loop_TOP_LOOP38022_U0_in_data_we1),
    .filter_data_address0(dataflow_in_loop_TOP_LOOP38022_U0_filter_data_address0),
    .filter_data_ce0(dataflow_in_loop_TOP_LOOP38022_U0_filter_data_ce0),
    .filter_data_d0(dataflow_in_loop_TOP_LOOP38022_U0_filter_data_d0),
    .filter_data_q0(filter_data_q0),
    .filter_data_we0(dataflow_in_loop_TOP_LOOP38022_U0_filter_data_we0),
    .filter_data_address1(dataflow_in_loop_TOP_LOOP38022_U0_filter_data_address1),
    .filter_data_ce1(dataflow_in_loop_TOP_LOOP38022_U0_filter_data_ce1),
    .filter_data_d1(dataflow_in_loop_TOP_LOOP38022_U0_filter_data_d1),
    .filter_data_q1(16'd0),
    .filter_data_we1(dataflow_in_loop_TOP_LOOP38022_U0_filter_data_we1),
    .adjustments_address0(dataflow_in_loop_TOP_LOOP38022_U0_adjustments_address0),
    .adjustments_ce0(dataflow_in_loop_TOP_LOOP38022_U0_adjustments_ce0),
    .adjustments_d0(dataflow_in_loop_TOP_LOOP38022_U0_adjustments_d0),
    .adjustments_q0(adjustments_q0),
    .adjustments_we0(dataflow_in_loop_TOP_LOOP38022_U0_adjustments_we0),
    .adjustments_address1(dataflow_in_loop_TOP_LOOP38022_U0_adjustments_address1),
    .adjustments_ce1(dataflow_in_loop_TOP_LOOP38022_U0_adjustments_ce1),
    .adjustments_d1(dataflow_in_loop_TOP_LOOP38022_U0_adjustments_d1),
    .adjustments_q1(48'd0),
    .adjustments_we1(dataflow_in_loop_TOP_LOOP38022_U0_adjustments_we1),
    .out_data_address0(dataflow_in_loop_TOP_LOOP38022_U0_out_data_address0),
    .out_data_ce0(dataflow_in_loop_TOP_LOOP38022_U0_out_data_ce0),
    .out_data_d0(dataflow_in_loop_TOP_LOOP38022_U0_out_data_d0),
    .out_data_q0(64'd0),
    .out_data_we0(dataflow_in_loop_TOP_LOOP38022_U0_out_data_we0),
    .out_data_address1(dataflow_in_loop_TOP_LOOP38022_U0_out_data_address1),
    .out_data_ce1(dataflow_in_loop_TOP_LOOP38022_U0_out_data_ce1),
    .out_data_d1(dataflow_in_loop_TOP_LOOP38022_U0_out_data_d1),
    .out_data_q1(64'd0),
    .out_data_we1(dataflow_in_loop_TOP_LOOP38022_U0_out_data_we1),
    .ap_start(dataflow_in_loop_TOP_LOOP38022_U0_ap_start),
    .in_data_empty_n(1'b0),
    .in_data_read(dataflow_in_loop_TOP_LOOP38022_U0_in_data_read),
    .out_data_full_n(out_data_full_n),
    .out_data_write(dataflow_in_loop_TOP_LOOP38022_U0_out_data_write),
    .ap_done(dataflow_in_loop_TOP_LOOP38022_U0_ap_done),
    .ap_ready(dataflow_in_loop_TOP_LOOP38022_U0_ap_ready),
    .ap_idle(dataflow_in_loop_TOP_LOOP38022_U0_ap_idle),
    .ap_continue(dataflow_in_loop_TOP_LOOP38022_U0_ap_continue)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        loop_dataflow_input_count <= 19'd0;
    end else begin
        if ((~(loop_dataflow_input_count == bound_minus_1) & (dataflow_in_loop_TOP_LOOP38022_U0_ap_ready == 1'b1) & (ap_start == 1'b1))) begin
            loop_dataflow_input_count <= (loop_dataflow_input_count + 19'd1);
        end else if (((dataflow_in_loop_TOP_LOOP38022_U0_ap_ready == 1'b1) & (loop_dataflow_input_count == bound_minus_1) & (ap_start == 1'b1))) begin
            loop_dataflow_input_count <= 19'd0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        loop_dataflow_output_count <= 19'd0;
    end else begin
        if ((~(loop_dataflow_output_count == bound_minus_1) & (dataflow_in_loop_TOP_LOOP38022_U0_ap_continue == 1'b1) & (dataflow_in_loop_TOP_LOOP38022_U0_ap_done == 1'b1))) begin
            loop_dataflow_output_count <= (loop_dataflow_output_count + 19'd1);
        end else if (((dataflow_in_loop_TOP_LOOP38022_U0_ap_continue == 1'b1) & (dataflow_in_loop_TOP_LOOP38022_U0_ap_done == 1'b1) & (loop_dataflow_output_count == bound_minus_1))) begin
            loop_dataflow_output_count <= 19'd0;
        end
    end
end

always @ (*) begin
    if (((dataflow_in_loop_TOP_LOOP38022_U0_ap_done == 1'b1) & (loop_dataflow_output_count == bound_minus_1))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = 1'b0;
    end
end

always @ (*) begin
    if (((dataflow_in_loop_TOP_LOOP38022_U0_ap_idle == 1'b1) & (loop_dataflow_output_count == 19'd0) & (ap_start == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((dataflow_in_loop_TOP_LOOP38022_U0_ap_ready == 1'b1) & (loop_dataflow_input_count == bound_minus_1) & (ap_start == 1'b1))) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((~(loop_dataflow_output_count == bound_minus_1) | (ap_continue == 1'b1))) begin
        dataflow_in_loop_TOP_LOOP38022_U0_ap_continue = 1'b1;
    end else begin
        dataflow_in_loop_TOP_LOOP38022_U0_ap_continue = 1'b0;
    end
end

assign adjustments_address0 = dataflow_in_loop_TOP_LOOP38022_U0_adjustments_address0;

assign adjustments_address1 = 5'd0;

assign adjustments_ce0 = dataflow_in_loop_TOP_LOOP38022_U0_adjustments_ce0;

assign adjustments_ce1 = 1'b0;

assign adjustments_d0 = 48'd0;

assign adjustments_d1 = 48'd0;

assign adjustments_we0 = 1'b0;

assign adjustments_we1 = 1'b0;

assign ap_sync_continue = ap_continue;

assign ap_sync_done = dataflow_in_loop_TOP_LOOP38022_U0_ap_done;

assign ap_sync_ready = dataflow_in_loop_TOP_LOOP38022_U0_ap_ready;

assign bound_minus_1 = (19'd401408 - 19'd1);

assign dataflow_in_loop_TOP_LOOP38022_U0_ap_start = ap_start;

assign dataflow_in_loop_TOP_LOOP38022_U0_in_data_full_n = in_data_empty_n;

assign dataflow_in_loop_TOP_LOOP38022_U0_in_data_write = 1'b0;

assign dataflow_in_loop_TOP_LOOP38022_U0_start_full_n = 1'b1;

assign dataflow_in_loop_TOP_LOOP38022_U0_start_write = 1'b0;

assign filter_data_address0 = dataflow_in_loop_TOP_LOOP38022_U0_filter_data_address0;

assign filter_data_address1 = 13'd0;

assign filter_data_ce0 = dataflow_in_loop_TOP_LOOP38022_U0_filter_data_ce0;

assign filter_data_ce1 = 1'b0;

assign filter_data_d0 = 16'd0;

assign filter_data_d1 = 16'd0;

assign filter_data_we0 = 1'b0;

assign filter_data_we1 = 1'b0;

assign in_data_address0 = dataflow_in_loop_TOP_LOOP38022_U0_in_data_address0;

assign in_data_address1 = 16'd0;

assign in_data_ce0 = dataflow_in_loop_TOP_LOOP38022_U0_in_data_ce0;

assign in_data_ce1 = 1'b0;

assign in_data_d0 = 64'd0;

assign in_data_d1 = 64'd0;

assign in_data_read = dataflow_in_loop_TOP_LOOP38022_U0_in_data_write;

assign in_data_we0 = 1'b0;

assign in_data_we1 = 1'b0;

assign out_data_address0 = 15'd0;

assign out_data_address1 = dataflow_in_loop_TOP_LOOP38022_U0_out_data_address1;

assign out_data_ce0 = 1'b0;

assign out_data_ce1 = dataflow_in_loop_TOP_LOOP38022_U0_out_data_ce1;

assign out_data_d0 = 64'd0;

assign out_data_d1 = dataflow_in_loop_TOP_LOOP38022_U0_out_data_d1;

assign out_data_we0 = 1'b0;

assign out_data_we1 = dataflow_in_loop_TOP_LOOP38022_U0_out_data_we1;

assign out_data_write = dataflow_in_loop_TOP_LOOP38022_U0_out_data_write;

endmodule //td_fused_top_tdf2_113
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf2_accum_1 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        accum_in_0_address0,
        accum_in_0_ce0,
        accum_in_0_q0,
        accum_in_0_address1,
        accum_in_0_ce1,
        accum_in_0_q1,
        accum_out_address0,
        accum_out_ce0,
        accum_out_we0,
        accum_out_d0,
        accum_out_address1,
        accum_out_ce1,
        accum_out_we1,
        accum_out_d1
);

parameter    ap_ST_fsm_state1 = 8'd1;
parameter    ap_ST_fsm_pp0_stage0 = 8'd2;
parameter    ap_ST_fsm_pp0_stage1 = 8'd4;
parameter    ap_ST_fsm_pp0_stage2 = 8'd8;
parameter    ap_ST_fsm_pp0_stage3 = 8'd16;
parameter    ap_ST_fsm_state12 = 8'd32;
parameter    ap_ST_fsm_state13 = 8'd64;
parameter    ap_ST_fsm_state14 = 8'd128;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [7:0] accum_in_0_address0;
output   accum_in_0_ce0;
input  [15:0] accum_in_0_q0;
output  [7:0] accum_in_0_address1;
output   accum_in_0_ce1;
input  [15:0] accum_in_0_q1;
output  [2:0] accum_out_address0;
output   accum_out_ce0;
output   accum_out_we0;
output  [15:0] accum_out_d0;
output  [2:0] accum_out_address1;
output   accum_out_ce1;
output   accum_out_we1;
output  [15:0] accum_out_d1;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg[7:0] accum_in_0_address0;
reg accum_in_0_ce0;
reg[7:0] accum_in_0_address1;
reg accum_in_0_ce1;
reg accum_out_ce0;
reg accum_out_we0;
reg accum_out_ce1;
reg accum_out_we1;

reg    ap_done_reg;
  reg   [7:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg   [7:0] x_reg_168;
reg   [15:0] psum_7_08_reg_180;
reg   [15:0] psum_6_07_reg_192;
reg   [15:0] psum_5_06_reg_204;
reg   [15:0] psum_4_05_reg_216;
reg   [15:0] psum_3_04_reg_228;
reg   [15:0] psum_2_03_reg_240;
reg   [15:0] psum_1_02_reg_252;
reg   [15:0] psum_0_01_reg_264;
wire   [0:0] icmp_ln49_fu_321_p2;
reg   [0:0] icmp_ln49_reg_492;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state6_pp0_stage0_iter1;
wire    ap_block_state10_pp0_stage0_iter2;
wire    ap_block_pp0_stage0_11001;
reg   [0:0] icmp_ln49_reg_492_pp0_iter1_reg;
reg   [0:0] icmp_ln49_reg_492_pp0_iter2_reg;
reg   [15:0] accum_in_0_load_reg_506;
wire    ap_CS_fsm_pp0_stage1;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_state3_pp0_stage1_iter0;
wire    ap_block_state7_pp0_stage1_iter1;
wire    ap_block_state11_pp0_stage1_iter2;
wire    ap_block_pp0_stage1_11001;
reg   [15:0] accum_in_0_load_50_reg_511;
reg   [15:0] accum_in_0_load_51_reg_526;
wire    ap_CS_fsm_pp0_stage2;
wire    ap_block_state4_pp0_stage2_iter0;
wire    ap_block_state8_pp0_stage2_iter1;
wire    ap_block_pp0_stage2_11001;
reg   [15:0] accum_in_0_load_52_reg_531;
wire   [7:0] add_ln49_fu_387_p2;
reg   [7:0] add_ln49_reg_546;
wire    ap_CS_fsm_pp0_stage3;
wire    ap_block_state5_pp0_stage3_iter0;
wire    ap_block_state9_pp0_stage3_iter1;
wire    ap_block_pp0_stage3_11001;
reg   [15:0] accum_in_0_load_53_reg_551;
reg   [15:0] accum_in_0_load_54_reg_556;
reg   [15:0] accum_in_0_load_55_reg_571;
reg    ap_enable_reg_pp0_iter1;
reg   [15:0] accum_in_0_load_56_reg_576;
wire   [15:0] grp_fu_305_p2;
wire   [15:0] grp_fu_310_p2;
reg    ap_enable_reg_pp0_iter2;
wire   [3:0] add_ln57_fu_432_p2;
wire    ap_CS_fsm_state13;
wire   [0:0] tmp_fu_415_p3;
reg    ap_block_state1;
wire    ap_block_pp0_stage2_subdone;
reg    ap_condition_pp0_exit_iter0_state4;
wire    ap_block_pp0_stage3_subdone;
wire    ap_block_pp0_stage1_subdone;
reg   [7:0] ap_phi_mux_x_phi_fu_172_p4;
wire    ap_block_pp0_stage0;
wire   [15:0] ap_phi_mux_psum_7_08_phi_fu_184_p4;
wire    ap_block_pp0_stage1;
wire   [15:0] ap_phi_mux_psum_6_07_phi_fu_196_p4;
wire   [15:0] ap_phi_mux_psum_5_06_phi_fu_208_p4;
wire   [15:0] ap_phi_mux_psum_4_05_phi_fu_220_p4;
wire   [15:0] ap_phi_mux_psum_3_04_phi_fu_232_p4;
wire    ap_block_pp0_stage3;
wire   [15:0] ap_phi_mux_psum_2_03_phi_fu_244_p4;
wire    ap_block_pp0_stage2;
reg   [3:0] q_reg_276;
wire    ap_CS_fsm_state12;
reg   [15:0] ap_phi_mux_phi_ln69_phi_fu_290_p8;
wire   [2:0] trunc_ln57_fu_428_p1;
wire   [63:0] zext_ln49_fu_327_p1;
wire   [63:0] zext_ln53_fu_338_p1;
wire   [63:0] zext_ln53_13_fu_349_p1;
wire   [63:0] zext_ln53_14_fu_360_p1;
wire   [63:0] zext_ln53_15_fu_371_p1;
wire   [63:0] zext_ln53_16_fu_382_p1;
wire   [63:0] zext_ln53_17_fu_399_p1;
wire   [63:0] zext_ln53_18_fu_410_p1;
wire   [63:0] zext_ln57_fu_423_p1;
wire   [63:0] zext_ln57_3_fu_444_p1;
reg   [15:0] grp_fu_305_p0;
reg   [15:0] grp_fu_305_p1;
reg   [15:0] grp_fu_310_p0;
reg   [15:0] grp_fu_310_p1;
wire   [7:0] or_ln53_fu_332_p2;
wire   [7:0] or_ln53_13_fu_343_p2;
wire   [7:0] or_ln53_14_fu_354_p2;
wire   [7:0] or_ln53_15_fu_365_p2;
wire   [7:0] or_ln53_16_fu_376_p2;
wire   [7:0] or_ln53_17_fu_393_p2;
wire   [7:0] or_ln53_18_fu_404_p2;
wire   [2:0] or_ln57_fu_438_p2;
wire   [0:0] icmp_ln69_fu_449_p2;
wire   [0:0] icmp_ln69_5_fu_463_p2;
wire   [15:0] select_ln69_fu_455_p3;
wire   [0:0] icmp_ln69_6_fu_477_p2;
wire   [15:0] select_ln69_5_fu_469_p3;
wire    ap_CS_fsm_state14;
reg   [7:0] ap_NS_fsm;
wire    ap_block_pp0_stage0_subdone;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
reg    ap_condition_514;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 8'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
end

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U96(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(grp_fu_305_p0),
    .din1(grp_fu_305_p1),
    .dout(grp_fu_305_p2)
);

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U97(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(grp_fu_310_p0),
    .din1(grp_fu_310_p1),
    .dout(grp_fu_310_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state14)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage2_subdone) & (1'b1 == ap_condition_pp0_exit_iter0_state4) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage3_subdone) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b0)) | ((1'b0 == ap_block_pp0_stage3_subdone) & (1'b1 == ap_CS_fsm_pp0_stage3)))) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end else if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter2 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state12)) begin
        q_reg_276 <= 4'd0;
    end else if (((tmp_fu_415_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state13))) begin
        q_reg_276 <= add_ln57_fu_432_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln49_reg_492 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        x_reg_168 <= add_ln49_reg_546;
    end else if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        x_reg_168 <= 8'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage1_11001) & (icmp_ln49_reg_492 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
        accum_in_0_load_50_reg_511 <= accum_in_0_q0;
        accum_in_0_load_reg_506 <= accum_in_0_q1;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2_11001) & (icmp_ln49_reg_492 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
        accum_in_0_load_51_reg_526 <= accum_in_0_q1;
        accum_in_0_load_52_reg_531 <= accum_in_0_q0;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage3_11001) & (icmp_ln49_reg_492 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
        accum_in_0_load_53_reg_551 <= accum_in_0_q1;
        accum_in_0_load_54_reg_556 <= accum_in_0_q0;
        add_ln49_reg_546 <= add_ln49_fu_387_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln49_reg_492 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        accum_in_0_load_55_reg_571 <= accum_in_0_q1;
        accum_in_0_load_56_reg_576 <= accum_in_0_q0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln49_reg_492 <= icmp_ln49_fu_321_p2;
        icmp_ln49_reg_492_pp0_iter1_reg <= icmp_ln49_reg_492;
        icmp_ln49_reg_492_pp0_iter2_reg <= icmp_ln49_reg_492_pp0_iter1_reg;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln49_reg_492_pp0_iter1_reg == 1'd1) & (1'b0 == ap_block_pp0_stage2_11001) & (1'b1 == ap_CS_fsm_pp0_stage2) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        psum_0_01_reg_264 <= grp_fu_305_p2;
        psum_1_02_reg_252 <= grp_fu_310_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln49_reg_492_pp0_iter1_reg == 1'd1) & (1'b0 == ap_block_pp0_stage3_11001) & (1'b1 == ap_CS_fsm_pp0_stage3) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        psum_2_03_reg_240 <= grp_fu_305_p2;
        psum_3_04_reg_228 <= grp_fu_310_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln49_reg_492_pp0_iter1_reg == 1'd1) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        psum_4_05_reg_216 <= grp_fu_305_p2;
        psum_5_06_reg_204 <= grp_fu_310_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln49_reg_492_pp0_iter2_reg == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        psum_6_07_reg_192 <= grp_fu_305_p2;
        psum_7_08_reg_180 <= grp_fu_310_p2;
    end
end

always @ (*) begin
    if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
        if (((1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            accum_in_0_address0 = zext_ln53_18_fu_410_p1;
        end else if (((1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            accum_in_0_address0 = zext_ln53_16_fu_382_p1;
        end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            accum_in_0_address0 = zext_ln53_14_fu_360_p1;
        end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            accum_in_0_address0 = zext_ln53_fu_338_p1;
        end else begin
            accum_in_0_address0 = 'bx;
        end
    end else begin
        accum_in_0_address0 = 'bx;
    end
end

always @ (*) begin
    if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
        if (((1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            accum_in_0_address1 = zext_ln53_17_fu_399_p1;
        end else if (((1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            accum_in_0_address1 = zext_ln53_15_fu_371_p1;
        end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            accum_in_0_address1 = zext_ln53_13_fu_349_p1;
        end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            accum_in_0_address1 = zext_ln49_fu_327_p1;
        end else begin
            accum_in_0_address1 = 'bx;
        end
    end else begin
        accum_in_0_address1 = 'bx;
    end
end

always @ (*) begin
    if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage3_11001) & (1'b1 == ap_CS_fsm_pp0_stage3)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2_11001) & (1'b1 == ap_CS_fsm_pp0_stage2)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1)))) begin
        accum_in_0_ce0 = 1'b1;
    end else begin
        accum_in_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage3_11001) & (1'b1 == ap_CS_fsm_pp0_stage3)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2_11001) & (1'b1 == ap_CS_fsm_pp0_stage2)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1)))) begin
        accum_in_0_ce1 = 1'b1;
    end else begin
        accum_in_0_ce1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state13)) begin
        accum_out_ce0 = 1'b1;
    end else begin
        accum_out_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state13)) begin
        accum_out_ce1 = 1'b1;
    end else begin
        accum_out_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((tmp_fu_415_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state13))) begin
        accum_out_we0 = 1'b1;
    end else begin
        accum_out_we0 = 1'b0;
    end
end

always @ (*) begin
    if (((tmp_fu_415_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state13))) begin
        accum_out_we1 = 1'b1;
    end else begin
        accum_out_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((icmp_ln49_reg_492 == 1'd0)) begin
        ap_condition_pp0_exit_iter0_state4 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state4 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state14)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((tmp_fu_415_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state13))) begin
        if ((trunc_ln57_fu_428_p1 == 3'd0)) begin
            ap_phi_mux_phi_ln69_phi_fu_290_p8 = psum_0_01_reg_264;
        end else if ((1'b1 == ap_condition_514)) begin
            ap_phi_mux_phi_ln69_phi_fu_290_p8 = psum_6_07_reg_192;
        end else if ((trunc_ln57_fu_428_p1 == 3'd4)) begin
            ap_phi_mux_phi_ln69_phi_fu_290_p8 = psum_4_05_reg_216;
        end else if ((trunc_ln57_fu_428_p1 == 3'd2)) begin
            ap_phi_mux_phi_ln69_phi_fu_290_p8 = psum_2_03_reg_240;
        end else begin
            ap_phi_mux_phi_ln69_phi_fu_290_p8 = 'bx;
        end
    end else begin
        ap_phi_mux_phi_ln69_phi_fu_290_p8 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0) & (icmp_ln49_reg_492 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_x_phi_fu_172_p4 = add_ln49_reg_546;
    end else begin
        ap_phi_mux_x_phi_fu_172_p4 = x_reg_168;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state14)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_305_p0 = ap_phi_mux_psum_6_07_phi_fu_196_p4;
    end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_305_p0 = ap_phi_mux_psum_4_05_phi_fu_220_p4;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
        grp_fu_305_p0 = ap_phi_mux_psum_2_03_phi_fu_244_p4;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
        grp_fu_305_p0 = grp_fu_305_p2;
    end else begin
        grp_fu_305_p0 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_305_p1 = accum_in_0_load_55_reg_571;
    end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_305_p1 = accum_in_0_load_53_reg_551;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
        grp_fu_305_p1 = accum_in_0_load_51_reg_526;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
        grp_fu_305_p1 = accum_in_0_load_reg_506;
    end else begin
        grp_fu_305_p1 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_310_p0 = ap_phi_mux_psum_7_08_phi_fu_184_p4;
    end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_310_p0 = ap_phi_mux_psum_5_06_phi_fu_208_p4;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
        grp_fu_310_p0 = ap_phi_mux_psum_3_04_phi_fu_232_p4;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
        grp_fu_310_p0 = grp_fu_310_p2;
    end else begin
        grp_fu_310_p0 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_310_p1 = accum_in_0_load_56_reg_576;
    end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_310_p1 = accum_in_0_load_54_reg_556;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
        grp_fu_310_p1 = accum_in_0_load_52_reg_531;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
        grp_fu_310_p1 = accum_in_0_load_50_reg_511;
    end else begin
        grp_fu_310_p1 = 'bx;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_pp0_stage1 : begin
            if ((~((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter2 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0)) & (1'b0 == ap_block_pp0_stage1_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage2;
            end else if (((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter2 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
                ap_NS_fsm = ap_ST_fsm_state12;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end
        end
        ap_ST_fsm_pp0_stage2 : begin
            if ((~((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2_subdone) & (icmp_ln49_reg_492 == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b0)) & (1'b0 == ap_block_pp0_stage2_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage3;
            end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2_subdone) & (icmp_ln49_reg_492 == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
                ap_NS_fsm = ap_ST_fsm_state12;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage2;
            end
        end
        ap_ST_fsm_pp0_stage3 : begin
            if ((1'b0 == ap_block_pp0_stage3_subdone)) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage3;
            end
        end
        ap_ST_fsm_state12 : begin
            ap_NS_fsm = ap_ST_fsm_state13;
        end
        ap_ST_fsm_state13 : begin
            if (((tmp_fu_415_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state13))) begin
                ap_NS_fsm = ap_ST_fsm_state13;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state14;
            end
        end
        ap_ST_fsm_state14 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign accum_out_address0 = zext_ln57_3_fu_444_p1;

assign accum_out_address1 = zext_ln57_fu_423_p1;

assign accum_out_d0 = ((icmp_ln69_6_fu_477_p2[0:0] == 1'b1) ? psum_5_06_reg_204 : select_ln69_5_fu_469_p3);

assign accum_out_d1 = ap_phi_mux_phi_ln69_phi_fu_290_p8;

assign add_ln49_fu_387_p2 = (x_reg_168 + 8'd8);

assign add_ln57_fu_432_p2 = (q_reg_276 + 4'd2);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_pp0_stage1 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_pp0_stage2 = ap_CS_fsm[32'd3];

assign ap_CS_fsm_pp0_stage3 = ap_CS_fsm[32'd4];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state12 = ap_CS_fsm[32'd5];

assign ap_CS_fsm_state13 = ap_CS_fsm[32'd6];

assign ap_CS_fsm_state14 = ap_CS_fsm[32'd7];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1_subdone = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage2 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage2_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage2_subdone = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage3 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage3_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage3_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((ap_done_reg == 1'b1) | (ap_start == 1'b0));
end

assign ap_block_state10_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state11_pp0_stage1_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage1_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage2_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage3_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage1_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage2_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state9_pp0_stage3_iter1 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_condition_514 = (~(trunc_ln57_fu_428_p1 == 3'd0) & ~(trunc_ln57_fu_428_p1 == 3'd4) & ~(trunc_ln57_fu_428_p1 == 3'd2));
end

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign ap_phi_mux_psum_2_03_phi_fu_244_p4 = grp_fu_305_p2;

assign ap_phi_mux_psum_3_04_phi_fu_232_p4 = grp_fu_310_p2;

assign ap_phi_mux_psum_4_05_phi_fu_220_p4 = grp_fu_305_p2;

assign ap_phi_mux_psum_5_06_phi_fu_208_p4 = grp_fu_310_p2;

assign ap_phi_mux_psum_6_07_phi_fu_196_p4 = grp_fu_305_p2;

assign ap_phi_mux_psum_7_08_phi_fu_184_p4 = grp_fu_310_p2;

assign icmp_ln49_fu_321_p2 = ((ap_phi_mux_x_phi_fu_172_p4 < 8'd144) ? 1'b1 : 1'b0);

assign icmp_ln69_5_fu_463_p2 = ((or_ln57_fu_438_p2 == 3'd3) ? 1'b1 : 1'b0);

assign icmp_ln69_6_fu_477_p2 = ((or_ln57_fu_438_p2 == 3'd5) ? 1'b1 : 1'b0);

assign icmp_ln69_fu_449_p2 = ((or_ln57_fu_438_p2 == 3'd1) ? 1'b1 : 1'b0);

assign or_ln53_13_fu_343_p2 = (x_reg_168 | 8'd2);

assign or_ln53_14_fu_354_p2 = (x_reg_168 | 8'd3);

assign or_ln53_15_fu_365_p2 = (x_reg_168 | 8'd4);

assign or_ln53_16_fu_376_p2 = (x_reg_168 | 8'd5);

assign or_ln53_17_fu_393_p2 = (x_reg_168 | 8'd6);

assign or_ln53_18_fu_404_p2 = (x_reg_168 | 8'd7);

assign or_ln53_fu_332_p2 = (ap_phi_mux_x_phi_fu_172_p4 | 8'd1);

assign or_ln57_fu_438_p2 = (trunc_ln57_fu_428_p1 | 3'd1);

assign select_ln69_5_fu_469_p3 = ((icmp_ln69_5_fu_463_p2[0:0] == 1'b1) ? psum_3_04_reg_228 : select_ln69_fu_455_p3);

assign select_ln69_fu_455_p3 = ((icmp_ln69_fu_449_p2[0:0] == 1'b1) ? psum_1_02_reg_252 : psum_7_08_reg_180);

assign tmp_fu_415_p3 = q_reg_276[32'd3];

assign trunc_ln57_fu_428_p1 = q_reg_276[2:0];

assign zext_ln49_fu_327_p1 = ap_phi_mux_x_phi_fu_172_p4;

assign zext_ln53_13_fu_349_p1 = or_ln53_13_fu_343_p2;

assign zext_ln53_14_fu_360_p1 = or_ln53_14_fu_354_p2;

assign zext_ln53_15_fu_371_p1 = or_ln53_15_fu_365_p2;

assign zext_ln53_16_fu_382_p1 = or_ln53_16_fu_376_p2;

assign zext_ln53_17_fu_399_p1 = or_ln53_17_fu_393_p2;

assign zext_ln53_18_fu_410_p1 = or_ln53_18_fu_404_p2;

assign zext_ln53_fu_338_p1 = or_ln53_fu_332_p2;

assign zext_ln57_3_fu_444_p1 = or_ln57_fu_438_p2;

assign zext_ln57_fu_423_p1 = q_reg_276;

endmodule //td_fused_top_tdf2_accum_1
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf2_accum_2 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        accum_in_16,
        accum_in_16_ap_vld,
        accum_in_address0,
        accum_in_ce0,
        accum_in_q0
);

parameter    ap_ST_fsm_state1 = 7'd1;
parameter    ap_ST_fsm_state2 = 7'd2;
parameter    ap_ST_fsm_state3 = 7'd4;
parameter    ap_ST_fsm_state4 = 7'd8;
parameter    ap_ST_fsm_state5 = 7'd16;
parameter    ap_ST_fsm_state6 = 7'd32;
parameter    ap_ST_fsm_state7 = 7'd64;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [15:0] accum_in_16;
output   accum_in_16_ap_vld;
output  [2:0] accum_in_address0;
output   accum_in_ce0;
input  [15:0] accum_in_q0;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg[15:0] accum_in_16;
reg accum_in_16_ap_vld;
reg accum_in_ce0;

reg    ap_done_reg;
  reg   [6:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
wire   [3:0] add_ln81_fu_74_p2;
reg   [3:0] add_ln81_reg_91;
wire    ap_CS_fsm_state2;
wire   [0:0] icmp_ln81_fu_85_p2;
wire    ap_CS_fsm_state3;
wire   [15:0] grp_fu_68_p2;
wire    ap_CS_fsm_state7;
reg   [3:0] i_1_1_reg_44;
reg    ap_block_state1;
reg   [15:0] sum_01_reg_55;
wire   [63:0] zext_ln81_fu_80_p1;
reg   [15:0] accum_in_16_preg;
reg   [6:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 7'd1;
#0 accum_in_16_preg = 16'd0;
end

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U100(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(sum_01_reg_55),
    .din1(accum_in_q0),
    .dout(grp_fu_68_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        accum_in_16_preg <= 16'd0;
    end else begin
        if (((icmp_ln81_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
            accum_in_16_preg <= sum_01_reg_55;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if (((icmp_ln81_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        i_1_1_reg_44 <= 4'd0;
    end else if ((1'b1 == ap_CS_fsm_state7)) begin
        i_1_1_reg_44 <= add_ln81_reg_91;
    end
end

always @ (posedge ap_clk) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        sum_01_reg_55 <= 16'd0;
    end else if ((1'b1 == ap_CS_fsm_state7)) begin
        sum_01_reg_55 <= grp_fu_68_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        add_ln81_reg_91 <= add_ln81_fu_74_p2;
    end
end

always @ (*) begin
    if (((icmp_ln81_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        accum_in_16 = sum_01_reg_55;
    end else begin
        accum_in_16 = accum_in_16_preg;
    end
end

always @ (*) begin
    if (((icmp_ln81_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        accum_in_16_ap_vld = 1'b1;
    end else begin
        accum_in_16_ap_vld = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        accum_in_ce0 = 1'b1;
    end else begin
        accum_in_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln81_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln81_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_state2 : begin
            if (((icmp_ln81_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end
        end
        ap_ST_fsm_state3 : begin
            ap_NS_fsm = ap_ST_fsm_state4;
        end
        ap_ST_fsm_state4 : begin
            ap_NS_fsm = ap_ST_fsm_state5;
        end
        ap_ST_fsm_state5 : begin
            ap_NS_fsm = ap_ST_fsm_state6;
        end
        ap_ST_fsm_state6 : begin
            ap_NS_fsm = ap_ST_fsm_state7;
        end
        ap_ST_fsm_state7 : begin
            ap_NS_fsm = ap_ST_fsm_state2;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign accum_in_address0 = zext_ln81_fu_80_p1;

assign add_ln81_fu_74_p2 = (i_1_1_reg_44 + 4'd1);

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state7 = ap_CS_fsm[32'd6];

always @ (*) begin
    ap_block_state1 = ((ap_done_reg == 1'b1) | (ap_start == 1'b0));
end

assign icmp_ln81_fu_85_p2 = ((i_1_1_reg_44 == 4'd8) ? 1'b1 : 1'b0);

assign zext_ln81_fu_80_p1 = i_1_1_reg_44;

endmodule //td_fused_top_tdf2_accum_2
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_tdf2_adjustments_ram (addr0, ce0, q0, addr1, ce1, d1, we1,  clk);

parameter DWIDTH = 48;
parameter AWIDTH = 5;
parameter MEM_SIZE = 32;

input[AWIDTH-1:0] addr0;
input ce0;
output wire[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
input clk;

 reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];
wire [AWIDTH-1:0] addr0_t0; 
reg [AWIDTH-1:0] addr0_t1; 
reg [DWIDTH-1:0] q0_t0;
reg [DWIDTH-1:0] q0_t1;
wire [AWIDTH-1:0] addr1_t0; 
reg [AWIDTH-1:0] addr1_t1; 
wire [DWIDTH-1:0] d1_t0; 
wire we1_t0; 
reg [DWIDTH-1:0] d1_t1; 
reg we1_t1; 


assign addr0_t0 = addr0;
assign q0 = q0_t1;
assign addr1_t0 = addr1;
assign d1_t0 = d1;
assign we1_t0 = we1;

always @(posedge clk)  
begin
    if (ce0) 
    begin
        addr0_t1 <= addr0_t0; 
        q0_t1 <= q0_t0;
    end
    if (ce1) 
    begin
        addr1_t1 <= addr1_t0; 
        d1_t1 <= d1_t0;
        we1_t1 <= we1_t0;
    end
end


always @(posedge clk)  
begin 
    if (ce0) begin
        q0_t0 <= ram[addr0_t1];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1_t1) 
            ram[addr1_t1] <= d1_t1; 
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_tdf2_adjustments(
    reset,
    clk,
    address0,
    ce0,
    q0,
    address1,
    ce1,
    we1,
    d1);

parameter DataWidth = 32'd48;
parameter AddressRange = 32'd32;
parameter AddressWidth = 32'd5;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;



td_fused_top_tdf2_adjustments_ram td_fused_top_tdf2_adjustments_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 )
);

endmodule

// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf2_adjust (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        sums_read,
        adjustments_address0,
        adjustments_ce0,
        adjustments_q0,
        input_indices_23_dout,
        input_indices_23_empty_n,
        input_indices_23_read,
        ap_return
);

parameter    ap_ST_fsm_state1 = 17'd1;
parameter    ap_ST_fsm_state2 = 17'd2;
parameter    ap_ST_fsm_state3 = 17'd4;
parameter    ap_ST_fsm_state4 = 17'd8;
parameter    ap_ST_fsm_state5 = 17'd16;
parameter    ap_ST_fsm_state6 = 17'd32;
parameter    ap_ST_fsm_state7 = 17'd64;
parameter    ap_ST_fsm_state8 = 17'd128;
parameter    ap_ST_fsm_state9 = 17'd256;
parameter    ap_ST_fsm_state10 = 17'd512;
parameter    ap_ST_fsm_state11 = 17'd1024;
parameter    ap_ST_fsm_state12 = 17'd2048;
parameter    ap_ST_fsm_state13 = 17'd4096;
parameter    ap_ST_fsm_state14 = 17'd8192;
parameter    ap_ST_fsm_state15 = 17'd16384;
parameter    ap_ST_fsm_state16 = 17'd32768;
parameter    ap_ST_fsm_state17 = 17'd65536;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
input  [15:0] sums_read;
output  [4:0] adjustments_address0;
output   adjustments_ce0;
input  [47:0] adjustments_q0;
input  [4:0] input_indices_23_dout;
input   input_indices_23_empty_n;
output   input_indices_23_read;
output  [15:0] ap_return;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg adjustments_ce0;
reg input_indices_23_read;

reg    ap_done_reg;
  reg   [16:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    input_indices_23_blk_n;
wire    ap_CS_fsm_state4;
reg   [15:0] tmp_69_i_i_reg_167;
reg   [15:0] tmp_70_i_i_reg_172;
wire   [15:0] grp_fu_81_p2;
reg   [15:0] sub_i_i_i_reg_177;
wire    ap_CS_fsm_state8;
wire    ap_CS_fsm_state9;
wire   [15:0] grp_fu_86_p2;
reg   [15:0] mul_i_i_i_reg_187;
wire    ap_CS_fsm_state12;
wire    ap_CS_fsm_state13;
wire   [63:0] zext_ln220_fu_90_p1;
reg    ap_block_state1;
wire    ap_CS_fsm_state2;
wire    ap_CS_fsm_state3;
wire   [15:0] grp_fu_77_p1;
wire   [15:0] grp_fu_81_p1;
wire   [15:0] grp_fu_86_p1;
wire   [15:0] trunc_ln220_fu_95_p1;
wire   [15:0] grp_fu_77_p2;
wire    ap_CS_fsm_state17;
wire   [15:0] bitcast_ln648_fu_132_p1;
wire   [0:0] tmp_fu_136_p3;
reg   [16:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 17'd1;
end

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U104(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(mul_i_i_i_reg_187),
    .din1(grp_fu_77_p1),
    .dout(grp_fu_77_p2)
);

td_fused_top_hsub_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hsub_16ns_16ns_16_5_full_dsp_1_U105(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(sums_read),
    .din1(grp_fu_81_p1),
    .dout(grp_fu_81_p2)
);

td_fused_top_hmul_16ns_16ns_16_4_max_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hmul_16ns_16ns_16_4_max_dsp_1_U106(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(sub_i_i_i_reg_177),
    .din1(grp_fu_86_p1),
    .dout(grp_fu_86_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state17)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state12)) begin
        mul_i_i_i_reg_187 <= grp_fu_86_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state8)) begin
        sub_i_i_i_reg_177 <= grp_fu_81_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        tmp_69_i_i_reg_167 <= {{adjustments_q0[31:16]}};
        tmp_70_i_i_reg_172 <= {{adjustments_q0[47:32]}};
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state2) | (~((input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1)))) begin
        adjustments_ce0 = 1'b1;
    end else begin
        adjustments_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state17)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state17)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        input_indices_23_blk_n = input_indices_23_empty_n;
    end else begin
        input_indices_23_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        input_indices_23_read = 1'b1;
    end else begin
        input_indices_23_read = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_state2 : begin
            ap_NS_fsm = ap_ST_fsm_state3;
        end
        ap_ST_fsm_state3 : begin
            ap_NS_fsm = ap_ST_fsm_state4;
        end
        ap_ST_fsm_state4 : begin
            ap_NS_fsm = ap_ST_fsm_state5;
        end
        ap_ST_fsm_state5 : begin
            ap_NS_fsm = ap_ST_fsm_state6;
        end
        ap_ST_fsm_state6 : begin
            ap_NS_fsm = ap_ST_fsm_state7;
        end
        ap_ST_fsm_state7 : begin
            ap_NS_fsm = ap_ST_fsm_state8;
        end
        ap_ST_fsm_state8 : begin
            ap_NS_fsm = ap_ST_fsm_state9;
        end
        ap_ST_fsm_state9 : begin
            ap_NS_fsm = ap_ST_fsm_state10;
        end
        ap_ST_fsm_state10 : begin
            ap_NS_fsm = ap_ST_fsm_state11;
        end
        ap_ST_fsm_state11 : begin
            ap_NS_fsm = ap_ST_fsm_state12;
        end
        ap_ST_fsm_state12 : begin
            ap_NS_fsm = ap_ST_fsm_state13;
        end
        ap_ST_fsm_state13 : begin
            ap_NS_fsm = ap_ST_fsm_state14;
        end
        ap_ST_fsm_state14 : begin
            ap_NS_fsm = ap_ST_fsm_state15;
        end
        ap_ST_fsm_state15 : begin
            ap_NS_fsm = ap_ST_fsm_state16;
        end
        ap_ST_fsm_state16 : begin
            ap_NS_fsm = ap_ST_fsm_state17;
        end
        ap_ST_fsm_state17 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign adjustments_address0 = zext_ln220_fu_90_p1;

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state12 = ap_CS_fsm[32'd11];

assign ap_CS_fsm_state13 = ap_CS_fsm[32'd12];

assign ap_CS_fsm_state17 = ap_CS_fsm[32'd16];

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

assign ap_CS_fsm_state8 = ap_CS_fsm[32'd7];

assign ap_CS_fsm_state9 = ap_CS_fsm[32'd8];

always @ (*) begin
    ap_block_state1 = ((input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0));
end

assign ap_return = ((tmp_fu_136_p3[0:0] == 1'b1) ? 16'd0 : grp_fu_77_p2);

assign bitcast_ln648_fu_132_p1 = grp_fu_77_p2;

assign grp_fu_77_p1 = tmp_70_i_i_reg_172;

assign grp_fu_81_p1 = trunc_ln220_fu_95_p1;

assign grp_fu_86_p1 = tmp_69_i_i_reg_167;

assign tmp_fu_136_p3 = bitcast_ln648_fu_132_p1[32'd15];

assign trunc_ln220_fu_95_p1 = adjustments_q0[15:0];

assign zext_ln220_fu_90_p1 = input_indices_23_dout;

endmodule //td_fused_top_tdf2_adjust
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf2_dot_product (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        ifmap_vec_address0,
        ifmap_vec_ce0,
        ifmap_vec_q0,
        weight_vecs_0_address0,
        weight_vecs_0_ce0,
        weight_vecs_0_q0,
        products_0_address0,
        products_0_ce0,
        products_0_we0,
        products_0_d0
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state10 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [7:0] ifmap_vec_address0;
output   ifmap_vec_ce0;
input  [15:0] ifmap_vec_q0;
output  [7:0] weight_vecs_0_address0;
output   weight_vecs_0_ce0;
input  [15:0] weight_vecs_0_q0;
output  [7:0] products_0_address0;
output   products_0_ce0;
output   products_0_we0;
output  [15:0] products_0_d0;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg ifmap_vec_ce0;
reg weight_vecs_0_ce0;
reg products_0_ce0;
reg products_0_we0;

reg    ap_done_reg;
  reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg   [7:0] indvar_flatten17_reg_97;
reg   [6:0] indvar_flatten_reg_108;
reg   [1:0] jj_reg_119;
reg   [4:0] ic_reg_131;
reg   [1:0] ii_reg_142;
wire   [7:0] add_ln147_5_fu_157_p2;
wire    ap_CS_fsm_pp0_stage0;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
wire    ap_block_state4_pp0_stage0_iter2;
wire    ap_block_state5_pp0_stage0_iter3;
wire    ap_block_state6_pp0_stage0_iter4;
wire    ap_block_state7_pp0_stage0_iter5;
wire    ap_block_state8_pp0_stage0_iter6;
wire    ap_block_state9_pp0_stage0_iter7;
wire    ap_block_pp0_stage0_11001;
wire   [0:0] icmp_ln147_fu_163_p2;
reg   [0:0] icmp_ln147_reg_408;
reg   [0:0] icmp_ln147_reg_408_pp0_iter1_reg;
reg   [0:0] icmp_ln147_reg_408_pp0_iter2_reg;
reg   [0:0] icmp_ln147_reg_408_pp0_iter3_reg;
reg   [0:0] icmp_ln147_reg_408_pp0_iter4_reg;
reg   [0:0] icmp_ln147_reg_408_pp0_iter5_reg;
reg   [0:0] icmp_ln147_reg_408_pp0_iter6_reg;
wire   [0:0] icmp_ln148_fu_169_p2;
reg   [0:0] icmp_ln148_reg_412;
wire   [0:0] and_ln147_fu_195_p2;
reg   [0:0] and_ln147_reg_419;
wire   [1:0] add_ln148_fu_201_p2;
reg   [1:0] add_ln148_reg_424;
wire   [4:0] select_ln148_fu_213_p3;
reg   [4:0] select_ln148_reg_429;
wire   [1:0] select_ln148_13_fu_221_p3;
reg   [1:0] select_ln148_13_reg_434;
wire   [3:0] trunc_ln150_fu_229_p1;
reg   [3:0] trunc_ln150_reg_440;
reg   [3:0] trunc_ln150_reg_440_pp0_iter1_reg;
reg   [3:0] trunc_ln150_reg_440_pp0_iter2_reg;
reg   [3:0] trunc_ln150_reg_440_pp0_iter3_reg;
reg   [3:0] trunc_ln150_reg_440_pp0_iter4_reg;
reg   [3:0] trunc_ln150_reg_440_pp0_iter5_reg;
reg   [3:0] trunc_ln150_reg_440_pp0_iter6_reg;
wire   [4:0] add_ln149_fu_233_p2;
wire   [6:0] select_ln148_15_fu_245_p3;
wire   [1:0] select_ln147_14_fu_287_p3;
reg   [1:0] select_ln147_14_reg_455;
reg    ap_enable_reg_pp0_iter1;
wire   [3:0] select_ln148_14_fu_370_p3;
reg   [3:0] select_ln148_14_reg_460;
reg   [3:0] select_ln148_14_reg_460_pp0_iter2_reg;
reg   [3:0] select_ln148_14_reg_460_pp0_iter3_reg;
reg   [3:0] select_ln148_14_reg_460_pp0_iter4_reg;
reg   [3:0] select_ln148_14_reg_460_pp0_iter5_reg;
reg   [3:0] select_ln148_14_reg_460_pp0_iter6_reg;
reg   [15:0] ifmap_vec_load_reg_475;
reg   [15:0] weight_vecs_0_load_reg_480;
wire   [15:0] grp_fu_153_p2;
reg   [15:0] mul_reg_485;
reg    ap_block_state1;
wire    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_flush_enable;
reg    ap_enable_reg_pp0_iter2;
reg    ap_condition_pp0_exit_iter1_state3;
reg    ap_enable_reg_pp0_iter3;
reg    ap_enable_reg_pp0_iter4;
reg    ap_enable_reg_pp0_iter5;
reg    ap_enable_reg_pp0_iter6;
reg    ap_enable_reg_pp0_iter7;
reg   [1:0] ap_phi_mux_jj_phi_fu_123_p4;
wire    ap_block_pp0_stage0;
reg   [1:0] ap_phi_mux_ii_phi_fu_146_p4;
wire   [63:0] p_cast25_fu_386_p1;
wire   [63:0] idxprom30_fu_398_p1;
wire   [0:0] icmp_ln149_fu_189_p2;
wire   [0:0] xor_ln147_fu_183_p2;
wire   [1:0] select_ln147_fu_175_p3;
wire   [0:0] or_ln148_fu_207_p2;
wire   [6:0] add_ln148_5_fu_239_p2;
wire   [3:0] shl_ln_fu_257_p3;
wire   [3:0] zext_ln150_fu_253_p1;
wire   [3:0] sub_ln150_fu_265_p2;
wire   [3:0] zext_ln150_5_fu_271_p1;
wire   [1:0] add_ln147_fu_281_p2;
wire   [3:0] tmp_fu_298_p3;
wire   [3:0] select_ln147_18_cast_fu_294_p1;
wire   [3:0] shl_ln150_mid1_fu_316_p3;
wire   [3:0] zext_ln150_10_fu_312_p1;
wire   [3:0] sub_ln150_5_fu_324_p2;
wire   [3:0] add_ln150_fu_275_p2;
wire   [3:0] empty_112_fu_306_p2;
wire   [3:0] select_ln148_17_cast_fu_344_p1;
wire   [3:0] empty_113_fu_347_p2;
wire   [3:0] select_ln147_15_fu_330_p3;
wire   [3:0] zext_ln150_11_fu_361_p1;
wire   [3:0] add_ln150_5_fu_364_p2;
wire   [3:0] select_ln147_16_fu_337_p3;
wire   [7:0] tmp_128_cast_fu_353_p3;
wire   [7:0] select_ln148_cast_fu_377_p1;
wire   [7:0] empty_114_fu_380_p2;
wire   [7:0] p_fu_392_p3;
wire    ap_CS_fsm_state10;
reg   [2:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
#0 ap_enable_reg_pp0_iter4 = 1'b0;
#0 ap_enable_reg_pp0_iter5 = 1'b0;
#0 ap_enable_reg_pp0_iter6 = 1'b0;
#0 ap_enable_reg_pp0_iter7 = 1'b0;
end

td_fused_top_hmul_16ns_16ns_16_4_max_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hmul_16ns_16ns_16_4_max_dsp_1_U92(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(ifmap_vec_load_reg_475),
    .din1(weight_vecs_0_load_reg_480),
    .dout(grp_fu_153_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state10)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if ((1'b1 == ap_condition_pp0_flush_enable)) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            if ((1'b1 == ap_condition_pp0_exit_iter1_state3)) begin
                ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter0;
            end else if ((1'b1 == 1'b1)) begin
                ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
            end
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter4 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter5 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter5 <= ap_enable_reg_pp0_iter4;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter6 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter6 <= ap_enable_reg_pp0_iter5;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter7 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter7 <= ap_enable_reg_pp0_iter6;
        end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter7 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_fu_163_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ic_reg_131 <= add_ln149_fu_233_p2;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ic_reg_131 <= 5'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_reg_408_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        ii_reg_142 <= select_ln147_14_reg_455;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ii_reg_142 <= 2'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_fu_163_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        indvar_flatten17_reg_97 <= add_ln147_5_fu_157_p2;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indvar_flatten17_reg_97 <= 8'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_fu_163_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        indvar_flatten_reg_108 <= select_ln148_15_fu_245_p3;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indvar_flatten_reg_108 <= 7'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_reg_408 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        jj_reg_119 <= select_ln148_13_reg_434;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        jj_reg_119 <= 2'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_fu_163_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        add_ln148_reg_424 <= add_ln148_fu_201_p2;
        and_ln147_reg_419 <= and_ln147_fu_195_p2;
        icmp_ln148_reg_412 <= icmp_ln148_fu_169_p2;
        select_ln148_reg_429 <= select_ln148_fu_213_p3;
        trunc_ln150_reg_440 <= trunc_ln150_fu_229_p1;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln147_reg_408 <= icmp_ln147_fu_163_p2;
        icmp_ln147_reg_408_pp0_iter1_reg <= icmp_ln147_reg_408;
        trunc_ln150_reg_440_pp0_iter1_reg <= trunc_ln150_reg_440;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        icmp_ln147_reg_408_pp0_iter2_reg <= icmp_ln147_reg_408_pp0_iter1_reg;
        icmp_ln147_reg_408_pp0_iter3_reg <= icmp_ln147_reg_408_pp0_iter2_reg;
        icmp_ln147_reg_408_pp0_iter4_reg <= icmp_ln147_reg_408_pp0_iter3_reg;
        icmp_ln147_reg_408_pp0_iter5_reg <= icmp_ln147_reg_408_pp0_iter4_reg;
        icmp_ln147_reg_408_pp0_iter6_reg <= icmp_ln147_reg_408_pp0_iter5_reg;
        select_ln148_14_reg_460_pp0_iter2_reg <= select_ln148_14_reg_460;
        select_ln148_14_reg_460_pp0_iter3_reg <= select_ln148_14_reg_460_pp0_iter2_reg;
        select_ln148_14_reg_460_pp0_iter4_reg <= select_ln148_14_reg_460_pp0_iter3_reg;
        select_ln148_14_reg_460_pp0_iter5_reg <= select_ln148_14_reg_460_pp0_iter4_reg;
        select_ln148_14_reg_460_pp0_iter6_reg <= select_ln148_14_reg_460_pp0_iter5_reg;
        trunc_ln150_reg_440_pp0_iter2_reg <= trunc_ln150_reg_440_pp0_iter1_reg;
        trunc_ln150_reg_440_pp0_iter3_reg <= trunc_ln150_reg_440_pp0_iter2_reg;
        trunc_ln150_reg_440_pp0_iter4_reg <= trunc_ln150_reg_440_pp0_iter3_reg;
        trunc_ln150_reg_440_pp0_iter5_reg <= trunc_ln150_reg_440_pp0_iter4_reg;
        trunc_ln150_reg_440_pp0_iter6_reg <= trunc_ln150_reg_440_pp0_iter5_reg;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_reg_408_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        ifmap_vec_load_reg_475 <= ifmap_vec_q0;
        weight_vecs_0_load_reg_480 <= weight_vecs_0_q0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_reg_408_pp0_iter5_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        mul_reg_485 <= grp_fu_153_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_reg_408 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        select_ln147_14_reg_455 <= select_ln147_14_fu_287_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_fu_163_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        select_ln148_13_reg_434 <= select_ln148_13_fu_221_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_reg_408 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        select_ln148_14_reg_460 <= select_ln148_14_fu_370_p3;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_condition_pp0_exit_iter1_state3 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter1_state3 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln147_fu_163_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_condition_pp0_flush_enable = 1'b1;
    end else begin
        ap_condition_pp0_flush_enable = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state10)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter7 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln147_reg_408_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        ap_phi_mux_ii_phi_fu_146_p4 = select_ln147_14_reg_455;
    end else begin
        ap_phi_mux_ii_phi_fu_146_p4 = ii_reg_142;
    end
end

always @ (*) begin
    if (((icmp_ln147_reg_408 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_jj_phi_fu_123_p4 = select_ln148_13_reg_434;
    end else begin
        ap_phi_mux_jj_phi_fu_123_p4 = jj_reg_119;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state10)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ifmap_vec_ce0 = 1'b1;
    end else begin
        ifmap_vec_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter7 == 1'b1))) begin
        products_0_ce0 = 1'b1;
    end else begin
        products_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln147_reg_408_pp0_iter6_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter7 == 1'b1))) begin
        products_0_we0 = 1'b1;
    end else begin
        products_0_we0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        weight_vecs_0_ce0 = 1'b1;
    end else begin
        weight_vecs_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((~((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b1)) & ~((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter7 == 1'b1) & (ap_enable_reg_pp0_iter6 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if ((((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter7 == 1'b1) & (ap_enable_reg_pp0_iter6 == 1'b0)) | ((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b1)))) begin
                ap_NS_fsm = ap_ST_fsm_state10;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state10 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln147_5_fu_157_p2 = (indvar_flatten17_reg_97 + 8'd1);

assign add_ln147_fu_281_p2 = (ap_phi_mux_ii_phi_fu_146_p4 + 2'd1);

assign add_ln148_5_fu_239_p2 = (indvar_flatten_reg_108 + 7'd1);

assign add_ln148_fu_201_p2 = (select_ln147_fu_175_p3 + 2'd1);

assign add_ln149_fu_233_p2 = (select_ln148_fu_213_p3 + 5'd1);

assign add_ln150_5_fu_364_p2 = (select_ln147_15_fu_330_p3 + zext_ln150_11_fu_361_p1);

assign add_ln150_fu_275_p2 = (sub_ln150_fu_265_p2 + zext_ln150_5_fu_271_p1);

assign and_ln147_fu_195_p2 = (xor_ln147_fu_183_p2 & icmp_ln149_fu_189_p2);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state10 = ap_CS_fsm[32'd2];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (ap_done_reg == 1'b1));
end

assign ap_block_state2_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter4 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage0_iter5 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage0_iter6 = ~(1'b1 == 1'b1);

assign ap_block_state9_pp0_stage0_iter7 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign empty_112_fu_306_p2 = (tmp_fu_298_p3 - select_ln147_18_cast_fu_294_p1);

assign empty_113_fu_347_p2 = (empty_112_fu_306_p2 + select_ln148_17_cast_fu_344_p1);

assign empty_114_fu_380_p2 = (tmp_128_cast_fu_353_p3 + select_ln148_cast_fu_377_p1);

assign icmp_ln147_fu_163_p2 = ((indvar_flatten17_reg_97 == 8'd144) ? 1'b1 : 1'b0);

assign icmp_ln148_fu_169_p2 = ((indvar_flatten_reg_108 == 7'd48) ? 1'b1 : 1'b0);

assign icmp_ln149_fu_189_p2 = ((ic_reg_131 == 5'd16) ? 1'b1 : 1'b0);

assign idxprom30_fu_398_p1 = p_fu_392_p3;

assign ifmap_vec_address0 = p_cast25_fu_386_p1;

assign or_ln148_fu_207_p2 = (icmp_ln148_fu_169_p2 | and_ln147_fu_195_p2);

assign p_cast25_fu_386_p1 = empty_114_fu_380_p2;

assign p_fu_392_p3 = {{select_ln148_14_reg_460_pp0_iter6_reg}, {trunc_ln150_reg_440_pp0_iter6_reg}};

assign products_0_address0 = idxprom30_fu_398_p1;

assign products_0_d0 = mul_reg_485;

assign select_ln147_14_fu_287_p3 = ((icmp_ln148_reg_412[0:0] == 1'b1) ? add_ln147_fu_281_p2 : ap_phi_mux_ii_phi_fu_146_p4);

assign select_ln147_15_fu_330_p3 = ((icmp_ln148_reg_412[0:0] == 1'b1) ? sub_ln150_5_fu_324_p2 : sub_ln150_fu_265_p2);

assign select_ln147_16_fu_337_p3 = ((icmp_ln148_reg_412[0:0] == 1'b1) ? sub_ln150_5_fu_324_p2 : add_ln150_fu_275_p2);

assign select_ln147_18_cast_fu_294_p1 = select_ln147_14_fu_287_p3;

assign select_ln147_fu_175_p3 = ((icmp_ln148_fu_169_p2[0:0] == 1'b1) ? 2'd0 : ap_phi_mux_jj_phi_fu_123_p4);

assign select_ln148_13_fu_221_p3 = ((and_ln147_fu_195_p2[0:0] == 1'b1) ? add_ln148_fu_201_p2 : select_ln147_fu_175_p3);

assign select_ln148_14_fu_370_p3 = ((and_ln147_reg_419[0:0] == 1'b1) ? add_ln150_5_fu_364_p2 : select_ln147_16_fu_337_p3);

assign select_ln148_15_fu_245_p3 = ((icmp_ln148_fu_169_p2[0:0] == 1'b1) ? 7'd1 : add_ln148_5_fu_239_p2);

assign select_ln148_17_cast_fu_344_p1 = select_ln148_13_reg_434;

assign select_ln148_cast_fu_377_p1 = select_ln148_reg_429;

assign select_ln148_fu_213_p3 = ((or_ln148_fu_207_p2[0:0] == 1'b1) ? 5'd0 : ic_reg_131);

assign shl_ln150_mid1_fu_316_p3 = {{add_ln147_fu_281_p2}, {2'd0}};

assign shl_ln_fu_257_p3 = {{ap_phi_mux_ii_phi_fu_146_p4}, {2'd0}};

assign sub_ln150_5_fu_324_p2 = (shl_ln150_mid1_fu_316_p3 - zext_ln150_10_fu_312_p1);

assign sub_ln150_fu_265_p2 = (shl_ln_fu_257_p3 - zext_ln150_fu_253_p1);

assign tmp_128_cast_fu_353_p3 = {{empty_113_fu_347_p2}, {4'd0}};

assign tmp_fu_298_p3 = {{select_ln147_14_fu_287_p3}, {2'd0}};

assign trunc_ln150_fu_229_p1 = select_ln148_fu_213_p3[3:0];

assign weight_vecs_0_address0 = p_cast25_fu_386_p1;

assign xor_ln147_fu_183_p2 = (icmp_ln148_fu_169_p2 ^ 1'd1);

assign zext_ln150_10_fu_312_p1 = add_ln147_fu_281_p2;

assign zext_ln150_11_fu_361_p1 = add_ln148_reg_424;

assign zext_ln150_5_fu_271_p1 = jj_reg_119;

assign zext_ln150_fu_253_p1 = ap_phi_mux_ii_phi_fu_146_p4;

endmodule //td_fused_top_tdf2_dot_product
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_tdf2_filters_ram (addr0, ce0, q0, addr1, ce1, d1, we1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 13;
parameter MEM_SIZE = 4608;

input[AWIDTH-1:0] addr0;
input ce0;
output wire[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
input clk;

 reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];
wire [AWIDTH-1:0] addr0_t0; 
reg [AWIDTH-1:0] addr0_t1; 
reg [DWIDTH-1:0] q0_t0;
reg [DWIDTH-1:0] q0_t1;
wire [AWIDTH-1:0] addr1_t0; 
reg [AWIDTH-1:0] addr1_t1; 
wire [DWIDTH-1:0] d1_t0; 
wire we1_t0; 
reg [DWIDTH-1:0] d1_t1; 
reg we1_t1; 


assign addr0_t0 = addr0;
assign q0 = q0_t1;
assign addr1_t0 = addr1;
assign d1_t0 = d1;
assign we1_t0 = we1;

always @(posedge clk)  
begin
    if (ce0) 
    begin
        addr0_t1 <= addr0_t0; 
        q0_t1 <= q0_t0;
    end
    if (ce1) 
    begin
        addr1_t1 <= addr1_t0; 
        d1_t1 <= d1_t0;
        we1_t1 <= we1_t0;
    end
end


always @(posedge clk)  
begin 
    if (ce0) begin
        q0_t0 <= ram[addr0_t1];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1_t1) 
            ram[addr1_t1] <= d1_t1; 
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_tdf2_filters(
    reset,
    clk,
    address0,
    ce0,
    q0,
    address1,
    ce1,
    we1,
    d1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd4608;
parameter AddressWidth = 32'd13;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;



td_fused_top_tdf2_filters_ram td_fused_top_tdf2_filters_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 )
);

endmodule

// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf2_get_next_ijk (
        ap_clk,
        ap_rst,
        ap_start,
        start_full_n,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        start_out,
        start_write,
        input_indices_2_out_din,
        input_indices_2_out_full_n,
        input_indices_2_out_write,
        input_indices_2_out1_din,
        input_indices_2_out1_full_n,
        input_indices_2_out1_write,
        output_indices_0_din,
        output_indices_0_full_n,
        output_indices_0_write,
        output_indices_1_din,
        output_indices_1_full_n,
        output_indices_1_write,
        resetMaximum_din,
        resetMaximum_full_n,
        resetMaximum_write,
        storeOutput_din,
        storeOutput_full_n,
        storeOutput_write,
        ap_return_0,
        ap_return_1
);

parameter    ap_ST_fsm_state1 = 1'd1;

input   ap_clk;
input   ap_rst;
input   ap_start;
input   start_full_n;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output   start_out;
output   start_write;
output  [4:0] input_indices_2_out_din;
input   input_indices_2_out_full_n;
output   input_indices_2_out_write;
output  [4:0] input_indices_2_out1_din;
input   input_indices_2_out1_full_n;
output   input_indices_2_out1_write;
output  [5:0] output_indices_0_din;
input   output_indices_0_full_n;
output   output_indices_0_write;
output  [11:0] output_indices_1_din;
input   output_indices_1_full_n;
output   output_indices_1_write;
output   resetMaximum_din;
input   resetMaximum_full_n;
output   resetMaximum_write;
output   storeOutput_din;
input   storeOutput_full_n;
output   storeOutput_write;
output  [15:0] ap_return_0;
output  [15:0] ap_return_1;

reg ap_done;
reg ap_idle;
reg start_write;
reg input_indices_2_out_write;
reg input_indices_2_out1_write;
reg output_indices_0_write;
reg output_indices_1_write;
reg resetMaximum_write;
reg storeOutput_write;

reg    real_start;
reg    start_once_reg;
reg    ap_done_reg;
  reg   [0:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    internal_ap_ready;
reg   [1:0] i_p_2;
reg   [1:0] j_p_2;
reg   [15:0] i_6;
reg   [15:0] j_6;
reg   [15:0] k_6;
reg   [15:0] i_out_2;
reg   [15:0] j_out_2;
reg    input_indices_2_out_blk_n;
reg    input_indices_2_out1_blk_n;
reg    output_indices_0_blk_n;
reg    output_indices_1_blk_n;
reg    resetMaximum_blk_n;
reg    storeOutput_blk_n;
wire   [1:0] select_ln142_fu_338_p3;
reg    ap_block_state1;
wire   [0:0] or_ln142_fu_312_p2;
wire   [1:0] select_ln142_9_fu_346_p3;
wire   [15:0] select_ln147_fu_278_p3;
wire   [0:0] and_ln142_3_fu_306_p2;
wire   [15:0] select_ln142_10_fu_360_p3;
wire   [0:0] and_ln132_fu_354_p2;
wire   [15:0] select_ln142_11_fu_388_p3;
wire   [0:0] and_ln135_fu_294_p2;
wire   [15:0] select_ln147_3_fu_286_p3;
wire   [15:0] select_ln142_12_fu_396_p3;
wire   [4:0] trunc_ln128_fu_182_p1;
wire   [1:0] or_ln124_fu_126_p2;
wire   [0:0] icmp_ln125_fu_139_p2;
wire   [0:0] icmp_ln125_3_fu_145_p2;
wire   [15:0] zext_ln126_fu_114_p1;
wire   [15:0] zext_ln127_fu_122_p1;
wire   [1:0] add_ln131_fu_206_p2;
wire   [1:0] add_ln134_fu_218_p2;
wire   [15:0] add_ln137_fu_230_p2;
wire   [15:0] add_ln141_fu_248_p2;
wire   [15:0] add_ln146_fu_266_p2;
wire   [0:0] icmp_ln147_fu_272_p2;
wire   [15:0] add_ln145_fu_260_p2;
wire   [0:0] icmp_ln132_fu_212_p2;
wire   [0:0] icmp_ln135_fu_224_p2;
wire   [0:0] icmp_ln138_fu_236_p2;
wire   [0:0] icmp_ln142_fu_254_p2;
wire   [0:0] and_ln142_fu_300_p2;
wire   [0:0] xor_ln135_fu_318_p2;
wire   [0:0] and_ln135_3_fu_324_p2;
wire   [1:0] select_ln135_fu_330_p3;
wire   [15:0] add_ln140_fu_242_p2;
wire   [0:0] xor_ln138_fu_368_p2;
wire   [0:0] and_ln138_fu_374_p2;
wire   [15:0] select_ln138_fu_380_p3;
wire   [15:0] add_ln126_fu_162_p2;
wire   [15:0] add_ln127_fu_172_p2;
reg   [0:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 start_once_reg = 1'b0;
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 1'd1;
#0 i_p_2 = 2'd0;
#0 j_p_2 = 2'd0;
#0 i_6 = 16'd0;
#0 j_6 = 16'd0;
#0 k_6 = 16'd0;
#0 i_out_2 = 16'd0;
#0 j_out_2 = 16'd0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        start_once_reg <= 1'b0;
    end else begin
        if (((real_start == 1'b1) & (internal_ap_ready == 1'b0))) begin
            start_once_reg <= 1'b1;
        end else if ((internal_ap_ready == 1'b1)) begin
            start_once_reg <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1) & (1'd1 == and_ln142_3_fu_306_p2))) begin
        i_6 <= select_ln147_fu_278_p3;
        i_out_2 <= select_ln147_3_fu_286_p3;
    end
end

always @ (posedge ap_clk) begin
    if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (or_ln142_fu_312_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1))) begin
        i_p_2 <= select_ln142_fu_338_p3;
    end
end

always @ (posedge ap_clk) begin
    if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1) & (1'd1 == and_ln132_fu_354_p2))) begin
        j_6 <= select_ln142_10_fu_360_p3;
        j_out_2 <= select_ln142_12_fu_396_p3;
    end
end

always @ (posedge ap_clk) begin
    if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        j_p_2 <= select_ln142_9_fu_346_p3;
    end
end

always @ (posedge ap_clk) begin
    if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1) & (1'd1 == and_ln135_fu_294_p2))) begin
        k_6 <= select_ln142_11_fu_388_p3;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((real_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        input_indices_2_out1_blk_n = input_indices_2_out1_full_n;
    end else begin
        input_indices_2_out1_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        input_indices_2_out1_write = 1'b1;
    end else begin
        input_indices_2_out1_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        input_indices_2_out_blk_n = input_indices_2_out_full_n;
    end else begin
        input_indices_2_out_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        input_indices_2_out_write = 1'b1;
    end else begin
        input_indices_2_out_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        internal_ap_ready = 1'b1;
    end else begin
        internal_ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        output_indices_0_blk_n = output_indices_0_full_n;
    end else begin
        output_indices_0_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        output_indices_0_write = 1'b1;
    end else begin
        output_indices_0_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        output_indices_1_blk_n = output_indices_1_full_n;
    end else begin
        output_indices_1_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        output_indices_1_write = 1'b1;
    end else begin
        output_indices_1_write = 1'b0;
    end
end

always @ (*) begin
    if (((start_full_n == 1'b0) & (start_once_reg == 1'b0))) begin
        real_start = 1'b0;
    end else begin
        real_start = ap_start;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        resetMaximum_blk_n = resetMaximum_full_n;
    end else begin
        resetMaximum_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        resetMaximum_write = 1'b1;
    end else begin
        resetMaximum_write = 1'b0;
    end
end

always @ (*) begin
    if (((real_start == 1'b1) & (start_once_reg == 1'b0))) begin
        start_write = 1'b1;
    end else begin
        start_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        storeOutput_blk_n = storeOutput_full_n;
    end else begin
        storeOutput_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        storeOutput_write = 1'b1;
    end else begin
        storeOutput_write = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln126_fu_162_p2 = (i_6 + zext_ln126_fu_114_p1);

assign add_ln127_fu_172_p2 = (j_6 + zext_ln127_fu_122_p1);

assign add_ln131_fu_206_p2 = (j_p_2 + 2'd1);

assign add_ln134_fu_218_p2 = (i_p_2 + 2'd1);

assign add_ln137_fu_230_p2 = (k_6 + 16'd1);

assign add_ln140_fu_242_p2 = (j_6 + 16'd2);

assign add_ln141_fu_248_p2 = (j_out_2 + 16'd1);

assign add_ln145_fu_260_p2 = (i_6 + 16'd2);

assign add_ln146_fu_266_p2 = (i_out_2 + 16'd1);

assign and_ln132_fu_354_p2 = (icmp_ln138_fu_236_p2 & and_ln135_fu_294_p2);

assign and_ln135_3_fu_324_p2 = (xor_ln135_fu_318_p2 & icmp_ln132_fu_212_p2);

assign and_ln135_fu_294_p2 = (icmp_ln135_fu_224_p2 & icmp_ln132_fu_212_p2);

assign and_ln138_fu_374_p2 = (xor_ln138_fu_368_p2 & and_ln135_fu_294_p2);

assign and_ln142_3_fu_306_p2 = (and_ln142_fu_300_p2 & and_ln135_fu_294_p2);

assign and_ln142_fu_300_p2 = (icmp_ln142_fu_254_p2 & icmp_ln138_fu_236_p2);

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

always @ (*) begin
    ap_block_state1 = ((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1));
end

assign ap_ready = internal_ap_ready;

assign ap_return_0 = add_ln126_fu_162_p2;

assign ap_return_1 = add_ln127_fu_172_p2;

assign icmp_ln125_3_fu_145_p2 = ((j_p_2 == 2'd1) ? 1'b1 : 1'b0);

assign icmp_ln125_fu_139_p2 = ((i_p_2 == 2'd1) ? 1'b1 : 1'b0);

assign icmp_ln132_fu_212_p2 = ((add_ln131_fu_206_p2 == 2'd2) ? 1'b1 : 1'b0);

assign icmp_ln135_fu_224_p2 = ((add_ln134_fu_218_p2 == 2'd2) ? 1'b1 : 1'b0);

assign icmp_ln138_fu_236_p2 = ((add_ln137_fu_230_p2 == 16'd32) ? 1'b1 : 1'b0);

assign icmp_ln142_fu_254_p2 = ((add_ln141_fu_248_p2 == 16'd56) ? 1'b1 : 1'b0);

assign icmp_ln147_fu_272_p2 = ((add_ln146_fu_266_p2 == 16'd56) ? 1'b1 : 1'b0);

assign input_indices_2_out1_din = trunc_ln128_fu_182_p1;

assign input_indices_2_out_din = trunc_ln128_fu_182_p1;

assign or_ln124_fu_126_p2 = (j_p_2 | i_p_2);

assign or_ln142_fu_312_p2 = (icmp_ln132_fu_212_p2 | and_ln142_3_fu_306_p2);

assign output_indices_0_din = i_out_2[5:0];

assign output_indices_1_din = j_out_2[11:0];

assign resetMaximum_din = ((or_ln124_fu_126_p2 == 2'd0) ? 1'b1 : 1'b0);

assign select_ln135_fu_330_p3 = ((and_ln135_3_fu_324_p2[0:0] == 1'b1) ? add_ln134_fu_218_p2 : 2'd0);

assign select_ln138_fu_380_p3 = ((and_ln138_fu_374_p2[0:0] == 1'b1) ? add_ln137_fu_230_p2 : 16'd0);

assign select_ln142_10_fu_360_p3 = ((and_ln142_3_fu_306_p2[0:0] == 1'b1) ? 16'd0 : add_ln140_fu_242_p2);

assign select_ln142_11_fu_388_p3 = ((and_ln142_3_fu_306_p2[0:0] == 1'b1) ? 16'd0 : select_ln138_fu_380_p3);

assign select_ln142_12_fu_396_p3 = ((and_ln142_3_fu_306_p2[0:0] == 1'b1) ? 16'd0 : add_ln141_fu_248_p2);

assign select_ln142_9_fu_346_p3 = ((or_ln142_fu_312_p2[0:0] == 1'b1) ? 2'd0 : add_ln131_fu_206_p2);

assign select_ln142_fu_338_p3 = ((and_ln142_3_fu_306_p2[0:0] == 1'b1) ? 2'd0 : select_ln135_fu_330_p3);

assign select_ln147_3_fu_286_p3 = ((icmp_ln147_fu_272_p2[0:0] == 1'b1) ? 16'd0 : add_ln146_fu_266_p2);

assign select_ln147_fu_278_p3 = ((icmp_ln147_fu_272_p2[0:0] == 1'b1) ? 16'd0 : add_ln145_fu_260_p2);

assign start_out = real_start;

assign storeOutput_din = (icmp_ln125_fu_139_p2 & icmp_ln125_3_fu_145_p2);

assign trunc_ln128_fu_182_p1 = k_6[4:0];

assign xor_ln135_fu_318_p2 = (icmp_ln135_fu_224_p2 ^ 1'd1);

assign xor_ln138_fu_368_p2 = (icmp_ln138_fu_236_p2 ^ 1'd1);

assign zext_ln126_fu_114_p1 = i_p_2;

assign zext_ln127_fu_122_p1 = j_p_2;

endmodule //td_fused_top_tdf2_get_next_ijk
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf2_poolOutputs (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        output_indices_04_dout,
        output_indices_04_empty_n,
        output_indices_04_read,
        output_indices_15_dout,
        output_indices_15_empty_n,
        output_indices_15_read,
        resetMaximum6_dout,
        resetMaximum6_empty_n,
        resetMaximum6_read,
        storeOutput7_dout,
        storeOutput7_empty_n,
        storeOutput7_read,
        p_read,
        out_data_address1,
        out_data_ce1,
        out_data_we1,
        out_data_d1
);

parameter    ap_ST_fsm_state1 = 4'd1;
parameter    ap_ST_fsm_state2 = 4'd2;
parameter    ap_ST_fsm_state3 = 4'd4;
parameter    ap_ST_fsm_state4 = 4'd8;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
input  [5:0] output_indices_04_dout;
input   output_indices_04_empty_n;
output   output_indices_04_read;
input  [11:0] output_indices_15_dout;
input   output_indices_15_empty_n;
output   output_indices_15_read;
input  [0:0] resetMaximum6_dout;
input   resetMaximum6_empty_n;
output   resetMaximum6_read;
input  [0:0] storeOutput7_dout;
input   storeOutput7_empty_n;
output   storeOutput7_read;
input  [15:0] p_read;
output  [14:0] out_data_address1;
output   out_data_ce1;
output   out_data_we1;
output  [63:0] out_data_d1;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg output_indices_04_read;
reg output_indices_15_read;
reg resetMaximum6_read;
reg storeOutput7_read;

reg    ap_done_reg;
  reg   [3:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg   [15:0] max_vals_4_0;
reg    output_indices_04_blk_n;
wire    ap_CS_fsm_state2;
reg    output_indices_15_blk_n;
reg    resetMaximum6_blk_n;
reg    storeOutput7_blk_n;
reg   [5:0] output_indices_04_read_reg_147;
reg   [11:0] output_indices_15_read_reg_152;
wire   [0:0] storeOutput7_read_read_fu_82_p2;
reg   [0:0] storeOutput7_read_reg_157;
wire    grp_tdf2_writeOutputs_unaligned_fu_88_ap_start;
wire    grp_tdf2_writeOutputs_unaligned_fu_88_ap_done;
wire    grp_tdf2_writeOutputs_unaligned_fu_88_ap_idle;
wire    grp_tdf2_writeOutputs_unaligned_fu_88_ap_ready;
wire   [14:0] grp_tdf2_writeOutputs_unaligned_fu_88_out_data_address1;
wire    grp_tdf2_writeOutputs_unaligned_fu_88_out_data_ce1;
wire    grp_tdf2_writeOutputs_unaligned_fu_88_out_data_we1;
wire   [63:0] grp_tdf2_writeOutputs_unaligned_fu_88_out_data_d1;
reg    grp_tdf2_writeOutputs_unaligned_fu_88_ap_start_reg;
wire    ap_CS_fsm_state3;
wire    ap_CS_fsm_state4;
reg    ap_block_state4_on_subcall_done;
wire   [15:0] select_ln24_fu_126_p3;
reg    ap_block_state2;
reg    ap_block_state1;
wire   [0:0] grp_fu_110_p2;
wire   [0:0] or_ln24_fu_120_p2;
reg    grp_fu_110_ce;
reg   [3:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 4'd1;
#0 max_vals_4_0 = 16'd0;
#0 grp_tdf2_writeOutputs_unaligned_fu_88_ap_start_reg = 1'b0;
end

td_fused_top_tdf2_writeOutputs_unaligned grp_tdf2_writeOutputs_unaligned_fu_88(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(grp_tdf2_writeOutputs_unaligned_fu_88_ap_start),
    .ap_done(grp_tdf2_writeOutputs_unaligned_fu_88_ap_done),
    .ap_idle(grp_tdf2_writeOutputs_unaligned_fu_88_ap_idle),
    .ap_ready(grp_tdf2_writeOutputs_unaligned_fu_88_ap_ready),
    .i(output_indices_04_read_reg_147),
    .j(output_indices_15_read_reg_152),
    .out_data_address1(grp_tdf2_writeOutputs_unaligned_fu_88_out_data_address1),
    .out_data_ce1(grp_tdf2_writeOutputs_unaligned_fu_88_out_data_ce1),
    .out_data_we1(grp_tdf2_writeOutputs_unaligned_fu_88_out_data_we1),
    .out_data_d1(grp_tdf2_writeOutputs_unaligned_fu_88_out_data_d1),
    .max_vals_4_0(max_vals_4_0)
);

td_fused_top_hcmp_16ns_16ns_1_2_no_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 1 ))
hcmp_16ns_16ns_1_2_no_dsp_1_U114(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(grp_fu_110_ce),
    .din0(max_vals_4_0),
    .din1(p_read),
    .opcode(5'd4),
    .dout(grp_fu_110_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_state4) & (1'b0 == ap_block_state4_on_subcall_done))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        grp_tdf2_writeOutputs_unaligned_fu_88_ap_start_reg <= 1'b0;
    end else begin
        if ((1'b1 == ap_CS_fsm_state3)) begin
            grp_tdf2_writeOutputs_unaligned_fu_88_ap_start_reg <= 1'b1;
        end else if ((grp_tdf2_writeOutputs_unaligned_fu_88_ap_ready == 1'b1)) begin
            grp_tdf2_writeOutputs_unaligned_fu_88_ap_start_reg <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((~((storeOutput7_empty_n == 1'b0) | (resetMaximum6_empty_n == 1'b0) | (output_indices_15_empty_n == 1'b0) | (output_indices_04_empty_n == 1'b0)) & (1'b1 == ap_CS_fsm_state2))) begin
        max_vals_4_0 <= select_ln24_fu_126_p3;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        output_indices_04_read_reg_147 <= output_indices_04_dout;
        output_indices_15_read_reg_152 <= output_indices_15_dout;
        storeOutput7_read_reg_157 <= storeOutput7_dout;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state4) & (1'b0 == ap_block_state4_on_subcall_done))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state4) & (1'b0 == ap_block_state4_on_subcall_done))) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1)) | (~((storeOutput7_empty_n == 1'b0) | (resetMaximum6_empty_n == 1'b0) | (output_indices_15_empty_n == 1'b0) | (output_indices_04_empty_n == 1'b0)) & (1'b1 == ap_CS_fsm_state2)))) begin
        grp_fu_110_ce = 1'b1;
    end else begin
        grp_fu_110_ce = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        output_indices_04_blk_n = output_indices_04_empty_n;
    end else begin
        output_indices_04_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((storeOutput7_empty_n == 1'b0) | (resetMaximum6_empty_n == 1'b0) | (output_indices_15_empty_n == 1'b0) | (output_indices_04_empty_n == 1'b0)) & (1'b1 == ap_CS_fsm_state2))) begin
        output_indices_04_read = 1'b1;
    end else begin
        output_indices_04_read = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        output_indices_15_blk_n = output_indices_15_empty_n;
    end else begin
        output_indices_15_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((storeOutput7_empty_n == 1'b0) | (resetMaximum6_empty_n == 1'b0) | (output_indices_15_empty_n == 1'b0) | (output_indices_04_empty_n == 1'b0)) & (1'b1 == ap_CS_fsm_state2))) begin
        output_indices_15_read = 1'b1;
    end else begin
        output_indices_15_read = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        resetMaximum6_blk_n = resetMaximum6_empty_n;
    end else begin
        resetMaximum6_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((storeOutput7_empty_n == 1'b0) | (resetMaximum6_empty_n == 1'b0) | (output_indices_15_empty_n == 1'b0) | (output_indices_04_empty_n == 1'b0)) & (1'b1 == ap_CS_fsm_state2))) begin
        resetMaximum6_read = 1'b1;
    end else begin
        resetMaximum6_read = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        storeOutput7_blk_n = storeOutput7_empty_n;
    end else begin
        storeOutput7_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((storeOutput7_empty_n == 1'b0) | (resetMaximum6_empty_n == 1'b0) | (output_indices_15_empty_n == 1'b0) | (output_indices_04_empty_n == 1'b0)) & (1'b1 == ap_CS_fsm_state2))) begin
        storeOutput7_read = 1'b1;
    end else begin
        storeOutput7_read = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_state2 : begin
            if ((~((storeOutput7_empty_n == 1'b0) | (resetMaximum6_empty_n == 1'b0) | (output_indices_15_empty_n == 1'b0) | (output_indices_04_empty_n == 1'b0)) & (storeOutput7_read_read_fu_82_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state2))) begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end else if ((~((storeOutput7_empty_n == 1'b0) | (resetMaximum6_empty_n == 1'b0) | (output_indices_15_empty_n == 1'b0) | (output_indices_04_empty_n == 1'b0)) & (storeOutput7_read_read_fu_82_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end
        end
        ap_ST_fsm_state3 : begin
            ap_NS_fsm = ap_ST_fsm_state4;
        end
        ap_ST_fsm_state4 : begin
            if (((1'b1 == ap_CS_fsm_state4) & (1'b0 == ap_block_state4_on_subcall_done))) begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (ap_done_reg == 1'b1));
end

always @ (*) begin
    ap_block_state2 = ((storeOutput7_empty_n == 1'b0) | (resetMaximum6_empty_n == 1'b0) | (output_indices_15_empty_n == 1'b0) | (output_indices_04_empty_n == 1'b0));
end

always @ (*) begin
    ap_block_state4_on_subcall_done = ((grp_tdf2_writeOutputs_unaligned_fu_88_ap_done == 1'b0) & (storeOutput7_read_reg_157 == 1'd1));
end

assign grp_tdf2_writeOutputs_unaligned_fu_88_ap_start = grp_tdf2_writeOutputs_unaligned_fu_88_ap_start_reg;

assign or_ln24_fu_120_p2 = (resetMaximum6_dout | grp_fu_110_p2);

assign out_data_address1 = grp_tdf2_writeOutputs_unaligned_fu_88_out_data_address1;

assign out_data_ce1 = grp_tdf2_writeOutputs_unaligned_fu_88_out_data_ce1;

assign out_data_d1 = grp_tdf2_writeOutputs_unaligned_fu_88_out_data_d1;

assign out_data_we1 = grp_tdf2_writeOutputs_unaligned_fu_88_out_data_we1;

assign select_ln24_fu_126_p3 = ((or_ln24_fu_120_p2[0:0] == 1'b1) ? p_read : max_vals_4_0);

assign storeOutput7_read_read_fu_82_p2 = storeOutput7_dout;

endmodule //td_fused_top_tdf2_poolOutputs
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf2_readFilters24 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        filter_data_address0,
        filter_data_ce0,
        filter_data_q0,
        input_indices_23_dout,
        input_indices_23_empty_n,
        input_indices_23_read,
        weight_vecs_0_address0,
        weight_vecs_0_ce0,
        weight_vecs_0_we0,
        weight_vecs_0_d0
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state7 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [12:0] filter_data_address0;
output   filter_data_ce0;
input  [15:0] filter_data_q0;
input  [4:0] input_indices_23_dout;
input   input_indices_23_empty_n;
output   input_indices_23_read;
output  [7:0] weight_vecs_0_address0;
output   weight_vecs_0_ce0;
output   weight_vecs_0_we0;
output  [15:0] weight_vecs_0_d0;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg filter_data_ce0;
reg input_indices_23_read;
reg weight_vecs_0_ce0;
reg weight_vecs_0_we0;

reg    ap_done_reg;
  reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    input_indices_23_blk_n;
reg   [7:0] indvar_flatten13_reg_123;
reg   [1:0] ii_reg_134;
reg   [6:0] indvar_flatten_reg_145;
reg   [1:0] jj_reg_156;
reg   [4:0] kk_reg_167;
wire   [8:0] sext_ln47_fu_200_p1;
reg   [8:0] sext_ln47_reg_408;
wire   [7:0] add_ln47_5_fu_204_p2;
wire    ap_CS_fsm_pp0_stage0;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
wire    ap_block_state4_pp0_stage0_iter2;
wire    ap_block_state5_pp0_stage0_iter3;
wire    ap_block_state6_pp0_stage0_iter4;
wire    ap_block_pp0_stage0_11001;
wire   [0:0] icmp_ln47_fu_210_p2;
reg   [0:0] icmp_ln47_reg_418;
reg   [0:0] icmp_ln47_reg_418_pp0_iter1_reg;
reg   [0:0] icmp_ln47_reg_418_pp0_iter2_reg;
reg   [0:0] icmp_ln47_reg_418_pp0_iter3_reg;
wire   [0:0] icmp_ln48_fu_222_p2;
reg   [0:0] icmp_ln48_reg_422;
wire   [1:0] select_ln47_5_fu_228_p3;
reg   [1:0] select_ln47_5_reg_429;
wire   [6:0] select_ln48_10_fu_242_p3;
wire   [1:0] select_ln48_9_fu_329_p3;
reg   [1:0] select_ln48_9_reg_442;
reg    ap_enable_reg_pp0_iter1;
wire   [7:0] add_ln55_20_fu_392_p2;
reg   [7:0] add_ln55_20_reg_452;
reg   [7:0] add_ln55_20_reg_452_pp0_iter2_reg;
reg   [7:0] add_ln55_20_reg_452_pp0_iter3_reg;
wire   [4:0] add_ln49_fu_398_p2;
reg    ap_block_state1;
wire    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_flush_enable;
reg    ap_enable_reg_pp0_iter2;
reg    ap_condition_pp0_exit_iter1_state3;
reg    ap_enable_reg_pp0_iter3;
reg    ap_enable_reg_pp0_iter4;
reg   [1:0] ap_phi_mux_ii_phi_fu_138_p4;
wire    ap_block_pp0_stage0;
reg   [1:0] ap_phi_mux_jj_phi_fu_160_p4;
wire   [63:0] zext_ln55_47_fu_387_p1;
wire   [63:0] zext_ln55_48_fu_404_p1;
wire   [6:0] tmp_fu_182_p3;
wire   [7:0] zext_ln55_40_fu_190_p1;
wire   [7:0] zext_ln55_fu_178_p1;
wire   [7:0] sub_ln55_fu_194_p2;
wire   [1:0] add_ln47_fu_216_p2;
wire   [6:0] add_ln48_5_fu_236_p2;
wire   [8:0] zext_ln55_42_fu_260_p1;
wire   [8:0] add_ln55_fu_263_p2;
wire   [8:0] shl_ln55_fu_268_p2;
wire   [3:0] tmp_s_fu_280_p3;
wire   [3:0] zext_ln55_41_fu_257_p1;
wire   [0:0] icmp_ln49_fu_298_p2;
wire   [0:0] xor_ln47_fu_293_p2;
wire   [1:0] select_ln47_fu_250_p3;
wire   [0:0] and_ln47_fu_304_p2;
wire   [0:0] or_ln48_fu_316_p2;
wire   [1:0] add_ln48_fu_310_p2;
wire   [8:0] sub_ln55_9_fu_274_p2;
wire   [8:0] zext_ln55_44_fu_341_p1;
wire   [8:0] add_ln55_17_fu_345_p2;
wire   [3:0] sub_ln55_10_fu_287_p2;
wire   [3:0] zext_ln55_43_fu_337_p1;
wire   [3:0] add_ln55_18_fu_359_p2;
wire   [4:0] select_ln48_fu_321_p3;
wire   [12:0] tmp_124_cast_fu_351_p3;
wire   [12:0] zext_ln55_46_fu_377_p1;
wire   [12:0] add_ln55_19_fu_381_p2;
wire   [7:0] tmp_126_cast_fu_365_p3;
wire   [7:0] zext_ln55_45_fu_373_p1;
wire    ap_CS_fsm_state7;
reg   [2:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
#0 ap_enable_reg_pp0_iter4 = 1'b0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state7)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if ((1'b1 == ap_condition_pp0_flush_enable)) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((~((ap_start == 1'b0) | (input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            if ((1'b1 == ap_condition_pp0_exit_iter1_state3)) begin
                ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter0;
            end else if ((1'b1 == 1'b1)) begin
                ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
            end
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter4 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
        end else if ((~((ap_start == 1'b0) | (input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter4 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln47_reg_418 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ii_reg_134 <= select_ln47_5_reg_429;
    end else if ((~((ap_start == 1'b0) | (input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ii_reg_134 <= 2'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_fu_210_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        indvar_flatten13_reg_123 <= add_ln47_5_fu_204_p2;
    end else if ((~((ap_start == 1'b0) | (input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indvar_flatten13_reg_123 <= 8'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_fu_210_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        indvar_flatten_reg_145 <= select_ln48_10_fu_242_p3;
    end else if ((~((ap_start == 1'b0) | (input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indvar_flatten_reg_145 <= 7'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_reg_418_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        jj_reg_156 <= select_ln48_9_reg_442;
    end else if ((~((ap_start == 1'b0) | (input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        jj_reg_156 <= 2'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln47_reg_418 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        kk_reg_167 <= add_ln49_fu_398_p2;
    end else if ((~((ap_start == 1'b0) | (input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        kk_reg_167 <= 5'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_reg_418 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        add_ln55_20_reg_452 <= add_ln55_20_fu_392_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        add_ln55_20_reg_452_pp0_iter2_reg <= add_ln55_20_reg_452;
        add_ln55_20_reg_452_pp0_iter3_reg <= add_ln55_20_reg_452_pp0_iter2_reg;
        icmp_ln47_reg_418_pp0_iter2_reg <= icmp_ln47_reg_418_pp0_iter1_reg;
        icmp_ln47_reg_418_pp0_iter3_reg <= icmp_ln47_reg_418_pp0_iter2_reg;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln47_reg_418 <= icmp_ln47_fu_210_p2;
        icmp_ln47_reg_418_pp0_iter1_reg <= icmp_ln47_reg_418;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_fu_210_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln48_reg_422 <= icmp_ln48_fu_222_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_fu_210_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        select_ln47_5_reg_429 <= select_ln47_5_fu_228_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln47_reg_418 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        select_ln48_9_reg_442 <= select_ln48_9_fu_329_p3;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state1)) begin
        sext_ln47_reg_408 <= sext_ln47_fu_200_p1;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_condition_pp0_exit_iter1_state3 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter1_state3 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln47_fu_210_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_condition_pp0_flush_enable = 1'b1;
    end else begin
        ap_condition_pp0_flush_enable = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state7)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln47_reg_418 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_phi_mux_ii_phi_fu_138_p4 = select_ln47_5_reg_429;
    end else begin
        ap_phi_mux_ii_phi_fu_138_p4 = ii_reg_134;
    end
end

always @ (*) begin
    if (((icmp_ln47_reg_418_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        ap_phi_mux_jj_phi_fu_160_p4 = select_ln48_9_reg_442;
    end else begin
        ap_phi_mux_jj_phi_fu_160_p4 = jj_reg_156;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state7)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter3 == 1'b1)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter4 == 1'b1)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1)))) begin
        filter_data_ce0 = 1'b1;
    end else begin
        filter_data_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        input_indices_23_blk_n = input_indices_23_empty_n;
    end else begin
        input_indices_23_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        input_indices_23_read = 1'b1;
    end else begin
        input_indices_23_read = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter4 == 1'b1))) begin
        weight_vecs_0_ce0 = 1'b1;
    end else begin
        weight_vecs_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln47_reg_418_pp0_iter3_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter4 == 1'b1))) begin
        weight_vecs_0_we0 = 1'b1;
    end else begin
        weight_vecs_0_we0 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_start == 1'b0) | (input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((~((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b0)) & ~((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter4 == 1'b1) & (ap_enable_reg_pp0_iter3 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if ((((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b0)) | ((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter4 == 1'b1) & (ap_enable_reg_pp0_iter3 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_state7;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state7 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln47_5_fu_204_p2 = (indvar_flatten13_reg_123 + 8'd1);

assign add_ln47_fu_216_p2 = (ap_phi_mux_ii_phi_fu_138_p4 + 2'd1);

assign add_ln48_5_fu_236_p2 = (indvar_flatten_reg_145 + 7'd1);

assign add_ln48_fu_310_p2 = (select_ln47_fu_250_p3 + 2'd1);

assign add_ln49_fu_398_p2 = (select_ln48_fu_321_p3 + 5'd1);

assign add_ln55_17_fu_345_p2 = (sub_ln55_9_fu_274_p2 + zext_ln55_44_fu_341_p1);

assign add_ln55_18_fu_359_p2 = (sub_ln55_10_fu_287_p2 + zext_ln55_43_fu_337_p1);

assign add_ln55_19_fu_381_p2 = (tmp_124_cast_fu_351_p3 + zext_ln55_46_fu_377_p1);

assign add_ln55_20_fu_392_p2 = (tmp_126_cast_fu_365_p3 + zext_ln55_45_fu_373_p1);

assign add_ln55_fu_263_p2 = ((sext_ln47_reg_408) + (zext_ln55_42_fu_260_p1));

assign and_ln47_fu_304_p2 = (xor_ln47_fu_293_p2 & icmp_ln49_fu_298_p2);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state7 = ap_CS_fsm[32'd2];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1));
end

assign ap_block_state2_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter4 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign filter_data_address0 = zext_ln55_47_fu_387_p1;

assign icmp_ln47_fu_210_p2 = ((indvar_flatten13_reg_123 == 8'd144) ? 1'b1 : 1'b0);

assign icmp_ln48_fu_222_p2 = ((indvar_flatten_reg_145 == 7'd48) ? 1'b1 : 1'b0);

assign icmp_ln49_fu_298_p2 = ((kk_reg_167 == 5'd16) ? 1'b1 : 1'b0);

assign or_ln48_fu_316_p2 = (icmp_ln48_reg_422 | and_ln47_fu_304_p2);

assign select_ln47_5_fu_228_p3 = ((icmp_ln48_fu_222_p2[0:0] == 1'b1) ? add_ln47_fu_216_p2 : ap_phi_mux_ii_phi_fu_138_p4);

assign select_ln47_fu_250_p3 = ((icmp_ln48_reg_422[0:0] == 1'b1) ? 2'd0 : ap_phi_mux_jj_phi_fu_160_p4);

assign select_ln48_10_fu_242_p3 = ((icmp_ln48_fu_222_p2[0:0] == 1'b1) ? 7'd1 : add_ln48_5_fu_236_p2);

assign select_ln48_9_fu_329_p3 = ((and_ln47_fu_304_p2[0:0] == 1'b1) ? add_ln48_fu_310_p2 : select_ln47_fu_250_p3);

assign select_ln48_fu_321_p3 = ((or_ln48_fu_316_p2[0:0] == 1'b1) ? 5'd0 : kk_reg_167);

assign sext_ln47_fu_200_p1 = (sub_ln55_fu_194_p2);

assign shl_ln55_fu_268_p2 = add_ln55_fu_263_p2 << 9'd2;

assign sub_ln55_10_fu_287_p2 = (tmp_s_fu_280_p3 - zext_ln55_41_fu_257_p1);

assign sub_ln55_9_fu_274_p2 = (shl_ln55_fu_268_p2 - add_ln55_fu_263_p2);

assign sub_ln55_fu_194_p2 = (zext_ln55_40_fu_190_p1 - zext_ln55_fu_178_p1);

assign tmp_124_cast_fu_351_p3 = {{add_ln55_17_fu_345_p2}, {4'd0}};

assign tmp_126_cast_fu_365_p3 = {{add_ln55_18_fu_359_p2}, {4'd0}};

assign tmp_fu_182_p3 = {{input_indices_23_dout}, {2'd0}};

assign tmp_s_fu_280_p3 = {{select_ln47_5_reg_429}, {2'd0}};

assign weight_vecs_0_address0 = zext_ln55_48_fu_404_p1;

assign weight_vecs_0_d0 = filter_data_q0;

assign xor_ln47_fu_293_p2 = (icmp_ln48_reg_422 ^ 1'd1);

assign zext_ln55_40_fu_190_p1 = tmp_fu_182_p3;

assign zext_ln55_41_fu_257_p1 = select_ln47_5_reg_429;

assign zext_ln55_42_fu_260_p1 = select_ln47_5_reg_429;

assign zext_ln55_43_fu_337_p1 = select_ln48_9_fu_329_p3;

assign zext_ln55_44_fu_341_p1 = select_ln48_9_fu_329_p3;

assign zext_ln55_45_fu_373_p1 = select_ln48_fu_321_p3;

assign zext_ln55_46_fu_377_p1 = select_ln48_fu_321_p3;

assign zext_ln55_47_fu_387_p1 = add_ln55_19_fu_381_p2;

assign zext_ln55_48_fu_404_p1 = add_ln55_20_reg_452_pp0_iter3_reg;

assign zext_ln55_fu_178_p1 = input_indices_23_dout;

endmodule //td_fused_top_tdf2_readFilters24
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf2_readInputs25 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        in_data_address0,
        in_data_ce0,
        in_data_q0,
        i_17,
        j_17,
        ifmap_vec_address0,
        ifmap_vec_ce0,
        ifmap_vec_we0,
        ifmap_vec_d0,
        ifmap_vec_address1,
        ifmap_vec_ce1,
        ifmap_vec_we1,
        ifmap_vec_d1
);

parameter    ap_ST_fsm_state1 = 4'd1;
parameter    ap_ST_fsm_pp0_stage0 = 4'd2;
parameter    ap_ST_fsm_pp0_stage1 = 4'd4;
parameter    ap_ST_fsm_state8 = 4'd8;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [15:0] in_data_address0;
output   in_data_ce0;
input  [63:0] in_data_q0;
input  [15:0] i_17;
input  [15:0] j_17;
output  [7:0] ifmap_vec_address0;
output   ifmap_vec_ce0;
output   ifmap_vec_we0;
output  [15:0] ifmap_vec_d0;
output  [7:0] ifmap_vec_address1;
output   ifmap_vec_ce1;
output   ifmap_vec_we1;
output  [15:0] ifmap_vec_d1;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg in_data_ce0;
reg[7:0] ifmap_vec_address0;
reg ifmap_vec_ce0;
reg ifmap_vec_we0;
reg[15:0] ifmap_vec_d0;
reg[7:0] ifmap_vec_address1;
reg ifmap_vec_ce1;
reg ifmap_vec_we1;
reg[15:0] ifmap_vec_d1;

reg    ap_done_reg;
  reg   [3:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg   [5:0] indvar_flatten47_reg_194;
reg   [1:0] ii_reg_206;
reg   [4:0] indvar_flatten_reg_218;
reg   [1:0] jj_reg_229;
reg   [4:0] kk_0_i_reg_241;
wire   [17:0] p_cast_i_fu_270_p1;
reg   [17:0] p_cast_i_reg_931;
wire   [13:0] trunc_ln22_fu_274_p1;
reg   [13:0] trunc_ln22_reg_937;
wire   [17:0] sext_ln22_fu_284_p1;
reg   [17:0] sext_ln22_reg_943;
wire   [6:0] p_cast_fu_288_p2;
reg   [6:0] p_cast_reg_949;
wire   [0:0] or_ln23_21_fu_308_p2;
reg   [0:0] or_ln23_21_reg_955;
wire   [13:0] p_mid137_fu_314_p2;
reg   [13:0] p_mid137_reg_960;
wire   [6:0] p_cast5_i_fu_333_p2;
reg   [6:0] p_cast5_i_reg_965;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state4_pp0_stage0_iter1;
wire    ap_block_state6_pp0_stage0_iter2;
wire    ap_block_pp0_stage0_11001;
wire   [0:0] is_padding_fu_373_p2;
reg   [0:0] is_padding_reg_971;
wire   [0:0] icmp_ln19_fu_379_p2;
reg   [0:0] icmp_ln19_reg_978;
reg   [0:0] icmp_ln19_reg_978_pp0_iter1_reg;
reg   [0:0] icmp_ln19_reg_978_pp0_iter2_reg;
wire   [1:0] add_ln19_fu_385_p2;
reg   [1:0] add_ln19_reg_982;
wire   [0:0] icmp_ln20_fu_391_p2;
reg   [0:0] icmp_ln20_reg_987;
wire   [1:0] select_ln19_fu_397_p3;
reg   [1:0] select_ln19_reg_999;
wire   [6:0] p_cast5_i_mid1_fu_418_p2;
reg   [6:0] p_cast5_i_mid1_reg_1004;
wire   [0:0] or_ln23_23_fu_437_p2;
reg   [0:0] or_ln23_23_reg_1010;
wire   [1:0] add_ln20_fu_442_p2;
reg   [1:0] add_ln20_reg_1017;
wire   [0:0] or_ln23_25_fu_477_p2;
reg   [0:0] or_ln23_25_reg_1023;
wire   [4:0] add_ln20_5_fu_483_p2;
reg   [4:0] add_ln20_5_reg_1030;
wire   [5:0] add_ln19_5_fu_489_p2;
reg   [5:0] add_ln19_5_reg_1035;
wire    ap_CS_fsm_pp0_stage1;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_state3_pp0_stage1_iter0;
wire    ap_block_state5_pp0_stage1_iter1;
wire    ap_block_state7_pp0_stage1_iter2;
wire    ap_block_pp0_stage1_11001;
wire   [1:0] select_ln19_25_fu_527_p3;
reg   [1:0] select_ln19_25_reg_1040;
wire   [4:0] select_ln20_fu_591_p3;
reg   [4:0] select_ln20_reg_1047;
wire   [1:0] select_ln20_21_fu_599_p3;
reg   [1:0] select_ln20_21_reg_1053;
wire   [0:0] select_ln20_22_fu_608_p3;
reg   [0:0] select_ln20_22_reg_1059;
reg   [0:0] select_ln20_22_reg_1059_pp0_iter1_reg;
wire   [3:0] empty_111_fu_704_p1;
reg   [3:0] empty_111_reg_1067;
reg   [3:0] empty_111_reg_1067_pp0_iter1_reg;
wire   [4:0] select_ln20_25_fu_731_p3;
reg   [4:0] select_ln20_25_reg_1079;
wire   [4:0] add_ln25_fu_737_p2;
reg   [4:0] add_ln25_reg_1084;
reg    ap_enable_reg_pp0_iter1;
wire   [5:0] add_ln33_fu_769_p2;
reg   [5:0] add_ln33_reg_1089;
wire   [7:0] add_ln33_5_fu_790_p2;
reg   [7:0] add_ln33_5_reg_1096;
wire   [15:0] select_ln33_23_fu_869_p3;
reg   [15:0] select_ln33_23_reg_1101;
wire   [15:0] select_ln33_24_fu_890_p3;
reg   [15:0] select_ln33_24_reg_1106;
reg    ap_block_state1;
wire    ap_block_pp0_stage1_subdone;
reg    ap_condition_pp0_exit_iter0_state3;
reg    ap_enable_reg_pp0_iter2;
reg   [5:0] ap_phi_mux_indvar_flatten47_phi_fu_198_p4;
wire    ap_block_pp0_stage0;
reg   [1:0] ap_phi_mux_ii_phi_fu_210_p4;
reg   [4:0] ap_phi_mux_indvar_flatten_phi_fu_222_p4;
reg   [1:0] ap_phi_mux_jj_phi_fu_233_p4;
reg   [4:0] ap_phi_mux_kk_0_i_phi_fu_245_p4;
wire    ap_block_pp0_stage1;
wire   [63:0] sext_ln32_fu_726_p1;
wire   [63:0] zext_ln33_21_fu_796_p1;
wire   [63:0] sext_ln33_fu_828_p1;
wire   [63:0] sext_ln33_9_fu_909_p1;
wire   [63:0] sext_ln33_10_fu_926_p1;
wire   [15:0] select_ln33_fu_808_p3;
wire   [15:0] select_ln33_22_fu_847_p3;
wire   [16:0] zext_ln19_fu_256_p1;
wire   [16:0] empty_106_fu_264_p2;
wire   [16:0] j_cast_i_fu_252_p1;
wire   [16:0] add_ln22_fu_278_p2;
wire   [6:0] empty_fu_260_p1;
wire   [0:0] tmp_fu_294_p3;
wire   [0:0] icmp_ln24_fu_302_p2;
wire   [17:0] ii_cast_i_fu_320_p1;
wire   [6:0] ii_cast_fu_324_p1;
wire   [17:0] empty_107_fu_328_p2;
wire   [17:0] zext_ln20_fu_344_p1;
wire   [17:0] add_ln22_5_fu_348_p2;
wire   [0:0] tmp_37_fu_353_p3;
wire   [0:0] icmp_ln24_5_fu_361_p2;
wire   [0:0] or_ln23_fu_367_p2;
wire   [0:0] empty_108_fu_338_p2;
wire   [17:0] ii_cast_i_mid1_fu_405_p1;
wire   [6:0] ii_cast_mid1_fu_409_p1;
wire   [17:0] p_mid111_fu_413_p2;
wire   [0:0] p_mid113_fu_423_p2;
wire   [17:0] zext_ln20_5_fu_448_p1;
wire   [17:0] add_ln22_6_fu_452_p2;
wire   [0:0] tmp_38_fu_457_p3;
wire   [0:0] icmp_ln24_6_fu_465_p2;
wire   [0:0] or_ln23_24_fu_471_p2;
wire   [0:0] select_ln19_27_fu_429_p3;
wire   [2:0] zext_ln22_fu_495_p1;
wire   [2:0] tmp2_fu_505_p2;
wire   [13:0] tmp2_cast_fu_511_p1;
wire   [13:0] empty_109_fu_515_p2;
wire   [6:0] row_coord_int_mid131_fu_543_p3;
wire   [6:0] row_coord_int_fu_499_p3;
wire   [13:0] col_coord_int_mid139_fu_549_p3;
wire   [13:0] col_coord_int_fu_520_p3;
wire   [0:0] icmp_ln25_fu_574_p2;
wire   [0:0] xor_ln19_fu_569_p2;
wire   [0:0] and_ln19_fu_580_p2;
wire   [0:0] or_ln20_fu_586_p2;
wire   [0:0] select_ln19_28_fu_538_p3;
wire   [6:0] select_ln19_26_fu_533_p3;
wire   [2:0] zext_ln22_5_fu_605_p1;
wire   [2:0] tmp2_mid1_fu_622_p2;
wire   [13:0] tmp2_cast_mid1_fu_628_p1;
wire   [13:0] p_mid1_fu_632_p2;
wire   [6:0] row_coord_int_mid1_fu_615_p3;
wire   [6:0] select_ln19_29_fu_555_p3;
wire   [6:0] select_ln20_23_fu_644_p3;
wire   [13:0] tmp_7_fu_652_p3;
wire   [10:0] tmp_8_fu_664_p3;
wire   [14:0] zext_ln32_fu_660_p1;
wire   [14:0] zext_ln32_22_fu_672_p1;
wire   [14:0] sub_ln32_fu_676_p2;
wire   [13:0] col_coord_int_mid1_fu_637_p3;
wire   [13:0] select_ln19_30_fu_562_p3;
wire   [13:0] select_ln20_24_fu_686_p3;
wire   [15:0] sext_ln20_fu_682_p1;
wire   [15:0] zext_ln32_23_fu_694_p1;
wire   [15:0] add_ln32_fu_698_p2;
wire   [1:0] lshr_ln_fu_708_p4;
wire   [17:0] tmp_39_fu_718_p3;
wire   [3:0] tmp_s_fu_745_p3;
wire   [4:0] zext_ln33_18_fu_752_p1;
wire   [4:0] zext_ln33_fu_742_p1;
wire   [4:0] sub_ln33_fu_756_p2;
wire   [5:0] sub_ln33_cast_fu_762_p1;
wire   [5:0] zext_ln33_19_fu_766_p1;
wire   [3:0] trunc_ln33_fu_775_p1;
wire   [7:0] tmp_113_cast_fu_779_p3;
wire   [7:0] zext_ln33_20_fu_787_p1;
wire   [15:0] trunc_ln32_fu_800_p1;
wire   [15:0] bitcast_ln32_fu_804_p1;
wire   [3:0] or_ln25_fu_816_p2;
wire   [9:0] tmp_40_fu_821_p3;
wire   [15:0] tmp_66_i_fu_833_p4;
wire   [15:0] bitcast_ln32_22_fu_843_p1;
wire   [15:0] tmp_67_i_fu_855_p4;
wire   [15:0] bitcast_ln32_23_fu_865_p1;
wire   [15:0] tmp_68_i_fu_876_p4;
wire   [15:0] bitcast_ln32_24_fu_886_p1;
wire   [3:0] or_ln25_15_fu_897_p2;
wire   [9:0] tmp_41_fu_902_p3;
wire   [3:0] or_ln25_16_fu_914_p2;
wire   [9:0] tmp_42_fu_919_p3;
wire    ap_CS_fsm_state8;
reg   [3:0] ap_NS_fsm;
wire    ap_block_pp0_stage0_subdone;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 4'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_condition_pp0_exit_iter0_state3) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            if ((1'b1 == ap_condition_pp0_exit_iter0_state3)) begin
                ap_enable_reg_pp0_iter1 <= (1'b1 ^ ap_condition_pp0_exit_iter0_state3);
            end else if ((1'b1 == 1'b1)) begin
                ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
            end
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter2 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln19_reg_978 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ii_reg_206 <= select_ln19_25_reg_1040;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ii_reg_206 <= 2'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln19_reg_978 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        indvar_flatten47_reg_194 <= add_ln19_5_reg_1035;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indvar_flatten47_reg_194 <= 6'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln19_reg_978 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        indvar_flatten_reg_218 <= select_ln20_25_reg_1079;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indvar_flatten_reg_218 <= 5'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln19_reg_978 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        jj_reg_229 <= select_ln20_21_reg_1053;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        jj_reg_229 <= 2'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln19_reg_978_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        kk_0_i_reg_241 <= add_ln25_reg_1084;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        kk_0_i_reg_241 <= 5'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
        add_ln19_5_reg_1035 <= add_ln19_5_fu_489_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln19_fu_379_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        add_ln19_reg_982 <= add_ln19_fu_385_p2;
        add_ln20_5_reg_1030 <= add_ln20_5_fu_483_p2;
        add_ln20_reg_1017 <= add_ln20_fu_442_p2;
        icmp_ln20_reg_987 <= icmp_ln20_fu_391_p2;
        or_ln23_23_reg_1010 <= or_ln23_23_fu_437_p2;
        or_ln23_25_reg_1023 <= or_ln23_25_fu_477_p2;
        p_cast5_i_mid1_reg_1004 <= p_cast5_i_mid1_fu_418_p2;
        select_ln19_reg_999 <= select_ln19_fu_397_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln19_reg_978 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        add_ln25_reg_1084 <= add_ln25_fu_737_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln19_reg_978_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
        add_ln33_5_reg_1096 <= add_ln33_5_fu_790_p2;
        add_ln33_reg_1089 <= add_ln33_fu_769_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln19_reg_978 == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
        empty_111_reg_1067 <= empty_111_fu_704_p1;
        select_ln20_22_reg_1059 <= select_ln20_22_fu_608_p3;
        select_ln20_reg_1047 <= select_ln20_fu_591_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
        empty_111_reg_1067_pp0_iter1_reg <= empty_111_reg_1067;
        select_ln20_22_reg_1059_pp0_iter1_reg <= select_ln20_22_reg_1059;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln19_reg_978 <= icmp_ln19_fu_379_p2;
        icmp_ln19_reg_978_pp0_iter1_reg <= icmp_ln19_reg_978;
        icmp_ln19_reg_978_pp0_iter2_reg <= icmp_ln19_reg_978_pp0_iter1_reg;
        is_padding_reg_971 <= is_padding_fu_373_p2;
        p_cast5_i_reg_965 <= p_cast5_i_fu_333_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state1)) begin
        or_ln23_21_reg_955 <= or_ln23_21_fu_308_p2;
        p_cast_i_reg_931 <= p_cast_i_fu_270_p1;
        p_cast_reg_949 <= p_cast_fu_288_p2;
        p_mid137_reg_960 <= p_mid137_fu_314_p2;
        sext_ln22_reg_943 <= sext_ln22_fu_284_p1;
        trunc_ln22_reg_937 <= trunc_ln22_fu_274_p1;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln19_reg_978 == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
        select_ln19_25_reg_1040 <= select_ln19_25_fu_527_p3;
        select_ln20_21_reg_1053 <= select_ln20_21_fu_599_p3;
        select_ln20_25_reg_1079 <= select_ln20_25_fu_731_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln19_reg_978_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        select_ln33_23_reg_1101 <= select_ln33_23_fu_869_p3;
        select_ln33_24_reg_1106 <= select_ln33_24_fu_890_p3;
    end
end

always @ (*) begin
    if ((icmp_ln19_reg_978 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state3 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state3 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state8)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln19_reg_978 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_ii_phi_fu_210_p4 = select_ln19_25_reg_1040;
    end else begin
        ap_phi_mux_ii_phi_fu_210_p4 = ii_reg_206;
    end
end

always @ (*) begin
    if (((icmp_ln19_reg_978 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_indvar_flatten47_phi_fu_198_p4 = add_ln19_5_reg_1035;
    end else begin
        ap_phi_mux_indvar_flatten47_phi_fu_198_p4 = indvar_flatten47_reg_194;
    end
end

always @ (*) begin
    if (((icmp_ln19_reg_978 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_indvar_flatten_phi_fu_222_p4 = select_ln20_25_reg_1079;
    end else begin
        ap_phi_mux_indvar_flatten_phi_fu_222_p4 = indvar_flatten_reg_218;
    end
end

always @ (*) begin
    if (((icmp_ln19_reg_978 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_jj_phi_fu_233_p4 = select_ln20_21_reg_1053;
    end else begin
        ap_phi_mux_jj_phi_fu_233_p4 = jj_reg_229;
    end
end

always @ (*) begin
    if (((icmp_ln19_reg_978_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_kk_0_i_phi_fu_245_p4 = add_ln25_reg_1084;
    end else begin
        ap_phi_mux_kk_0_i_phi_fu_245_p4 = kk_0_i_reg_241;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state8)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((ap_enable_reg_pp0_iter2 == 1'b1)) begin
        if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            ifmap_vec_address0 = sext_ln33_10_fu_926_p1;
        end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ifmap_vec_address0 = sext_ln33_fu_828_p1;
        end else begin
            ifmap_vec_address0 = 'bx;
        end
    end else begin
        ifmap_vec_address0 = 'bx;
    end
end

always @ (*) begin
    if ((ap_enable_reg_pp0_iter2 == 1'b1)) begin
        if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            ifmap_vec_address1 = sext_ln33_9_fu_909_p1;
        end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ifmap_vec_address1 = zext_ln33_21_fu_796_p1;
        end else begin
            ifmap_vec_address1 = 'bx;
        end
    end else begin
        ifmap_vec_address1 = 'bx;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1)) | ((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter2 == 1'b1)))) begin
        ifmap_vec_ce0 = 1'b1;
    end else begin
        ifmap_vec_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1)) | ((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter2 == 1'b1)))) begin
        ifmap_vec_ce1 = 1'b1;
    end else begin
        ifmap_vec_ce1 = 1'b0;
    end
end

always @ (*) begin
    if ((ap_enable_reg_pp0_iter2 == 1'b1)) begin
        if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            ifmap_vec_d0 = select_ln33_24_reg_1106;
        end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ifmap_vec_d0 = select_ln33_22_fu_847_p3;
        end else begin
            ifmap_vec_d0 = 'bx;
        end
    end else begin
        ifmap_vec_d0 = 'bx;
    end
end

always @ (*) begin
    if ((ap_enable_reg_pp0_iter2 == 1'b1)) begin
        if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            ifmap_vec_d1 = select_ln33_23_reg_1101;
        end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ifmap_vec_d1 = select_ln33_fu_808_p3;
        end else begin
            ifmap_vec_d1 = 'bx;
        end
    end else begin
        ifmap_vec_d1 = 'bx;
    end
end

always @ (*) begin
    if ((((icmp_ln19_reg_978_pp0_iter2_reg == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter2 == 1'b1)) | ((icmp_ln19_reg_978_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1)))) begin
        ifmap_vec_we0 = 1'b1;
    end else begin
        ifmap_vec_we0 = 1'b0;
    end
end

always @ (*) begin
    if ((((icmp_ln19_reg_978_pp0_iter2_reg == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter2 == 1'b1)) | ((icmp_ln19_reg_978_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1)))) begin
        ifmap_vec_we1 = 1'b1;
    end else begin
        ifmap_vec_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1)) | ((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1)) | ((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1)) | ((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1)))) begin
        in_data_ce0 = 1'b1;
    end else begin
        in_data_ce0 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_pp0_stage1 : begin
            if ((~((icmp_ln19_reg_978 == 1'd1) & (1'b0 == ap_block_pp0_stage1_subdone) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1)) & ~((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter2 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0)) & (1'b0 == ap_block_pp0_stage1_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if ((((icmp_ln19_reg_978 == 1'd1) & (1'b0 == ap_block_pp0_stage1_subdone) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1)) | ((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter2 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_state8;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end
        end
        ap_ST_fsm_state8 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln19_5_fu_489_p2 = (indvar_flatten47_reg_194 + 6'd1);

assign add_ln19_fu_385_p2 = (ap_phi_mux_ii_phi_fu_210_p4 + 2'd1);

assign add_ln20_5_fu_483_p2 = (ap_phi_mux_indvar_flatten_phi_fu_222_p4 + 5'd1);

assign add_ln20_fu_442_p2 = (select_ln19_fu_397_p3 + 2'd1);

assign add_ln22_5_fu_348_p2 = ((sext_ln22_reg_943) + (zext_ln20_fu_344_p1));

assign add_ln22_6_fu_452_p2 = ((sext_ln22_reg_943) + (zext_ln20_5_fu_448_p1));

assign add_ln22_fu_278_p2 = ((j_cast_i_fu_252_p1) + (17'd131071));

assign add_ln25_fu_737_p2 = (select_ln20_reg_1047 + 5'd4);

assign add_ln32_fu_698_p2 = ((sext_ln20_fu_682_p1) + (zext_ln32_23_fu_694_p1));

assign add_ln33_5_fu_790_p2 = (tmp_113_cast_fu_779_p3 + zext_ln33_20_fu_787_p1);

assign add_ln33_fu_769_p2 = ((sub_ln33_cast_fu_762_p1) + (zext_ln33_19_fu_766_p1));

assign and_ln19_fu_580_p2 = (xor_ln19_fu_569_p2 & icmp_ln25_fu_574_p2);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_pp0_stage1 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state8 = ap_CS_fsm[32'd3];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (ap_done_reg == 1'b1));
end

assign ap_block_state2_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage1_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage1_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage1_iter2 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign bitcast_ln32_22_fu_843_p1 = tmp_66_i_fu_833_p4;

assign bitcast_ln32_23_fu_865_p1 = tmp_67_i_fu_855_p4;

assign bitcast_ln32_24_fu_886_p1 = tmp_68_i_fu_876_p4;

assign bitcast_ln32_fu_804_p1 = trunc_ln32_fu_800_p1;

assign col_coord_int_fu_520_p3 = ((is_padding_reg_971[0:0] == 1'b1) ? 14'd0 : empty_109_fu_515_p2);

assign col_coord_int_mid139_fu_549_p3 = ((or_ln23_23_reg_1010[0:0] == 1'b1) ? 14'd0 : p_mid137_reg_960);

assign col_coord_int_mid1_fu_637_p3 = ((or_ln23_25_reg_1023[0:0] == 1'b1) ? 14'd0 : p_mid1_fu_632_p2);

assign empty_106_fu_264_p2 = ((zext_ln19_fu_256_p1) + (17'd131071));

assign empty_107_fu_328_p2 = ((p_cast_i_reg_931) + (ii_cast_i_fu_320_p1));

assign empty_108_fu_338_p2 = ((empty_107_fu_328_p2 > 18'd111) ? 1'b1 : 1'b0);

assign empty_109_fu_515_p2 = ((tmp2_cast_fu_511_p1) + (trunc_ln22_reg_937));

assign empty_111_fu_704_p1 = select_ln20_fu_591_p3[3:0];

assign empty_fu_260_p1 = i_17[6:0];

assign icmp_ln19_fu_379_p2 = ((ap_phi_mux_indvar_flatten47_phi_fu_198_p4 == 6'd36) ? 1'b1 : 1'b0);

assign icmp_ln20_fu_391_p2 = ((ap_phi_mux_indvar_flatten_phi_fu_222_p4 == 5'd12) ? 1'b1 : 1'b0);

assign icmp_ln24_5_fu_361_p2 = (((add_ln22_5_fu_348_p2) > (18'd111)) ? 1'b1 : 1'b0);

assign icmp_ln24_6_fu_465_p2 = (((add_ln22_6_fu_452_p2) > (18'd111)) ? 1'b1 : 1'b0);

assign icmp_ln24_fu_302_p2 = (((add_ln22_fu_278_p2) > (17'd111)) ? 1'b1 : 1'b0);

assign icmp_ln25_fu_574_p2 = ((ap_phi_mux_kk_0_i_phi_fu_245_p4 == 5'd16) ? 1'b1 : 1'b0);

assign ii_cast_fu_324_p1 = ap_phi_mux_ii_phi_fu_210_p4;

assign ii_cast_i_fu_320_p1 = ap_phi_mux_ii_phi_fu_210_p4;

assign ii_cast_i_mid1_fu_405_p1 = add_ln19_fu_385_p2;

assign ii_cast_mid1_fu_409_p1 = add_ln19_fu_385_p2;

assign in_data_address0 = sext_ln32_fu_726_p1;

assign is_padding_fu_373_p2 = (or_ln23_fu_367_p2 | empty_108_fu_338_p2);

assign j_cast_i_fu_252_p1 = j_17;

assign lshr_ln_fu_708_p4 = {{select_ln20_fu_591_p3[3:2]}};

assign or_ln20_fu_586_p2 = (icmp_ln20_reg_987 | and_ln19_fu_580_p2);

assign or_ln23_21_fu_308_p2 = (tmp_fu_294_p3 | icmp_ln24_fu_302_p2);

assign or_ln23_23_fu_437_p2 = (p_mid113_fu_423_p2 | or_ln23_21_reg_955);

assign or_ln23_24_fu_471_p2 = (tmp_38_fu_457_p3 | icmp_ln24_6_fu_465_p2);

assign or_ln23_25_fu_477_p2 = (select_ln19_27_fu_429_p3 | or_ln23_24_fu_471_p2);

assign or_ln23_fu_367_p2 = (tmp_37_fu_353_p3 | icmp_ln24_5_fu_361_p2);

assign or_ln25_15_fu_897_p2 = (empty_111_reg_1067_pp0_iter1_reg | 4'd2);

assign or_ln25_16_fu_914_p2 = (empty_111_reg_1067_pp0_iter1_reg | 4'd3);

assign or_ln25_fu_816_p2 = (empty_111_reg_1067_pp0_iter1_reg | 4'd1);

assign p_cast5_i_fu_333_p2 = (p_cast_reg_949 + ii_cast_fu_324_p1);

assign p_cast5_i_mid1_fu_418_p2 = (p_cast_reg_949 + ii_cast_mid1_fu_409_p1);

assign p_cast_fu_288_p2 = ((empty_fu_260_p1) + (7'd127));

assign p_cast_i_fu_270_p1 = (empty_106_fu_264_p2);

assign p_mid111_fu_413_p2 = ((p_cast_i_reg_931) + (ii_cast_i_mid1_fu_405_p1));

assign p_mid113_fu_423_p2 = ((p_mid111_fu_413_p2 > 18'd111) ? 1'b1 : 1'b0);

assign p_mid137_fu_314_p2 = ((trunc_ln22_fu_274_p1) + (14'd16383));

assign p_mid1_fu_632_p2 = ((tmp2_cast_mid1_fu_628_p1) + (trunc_ln22_reg_937));

assign row_coord_int_fu_499_p3 = ((is_padding_reg_971[0:0] == 1'b1) ? 7'd0 : p_cast5_i_reg_965);

assign row_coord_int_mid131_fu_543_p3 = ((or_ln23_23_reg_1010[0:0] == 1'b1) ? 7'd0 : p_cast5_i_mid1_reg_1004);

assign row_coord_int_mid1_fu_615_p3 = ((or_ln23_25_reg_1023[0:0] == 1'b1) ? 7'd0 : select_ln19_26_fu_533_p3);

assign select_ln19_25_fu_527_p3 = ((icmp_ln20_reg_987[0:0] == 1'b1) ? add_ln19_reg_982 : ii_reg_206);

assign select_ln19_26_fu_533_p3 = ((icmp_ln20_reg_987[0:0] == 1'b1) ? p_cast5_i_mid1_reg_1004 : p_cast5_i_reg_965);

assign select_ln19_27_fu_429_p3 = ((icmp_ln20_fu_391_p2[0:0] == 1'b1) ? p_mid113_fu_423_p2 : empty_108_fu_338_p2);

assign select_ln19_28_fu_538_p3 = ((icmp_ln20_reg_987[0:0] == 1'b1) ? or_ln23_23_reg_1010 : is_padding_reg_971);

assign select_ln19_29_fu_555_p3 = ((icmp_ln20_reg_987[0:0] == 1'b1) ? row_coord_int_mid131_fu_543_p3 : row_coord_int_fu_499_p3);

assign select_ln19_30_fu_562_p3 = ((icmp_ln20_reg_987[0:0] == 1'b1) ? col_coord_int_mid139_fu_549_p3 : col_coord_int_fu_520_p3);

assign select_ln19_fu_397_p3 = ((icmp_ln20_fu_391_p2[0:0] == 1'b1) ? 2'd0 : ap_phi_mux_jj_phi_fu_233_p4);

assign select_ln20_21_fu_599_p3 = ((and_ln19_fu_580_p2[0:0] == 1'b1) ? add_ln20_reg_1017 : select_ln19_reg_999);

assign select_ln20_22_fu_608_p3 = ((and_ln19_fu_580_p2[0:0] == 1'b1) ? or_ln23_25_reg_1023 : select_ln19_28_fu_538_p3);

assign select_ln20_23_fu_644_p3 = ((and_ln19_fu_580_p2[0:0] == 1'b1) ? row_coord_int_mid1_fu_615_p3 : select_ln19_29_fu_555_p3);

assign select_ln20_24_fu_686_p3 = ((and_ln19_fu_580_p2[0:0] == 1'b1) ? col_coord_int_mid1_fu_637_p3 : select_ln19_30_fu_562_p3);

assign select_ln20_25_fu_731_p3 = ((icmp_ln20_reg_987[0:0] == 1'b1) ? 5'd1 : add_ln20_5_reg_1030);

assign select_ln20_fu_591_p3 = ((or_ln20_fu_586_p2[0:0] == 1'b1) ? 5'd0 : ap_phi_mux_kk_0_i_phi_fu_245_p4);

assign select_ln33_22_fu_847_p3 = ((select_ln20_22_reg_1059_pp0_iter1_reg[0:0] == 1'b1) ? 16'd0 : bitcast_ln32_22_fu_843_p1);

assign select_ln33_23_fu_869_p3 = ((select_ln20_22_reg_1059_pp0_iter1_reg[0:0] == 1'b1) ? 16'd0 : bitcast_ln32_23_fu_865_p1);

assign select_ln33_24_fu_890_p3 = ((select_ln20_22_reg_1059_pp0_iter1_reg[0:0] == 1'b1) ? 16'd0 : bitcast_ln32_24_fu_886_p1);

assign select_ln33_fu_808_p3 = ((select_ln20_22_reg_1059_pp0_iter1_reg[0:0] == 1'b1) ? 16'd0 : bitcast_ln32_fu_804_p1);

assign sext_ln20_fu_682_p1 = (sub_ln32_fu_676_p2);

assign sext_ln22_fu_284_p1 = add_ln22_fu_278_p2;

assign sext_ln32_fu_726_p1 = (tmp_39_fu_718_p3);

assign sext_ln33_10_fu_926_p1 = (tmp_42_fu_919_p3);

assign sext_ln33_9_fu_909_p1 = (tmp_41_fu_902_p3);

assign sext_ln33_fu_828_p1 = (tmp_40_fu_821_p3);

assign sub_ln32_fu_676_p2 = (zext_ln32_fu_660_p1 - zext_ln32_22_fu_672_p1);

assign sub_ln33_cast_fu_762_p1 = (sub_ln33_fu_756_p2);

assign sub_ln33_fu_756_p2 = (zext_ln33_18_fu_752_p1 - zext_ln33_fu_742_p1);

assign tmp2_cast_fu_511_p1 = (tmp2_fu_505_p2);

assign tmp2_cast_mid1_fu_628_p1 = (tmp2_mid1_fu_622_p2);

assign tmp2_fu_505_p2 = ((zext_ln22_fu_495_p1) + (3'd7));

assign tmp2_mid1_fu_622_p2 = ((zext_ln22_5_fu_605_p1) + (3'd7));

assign tmp_113_cast_fu_779_p3 = {{trunc_ln33_fu_775_p1}, {4'd0}};

assign tmp_37_fu_353_p3 = add_ln22_5_fu_348_p2[32'd17];

assign tmp_38_fu_457_p3 = add_ln22_6_fu_452_p2[32'd17];

assign tmp_39_fu_718_p3 = {{add_ln32_fu_698_p2}, {lshr_ln_fu_708_p4}};

assign tmp_40_fu_821_p3 = {{add_ln33_reg_1089}, {or_ln25_fu_816_p2}};

assign tmp_41_fu_902_p3 = {{add_ln33_reg_1089}, {or_ln25_15_fu_897_p2}};

assign tmp_42_fu_919_p3 = {{add_ln33_reg_1089}, {or_ln25_16_fu_914_p2}};

assign tmp_66_i_fu_833_p4 = {{in_data_q0[31:16]}};

assign tmp_67_i_fu_855_p4 = {{in_data_q0[47:32]}};

assign tmp_68_i_fu_876_p4 = {{in_data_q0[63:48]}};

assign tmp_7_fu_652_p3 = {{select_ln20_23_fu_644_p3}, {7'd0}};

assign tmp_8_fu_664_p3 = {{select_ln20_23_fu_644_p3}, {4'd0}};

assign tmp_fu_294_p3 = add_ln22_fu_278_p2[32'd16];

assign tmp_s_fu_745_p3 = {{select_ln19_25_reg_1040}, {2'd0}};

assign trunc_ln22_fu_274_p1 = j_17[13:0];

assign trunc_ln32_fu_800_p1 = in_data_q0[15:0];

assign trunc_ln33_fu_775_p1 = add_ln33_fu_769_p2[3:0];

assign xor_ln19_fu_569_p2 = (icmp_ln20_reg_987 ^ 1'd1);

assign zext_ln19_fu_256_p1 = i_17;

assign zext_ln20_5_fu_448_p1 = add_ln20_fu_442_p2;

assign zext_ln20_fu_344_p1 = ap_phi_mux_jj_phi_fu_233_p4;

assign zext_ln22_5_fu_605_p1 = add_ln20_reg_1017;

assign zext_ln22_fu_495_p1 = jj_reg_229;

assign zext_ln32_22_fu_672_p1 = tmp_8_fu_664_p3;

assign zext_ln32_23_fu_694_p1 = select_ln20_24_fu_686_p3;

assign zext_ln32_fu_660_p1 = tmp_7_fu_652_p3;

assign zext_ln33_18_fu_752_p1 = tmp_s_fu_745_p3;

assign zext_ln33_19_fu_766_p1 = select_ln20_21_reg_1053;

assign zext_ln33_20_fu_787_p1 = select_ln20_reg_1047;

assign zext_ln33_21_fu_796_p1 = add_ln33_5_reg_1096;

assign zext_ln33_fu_742_p1 = select_ln19_25_reg_1040;

endmodule //td_fused_top_tdf2_readInputs25
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf2_writeOutputs_unaligned (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        i,
        j,
        out_data_address1,
        out_data_ce1,
        out_data_we1,
        out_data_d1,
        max_vals_4_0
);

parameter    ap_ST_fsm_state1 = 2'd1;
parameter    ap_ST_fsm_state2 = 2'd2;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
input  [5:0] i;
input  [11:0] j;
output  [14:0] out_data_address1;
output   out_data_ce1;
output   out_data_we1;
output  [63:0] out_data_d1;
input  [15:0] max_vals_4_0;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg out_data_ce1;
reg out_data_we1;

  reg   [1:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg   [15:0] outputCount_7;
reg   [15:0] outputChanIdx_7;
reg   [15:0] outputRow_9_0;
reg   [15:0] outputRow_9_1;
reg   [15:0] outputRow_9_2;
reg   [15:0] outputRow_9_3;
wire   [15:0] add_ln87_fu_175_p2;
wire   [0:0] icmp_ln88_fu_181_p2;
reg   [0:0] icmp_ln88_reg_295;
reg   [15:0] ap_phi_mux_empty_phi_fu_92_p4;
reg   [15:0] empty_reg_89;
wire    ap_CS_fsm_state2;
wire   [63:0] zext_ln94_14_fu_209_p1;
wire   [15:0] select_ln97_fu_267_p3;
wire   [1:0] trunc_ln86_fu_147_p1;
reg   [15:0] ap_sig_allocacmp_outputRow_9_0_load;
reg   [15:0] ap_sig_allocacmp_outputRow_9_1_load;
reg   [15:0] ap_sig_allocacmp_outputRow_9_2_load;
reg   [15:0] ap_sig_allocacmp_outputRow_9_3_load;
wire   [8:0] tmp_s_fu_107_p3;
wire   [11:0] tmp_fu_99_p3;
wire   [11:0] zext_ln94_fu_115_p1;
wire   [11:0] sub_ln94_fu_119_p2;
wire   [11:0] add_ln94_fu_125_p2;
wire   [4:0] trunc_ln94_fu_195_p1;
wire   [14:0] tmp_110_cast_fu_131_p3;
wire   [14:0] zext_ln94_13_fu_199_p1;
wire   [14:0] add_ln94_6_fu_203_p2;
wire   [15:0] bitcast_ln94_18_fu_238_p1;
wire   [15:0] bitcast_ln94_17_fu_230_p1;
wire   [15:0] bitcast_ln94_16_fu_222_p1;
wire   [15:0] bitcast_ln94_fu_214_p1;
wire   [15:0] add_ln96_fu_255_p2;
wire   [0:0] icmp_ln97_fu_261_p2;
reg   [1:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_CS_fsm = 2'd1;
#0 outputCount_7 = 16'd0;
#0 outputChanIdx_7 = 16'd0;
#0 outputRow_9_0 = 16'd0;
#0 outputRow_9_1 = 16'd0;
#0 outputRow_9_2 = 16'd0;
#0 outputRow_9_3 = 16'd0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln88_reg_295 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        empty_reg_89 <= 16'd0;
    end else if (((ap_start == 1'b1) & (icmp_ln88_fu_181_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state1))) begin
        empty_reg_89 <= add_ln87_fu_175_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state1)) begin
        icmp_ln88_reg_295 <= icmp_ln88_fu_181_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_start == 1'b1) & (icmp_ln88_fu_181_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1))) begin
        outputChanIdx_7 <= select_ln97_fu_267_p3;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        outputCount_7 <= ap_phi_mux_empty_phi_fu_92_p4;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_start == 1'b1) & (trunc_ln86_fu_147_p1 == 2'd0) & (1'b1 == ap_CS_fsm_state1))) begin
        outputRow_9_0 <= max_vals_4_0;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_start == 1'b1) & (trunc_ln86_fu_147_p1 == 2'd1) & (1'b1 == ap_CS_fsm_state1))) begin
        outputRow_9_1 <= max_vals_4_0;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_start == 1'b1) & (trunc_ln86_fu_147_p1 == 2'd2) & (1'b1 == ap_CS_fsm_state1))) begin
        outputRow_9_2 <= max_vals_4_0;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_start == 1'b1) & (trunc_ln86_fu_147_p1 == 2'd3) & (1'b1 == ap_CS_fsm_state1))) begin
        outputRow_9_3 <= max_vals_4_0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state2) | ((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1)))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = 1'b0;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln88_reg_295 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        ap_phi_mux_empty_phi_fu_92_p4 = 16'd0;
    end else begin
        ap_phi_mux_empty_phi_fu_92_p4 = empty_reg_89;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((trunc_ln86_fu_147_p1 == 2'd0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_sig_allocacmp_outputRow_9_0_load = max_vals_4_0;
    end else begin
        ap_sig_allocacmp_outputRow_9_0_load = outputRow_9_0;
    end
end

always @ (*) begin
    if (((trunc_ln86_fu_147_p1 == 2'd1) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_sig_allocacmp_outputRow_9_1_load = max_vals_4_0;
    end else begin
        ap_sig_allocacmp_outputRow_9_1_load = outputRow_9_1;
    end
end

always @ (*) begin
    if (((trunc_ln86_fu_147_p1 == 2'd2) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_sig_allocacmp_outputRow_9_2_load = max_vals_4_0;
    end else begin
        ap_sig_allocacmp_outputRow_9_2_load = outputRow_9_2;
    end
end

always @ (*) begin
    if (((trunc_ln86_fu_147_p1 == 2'd3) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_sig_allocacmp_outputRow_9_3_load = max_vals_4_0;
    end else begin
        ap_sig_allocacmp_outputRow_9_3_load = outputRow_9_3;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state2) | ((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)))) begin
        out_data_ce1 = 1'b1;
    end else begin
        out_data_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_start == 1'b1) & (icmp_ln88_fu_181_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1))) begin
        out_data_we1 = 1'b1;
    end else begin
        out_data_we1 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_state2 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln87_fu_175_p2 = (outputCount_7 + 16'd1);

assign add_ln94_6_fu_203_p2 = (tmp_110_cast_fu_131_p3 + zext_ln94_13_fu_199_p1);

assign add_ln94_fu_125_p2 = (sub_ln94_fu_119_p2 + j);

assign add_ln96_fu_255_p2 = (outputChanIdx_7 + 16'd1);

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign bitcast_ln94_16_fu_222_p1 = ap_sig_allocacmp_outputRow_9_1_load;

assign bitcast_ln94_17_fu_230_p1 = ap_sig_allocacmp_outputRow_9_2_load;

assign bitcast_ln94_18_fu_238_p1 = ap_sig_allocacmp_outputRow_9_3_load;

assign bitcast_ln94_fu_214_p1 = ap_sig_allocacmp_outputRow_9_0_load;

assign icmp_ln88_fu_181_p2 = ((add_ln87_fu_175_p2 == 16'd4) ? 1'b1 : 1'b0);

assign icmp_ln97_fu_261_p2 = ((add_ln96_fu_255_p2 == 16'd8) ? 1'b1 : 1'b0);

assign out_data_address1 = zext_ln94_14_fu_209_p1;

assign out_data_d1 = {{{{bitcast_ln94_18_fu_238_p1}, {bitcast_ln94_17_fu_230_p1}}, {bitcast_ln94_16_fu_222_p1}}, {bitcast_ln94_fu_214_p1}};

assign select_ln97_fu_267_p3 = ((icmp_ln97_fu_261_p2[0:0] == 1'b1) ? 16'd0 : add_ln96_fu_255_p2);

assign sub_ln94_fu_119_p2 = (tmp_fu_99_p3 - zext_ln94_fu_115_p1);

assign tmp_110_cast_fu_131_p3 = {{add_ln94_fu_125_p2}, {3'd0}};

assign tmp_fu_99_p3 = {{i}, {6'd0}};

assign tmp_s_fu_107_p3 = {{i}, {3'd0}};

assign trunc_ln86_fu_147_p1 = outputCount_7[1:0];

assign trunc_ln94_fu_195_p1 = outputChanIdx_7[4:0];

assign zext_ln94_13_fu_199_p1 = trunc_ln94_fu_195_p1;

assign zext_ln94_14_fu_209_p1 = add_ln94_6_fu_203_p2;

assign zext_ln94_fu_115_p1 = tmp_s_fu_107_p3;

endmodule //td_fused_top_tdf2_writeOutputs_unaligned
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf3_112 (
        in_data_address0,
        in_data_ce0,
        in_data_d0,
        in_data_q0,
        in_data_we0,
        in_data_address1,
        in_data_ce1,
        in_data_d1,
        in_data_q1,
        in_data_we1,
        out_data_address0,
        out_data_ce0,
        out_data_d0,
        out_data_q0,
        out_data_we0,
        out_data_address1,
        out_data_ce1,
        out_data_d1,
        out_data_q1,
        out_data_we1,
        filter_data_address0,
        filter_data_ce0,
        filter_data_d0,
        filter_data_q0,
        filter_data_we0,
        filter_data_address1,
        filter_data_ce1,
        filter_data_d1,
        filter_data_q1,
        filter_data_we1,
        adjustments_address0,
        adjustments_ce0,
        adjustments_d0,
        adjustments_q0,
        adjustments_we0,
        adjustments_address1,
        adjustments_ce1,
        adjustments_d1,
        adjustments_q1,
        adjustments_we1,
        ap_clk,
        ap_rst,
        in_data_empty_n,
        in_data_read,
        out_data_full_n,
        out_data_write,
        ap_start,
        ap_done,
        ap_ready,
        ap_idle,
        ap_continue
);


output  [14:0] in_data_address0;
output   in_data_ce0;
output  [63:0] in_data_d0;
input  [63:0] in_data_q0;
output   in_data_we0;
output  [14:0] in_data_address1;
output   in_data_ce1;
output  [63:0] in_data_d1;
input  [63:0] in_data_q1;
output   in_data_we1;
output  [13:0] out_data_address0;
output   out_data_ce0;
output  [63:0] out_data_d0;
input  [63:0] out_data_q0;
output   out_data_we0;
output  [13:0] out_data_address1;
output   out_data_ce1;
output  [63:0] out_data_d1;
input  [63:0] out_data_q1;
output   out_data_we1;
output  [8:0] filter_data_address0;
output   filter_data_ce0;
output  [15:0] filter_data_d0;
input  [15:0] filter_data_q0;
output   filter_data_we0;
output  [8:0] filter_data_address1;
output   filter_data_ce1;
output  [15:0] filter_data_d1;
input  [15:0] filter_data_q1;
output   filter_data_we1;
output  [3:0] adjustments_address0;
output   adjustments_ce0;
output  [47:0] adjustments_d0;
input  [47:0] adjustments_q0;
output   adjustments_we0;
output  [3:0] adjustments_address1;
output   adjustments_ce1;
output  [47:0] adjustments_d1;
input  [47:0] adjustments_q1;
output   adjustments_we1;
input   ap_clk;
input   ap_rst;
input   in_data_empty_n;
output   in_data_read;
input   out_data_full_n;
output   out_data_write;
input   ap_start;
output   ap_done;
output   ap_ready;
output   ap_idle;
input   ap_continue;

reg ap_done;
reg ap_ready;
reg ap_idle;

wire   [14:0] dataflow_in_loop_TOP_LOOP37928_U0_in_data_address0;
wire    dataflow_in_loop_TOP_LOOP37928_U0_in_data_ce0;
wire   [63:0] dataflow_in_loop_TOP_LOOP37928_U0_in_data_d0;
wire    dataflow_in_loop_TOP_LOOP37928_U0_in_data_we0;
wire   [14:0] dataflow_in_loop_TOP_LOOP37928_U0_in_data_address1;
wire    dataflow_in_loop_TOP_LOOP37928_U0_in_data_ce1;
wire   [63:0] dataflow_in_loop_TOP_LOOP37928_U0_in_data_d1;
wire    dataflow_in_loop_TOP_LOOP37928_U0_in_data_we1;
wire   [8:0] dataflow_in_loop_TOP_LOOP37928_U0_filter_data_address0;
wire    dataflow_in_loop_TOP_LOOP37928_U0_filter_data_ce0;
wire   [15:0] dataflow_in_loop_TOP_LOOP37928_U0_filter_data_d0;
wire    dataflow_in_loop_TOP_LOOP37928_U0_filter_data_we0;
wire   [8:0] dataflow_in_loop_TOP_LOOP37928_U0_filter_data_address1;
wire    dataflow_in_loop_TOP_LOOP37928_U0_filter_data_ce1;
wire   [15:0] dataflow_in_loop_TOP_LOOP37928_U0_filter_data_d1;
wire    dataflow_in_loop_TOP_LOOP37928_U0_filter_data_we1;
wire   [3:0] dataflow_in_loop_TOP_LOOP37928_U0_adjustments_address0;
wire    dataflow_in_loop_TOP_LOOP37928_U0_adjustments_ce0;
wire   [47:0] dataflow_in_loop_TOP_LOOP37928_U0_adjustments_d0;
wire    dataflow_in_loop_TOP_LOOP37928_U0_adjustments_we0;
wire   [3:0] dataflow_in_loop_TOP_LOOP37928_U0_adjustments_address1;
wire    dataflow_in_loop_TOP_LOOP37928_U0_adjustments_ce1;
wire   [47:0] dataflow_in_loop_TOP_LOOP37928_U0_adjustments_d1;
wire    dataflow_in_loop_TOP_LOOP37928_U0_adjustments_we1;
wire   [13:0] dataflow_in_loop_TOP_LOOP37928_U0_out_data_address0;
wire    dataflow_in_loop_TOP_LOOP37928_U0_out_data_ce0;
wire   [63:0] dataflow_in_loop_TOP_LOOP37928_U0_out_data_d0;
wire    dataflow_in_loop_TOP_LOOP37928_U0_out_data_we0;
wire   [13:0] dataflow_in_loop_TOP_LOOP37928_U0_out_data_address1;
wire    dataflow_in_loop_TOP_LOOP37928_U0_out_data_ce1;
wire   [63:0] dataflow_in_loop_TOP_LOOP37928_U0_out_data_d1;
wire    dataflow_in_loop_TOP_LOOP37928_U0_out_data_we1;
wire    dataflow_in_loop_TOP_LOOP37928_U0_ap_start;
wire    dataflow_in_loop_TOP_LOOP37928_U0_in_data_read;
wire    dataflow_in_loop_TOP_LOOP37928_U0_out_data_write;
wire    dataflow_in_loop_TOP_LOOP37928_U0_ap_done;
wire    dataflow_in_loop_TOP_LOOP37928_U0_ap_ready;
wire    dataflow_in_loop_TOP_LOOP37928_U0_ap_idle;
reg    dataflow_in_loop_TOP_LOOP37928_U0_ap_continue;
wire    dataflow_in_loop_TOP_LOOP37928_U0_in_data_full_n;
wire    dataflow_in_loop_TOP_LOOP37928_U0_in_data_write;
wire    ap_sync_continue;
wire    ap_sync_done;
wire    ap_sync_ready;
reg   [15:0] loop_dataflow_input_count;
reg   [15:0] loop_dataflow_output_count;
wire   [15:0] bound_minus_1;
wire    dataflow_in_loop_TOP_LOOP37928_U0_start_full_n;
wire    dataflow_in_loop_TOP_LOOP37928_U0_start_write;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 loop_dataflow_input_count = 16'd0;
#0 loop_dataflow_output_count = 16'd0;
end

td_fused_top_dataflow_in_loop_TOP_LOOP37928 dataflow_in_loop_TOP_LOOP37928_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .in_data_address0(dataflow_in_loop_TOP_LOOP37928_U0_in_data_address0),
    .in_data_ce0(dataflow_in_loop_TOP_LOOP37928_U0_in_data_ce0),
    .in_data_d0(dataflow_in_loop_TOP_LOOP37928_U0_in_data_d0),
    .in_data_q0(in_data_q0),
    .in_data_we0(dataflow_in_loop_TOP_LOOP37928_U0_in_data_we0),
    .in_data_address1(dataflow_in_loop_TOP_LOOP37928_U0_in_data_address1),
    .in_data_ce1(dataflow_in_loop_TOP_LOOP37928_U0_in_data_ce1),
    .in_data_d1(dataflow_in_loop_TOP_LOOP37928_U0_in_data_d1),
    .in_data_q1(64'd0),
    .in_data_we1(dataflow_in_loop_TOP_LOOP37928_U0_in_data_we1),
    .filter_data_address0(dataflow_in_loop_TOP_LOOP37928_U0_filter_data_address0),
    .filter_data_ce0(dataflow_in_loop_TOP_LOOP37928_U0_filter_data_ce0),
    .filter_data_d0(dataflow_in_loop_TOP_LOOP37928_U0_filter_data_d0),
    .filter_data_q0(filter_data_q0),
    .filter_data_we0(dataflow_in_loop_TOP_LOOP37928_U0_filter_data_we0),
    .filter_data_address1(dataflow_in_loop_TOP_LOOP37928_U0_filter_data_address1),
    .filter_data_ce1(dataflow_in_loop_TOP_LOOP37928_U0_filter_data_ce1),
    .filter_data_d1(dataflow_in_loop_TOP_LOOP37928_U0_filter_data_d1),
    .filter_data_q1(16'd0),
    .filter_data_we1(dataflow_in_loop_TOP_LOOP37928_U0_filter_data_we1),
    .adjustments_address0(dataflow_in_loop_TOP_LOOP37928_U0_adjustments_address0),
    .adjustments_ce0(dataflow_in_loop_TOP_LOOP37928_U0_adjustments_ce0),
    .adjustments_d0(dataflow_in_loop_TOP_LOOP37928_U0_adjustments_d0),
    .adjustments_q0(adjustments_q0),
    .adjustments_we0(dataflow_in_loop_TOP_LOOP37928_U0_adjustments_we0),
    .adjustments_address1(dataflow_in_loop_TOP_LOOP37928_U0_adjustments_address1),
    .adjustments_ce1(dataflow_in_loop_TOP_LOOP37928_U0_adjustments_ce1),
    .adjustments_d1(dataflow_in_loop_TOP_LOOP37928_U0_adjustments_d1),
    .adjustments_q1(48'd0),
    .adjustments_we1(dataflow_in_loop_TOP_LOOP37928_U0_adjustments_we1),
    .out_data_address0(dataflow_in_loop_TOP_LOOP37928_U0_out_data_address0),
    .out_data_ce0(dataflow_in_loop_TOP_LOOP37928_U0_out_data_ce0),
    .out_data_d0(dataflow_in_loop_TOP_LOOP37928_U0_out_data_d0),
    .out_data_q0(64'd0),
    .out_data_we0(dataflow_in_loop_TOP_LOOP37928_U0_out_data_we0),
    .out_data_address1(dataflow_in_loop_TOP_LOOP37928_U0_out_data_address1),
    .out_data_ce1(dataflow_in_loop_TOP_LOOP37928_U0_out_data_ce1),
    .out_data_d1(dataflow_in_loop_TOP_LOOP37928_U0_out_data_d1),
    .out_data_q1(64'd0),
    .out_data_we1(dataflow_in_loop_TOP_LOOP37928_U0_out_data_we1),
    .ap_start(dataflow_in_loop_TOP_LOOP37928_U0_ap_start),
    .in_data_empty_n(1'b0),
    .in_data_read(dataflow_in_loop_TOP_LOOP37928_U0_in_data_read),
    .out_data_full_n(out_data_full_n),
    .out_data_write(dataflow_in_loop_TOP_LOOP37928_U0_out_data_write),
    .ap_done(dataflow_in_loop_TOP_LOOP37928_U0_ap_done),
    .ap_ready(dataflow_in_loop_TOP_LOOP37928_U0_ap_ready),
    .ap_idle(dataflow_in_loop_TOP_LOOP37928_U0_ap_idle),
    .ap_continue(dataflow_in_loop_TOP_LOOP37928_U0_ap_continue)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        loop_dataflow_input_count <= 16'd0;
    end else begin
        if ((~(loop_dataflow_input_count == bound_minus_1) & (dataflow_in_loop_TOP_LOOP37928_U0_ap_ready == 1'b1) & (ap_start == 1'b1))) begin
            loop_dataflow_input_count <= (loop_dataflow_input_count + 16'd1);
        end else if (((dataflow_in_loop_TOP_LOOP37928_U0_ap_ready == 1'b1) & (loop_dataflow_input_count == bound_minus_1) & (ap_start == 1'b1))) begin
            loop_dataflow_input_count <= 16'd0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        loop_dataflow_output_count <= 16'd0;
    end else begin
        if ((~(loop_dataflow_output_count == bound_minus_1) & (dataflow_in_loop_TOP_LOOP37928_U0_ap_done == 1'b1) & (dataflow_in_loop_TOP_LOOP37928_U0_ap_continue == 1'b1))) begin
            loop_dataflow_output_count <= (loop_dataflow_output_count + 16'd1);
        end else if (((dataflow_in_loop_TOP_LOOP37928_U0_ap_done == 1'b1) & (loop_dataflow_output_count == bound_minus_1) & (dataflow_in_loop_TOP_LOOP37928_U0_ap_continue == 1'b1))) begin
            loop_dataflow_output_count <= 16'd0;
        end
    end
end

always @ (*) begin
    if (((dataflow_in_loop_TOP_LOOP37928_U0_ap_done == 1'b1) & (loop_dataflow_output_count == bound_minus_1))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = 1'b0;
    end
end

always @ (*) begin
    if (((dataflow_in_loop_TOP_LOOP37928_U0_ap_idle == 1'b1) & (loop_dataflow_output_count == 16'd0) & (ap_start == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((dataflow_in_loop_TOP_LOOP37928_U0_ap_ready == 1'b1) & (loop_dataflow_input_count == bound_minus_1) & (ap_start == 1'b1))) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((~(loop_dataflow_output_count == bound_minus_1) | (ap_continue == 1'b1))) begin
        dataflow_in_loop_TOP_LOOP37928_U0_ap_continue = 1'b1;
    end else begin
        dataflow_in_loop_TOP_LOOP37928_U0_ap_continue = 1'b0;
    end
end

assign adjustments_address0 = dataflow_in_loop_TOP_LOOP37928_U0_adjustments_address0;

assign adjustments_address1 = 4'd0;

assign adjustments_ce0 = dataflow_in_loop_TOP_LOOP37928_U0_adjustments_ce0;

assign adjustments_ce1 = 1'b0;

assign adjustments_d0 = 48'd0;

assign adjustments_d1 = 48'd0;

assign adjustments_we0 = 1'b0;

assign adjustments_we1 = 1'b0;

assign ap_sync_continue = ap_continue;

assign ap_sync_done = dataflow_in_loop_TOP_LOOP37928_U0_ap_done;

assign ap_sync_ready = dataflow_in_loop_TOP_LOOP37928_U0_ap_ready;

assign bound_minus_1 = (16'd50176 - 16'd1);

assign dataflow_in_loop_TOP_LOOP37928_U0_ap_start = ap_start;

assign dataflow_in_loop_TOP_LOOP37928_U0_in_data_full_n = in_data_empty_n;

assign dataflow_in_loop_TOP_LOOP37928_U0_in_data_write = 1'b0;

assign dataflow_in_loop_TOP_LOOP37928_U0_start_full_n = 1'b1;

assign dataflow_in_loop_TOP_LOOP37928_U0_start_write = 1'b0;

assign filter_data_address0 = dataflow_in_loop_TOP_LOOP37928_U0_filter_data_address0;

assign filter_data_address1 = 9'd0;

assign filter_data_ce0 = dataflow_in_loop_TOP_LOOP37928_U0_filter_data_ce0;

assign filter_data_ce1 = 1'b0;

assign filter_data_d0 = 16'd0;

assign filter_data_d1 = 16'd0;

assign filter_data_we0 = 1'b0;

assign filter_data_we1 = 1'b0;

assign in_data_address0 = dataflow_in_loop_TOP_LOOP37928_U0_in_data_address0;

assign in_data_address1 = 15'd0;

assign in_data_ce0 = dataflow_in_loop_TOP_LOOP37928_U0_in_data_ce0;

assign in_data_ce1 = 1'b0;

assign in_data_d0 = 64'd0;

assign in_data_d1 = 64'd0;

assign in_data_read = dataflow_in_loop_TOP_LOOP37928_U0_in_data_write;

assign in_data_we0 = 1'b0;

assign in_data_we1 = 1'b0;

assign out_data_address0 = 14'd0;

assign out_data_address1 = dataflow_in_loop_TOP_LOOP37928_U0_out_data_address1;

assign out_data_ce0 = 1'b0;

assign out_data_ce1 = dataflow_in_loop_TOP_LOOP37928_U0_out_data_ce1;

assign out_data_d0 = 64'd0;

assign out_data_d1 = dataflow_in_loop_TOP_LOOP37928_U0_out_data_d1;

assign out_data_we0 = 1'b0;

assign out_data_we1 = dataflow_in_loop_TOP_LOOP37928_U0_out_data_we1;

assign out_data_write = dataflow_in_loop_TOP_LOOP37928_U0_out_data_write;

endmodule //td_fused_top_tdf3_112
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf3_accum_1 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        accum_in_0_address0,
        accum_in_0_ce0,
        accum_in_0_q0,
        accum_in_0_address1,
        accum_in_0_ce1,
        accum_in_0_q1,
        accum_out_address0,
        accum_out_ce0,
        accum_out_we0,
        accum_out_d0,
        accum_out_address1,
        accum_out_ce1,
        accum_out_we1,
        accum_out_d1
);

parameter    ap_ST_fsm_state1 = 8'd1;
parameter    ap_ST_fsm_pp0_stage0 = 8'd2;
parameter    ap_ST_fsm_pp0_stage1 = 8'd4;
parameter    ap_ST_fsm_pp0_stage2 = 8'd8;
parameter    ap_ST_fsm_pp0_stage3 = 8'd16;
parameter    ap_ST_fsm_state11 = 8'd32;
parameter    ap_ST_fsm_state12 = 8'd64;
parameter    ap_ST_fsm_state13 = 8'd128;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [4:0] accum_in_0_address0;
output   accum_in_0_ce0;
input  [15:0] accum_in_0_q0;
output  [4:0] accum_in_0_address1;
output   accum_in_0_ce1;
input  [15:0] accum_in_0_q1;
output  [2:0] accum_out_address0;
output   accum_out_ce0;
output   accum_out_we0;
output  [15:0] accum_out_d0;
output  [2:0] accum_out_address1;
output   accum_out_ce1;
output   accum_out_we1;
output  [15:0] accum_out_d1;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg[4:0] accum_in_0_address0;
reg accum_in_0_ce0;
reg[4:0] accum_in_0_address1;
reg accum_in_0_ce1;
reg accum_out_ce0;
reg accum_out_we0;
reg accum_out_ce1;
reg accum_out_we1;

reg    ap_done_reg;
  reg   [7:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg   [5:0] x_reg_168;
reg   [15:0] psum_7_08_reg_180;
reg   [15:0] psum_6_07_reg_192;
reg   [15:0] psum_5_06_reg_204;
reg   [15:0] psum_4_05_reg_216;
reg   [15:0] psum_3_04_reg_228;
reg   [15:0] psum_2_03_reg_240;
reg   [15:0] psum_1_02_reg_252;
reg   [15:0] psum_0_01_reg_264;
wire   [0:0] tmp_fu_323_p3;
reg   [0:0] tmp_reg_494;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state6_pp0_stage0_iter1;
wire    ap_block_state10_pp0_stage0_iter2;
wire    ap_block_pp0_stage0_11001;
reg   [0:0] tmp_reg_494_pp0_iter1_reg;
wire   [4:0] trunc_ln25_fu_336_p1;
reg   [4:0] trunc_ln25_reg_498;
wire    ap_CS_fsm_pp0_stage1;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_state3_pp0_stage1_iter0;
wire    ap_block_state7_pp0_stage1_iter1;
wire    ap_block_pp0_stage1_11001;
wire    ap_CS_fsm_pp0_stage2;
wire    ap_block_state4_pp0_stage2_iter0;
wire    ap_block_state8_pp0_stage2_iter1;
wire    ap_block_pp0_stage2_11001;
wire   [5:0] add_ln25_fu_391_p2;
reg   [5:0] add_ln25_reg_558;
wire    ap_CS_fsm_pp0_stage3;
wire    ap_block_state5_pp0_stage3_iter0;
wire    ap_block_state9_pp0_stage3_iter1;
wire    ap_block_pp0_stage3_11001;
reg    ap_enable_reg_pp0_iter1;
wire   [15:0] grp_fu_305_p2;
wire   [15:0] grp_fu_311_p2;
reg    ap_enable_reg_pp0_iter2;
wire   [3:0] add_ln33_fu_434_p2;
wire    ap_CS_fsm_state12;
wire   [0:0] tmp_36_fu_417_p3;
reg    ap_block_state1;
wire    ap_block_pp0_stage1_subdone;
reg    ap_condition_pp0_exit_iter0_state3;
wire    ap_block_pp0_stage3_subdone;
wire    ap_block_pp0_stage0_subdone;
reg   [5:0] ap_phi_mux_x_phi_fu_172_p4;
wire    ap_block_pp0_stage0;
wire   [15:0] ap_phi_mux_psum_7_08_phi_fu_184_p4;
wire   [15:0] ap_phi_mux_psum_6_07_phi_fu_196_p4;
wire   [15:0] ap_phi_mux_psum_5_06_phi_fu_208_p4;
wire    ap_block_pp0_stage3;
wire   [15:0] ap_phi_mux_psum_4_05_phi_fu_220_p4;
wire   [15:0] ap_phi_mux_psum_3_04_phi_fu_232_p4;
wire    ap_block_pp0_stage2;
wire   [15:0] ap_phi_mux_psum_2_03_phi_fu_244_p4;
wire    ap_block_pp0_stage1;
reg   [3:0] q_reg_276;
wire    ap_CS_fsm_state11;
reg   [15:0] ap_phi_mux_phi_ln45_phi_fu_290_p8;
wire   [2:0] trunc_ln33_fu_430_p1;
wire   [63:0] zext_ln25_fu_331_p1;
wire   [63:0] zext_ln29_fu_346_p1;
wire   [63:0] zext_ln29_13_fu_356_p1;
wire   [63:0] zext_ln29_14_fu_366_p1;
wire   [63:0] zext_ln29_15_fu_376_p1;
wire   [63:0] zext_ln29_16_fu_386_p1;
wire   [63:0] zext_ln29_17_fu_402_p1;
wire   [63:0] zext_ln29_18_fu_412_p1;
wire   [63:0] zext_ln33_fu_425_p1;
wire   [63:0] zext_ln33_3_fu_446_p1;
reg   [15:0] grp_fu_305_p0;
reg   [15:0] grp_fu_311_p0;
wire   [4:0] or_ln29_fu_340_p2;
wire   [4:0] or_ln29_13_fu_351_p2;
wire   [4:0] or_ln29_14_fu_361_p2;
wire   [4:0] or_ln29_15_fu_371_p2;
wire   [4:0] or_ln29_16_fu_381_p2;
wire   [4:0] or_ln29_17_fu_397_p2;
wire   [4:0] or_ln29_18_fu_407_p2;
wire   [2:0] or_ln33_fu_440_p2;
wire   [0:0] icmp_ln45_fu_451_p2;
wire   [0:0] icmp_ln45_5_fu_465_p2;
wire   [15:0] select_ln45_fu_457_p3;
wire   [0:0] icmp_ln45_6_fu_479_p2;
wire   [15:0] select_ln45_5_fu_471_p3;
wire    ap_CS_fsm_state13;
reg   [7:0] ap_NS_fsm;
wire    ap_block_pp0_stage2_subdone;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
reg    ap_condition_499;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 8'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
end

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U162(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(grp_fu_305_p0),
    .din1(accum_in_0_q1),
    .dout(grp_fu_305_p2)
);

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U163(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(grp_fu_311_p0),
    .din1(accum_in_0_q0),
    .dout(grp_fu_311_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state13)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b1 == ap_condition_pp0_exit_iter0_state3))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage3_subdone) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b0)) | ((1'b0 == ap_block_pp0_stage3_subdone) & (1'b1 == ap_CS_fsm_pp0_stage3)))) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end else if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter2 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state11)) begin
        q_reg_276 <= 4'd0;
    end else if (((tmp_36_fu_417_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state12))) begin
        q_reg_276 <= add_ln33_fu_434_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (tmp_reg_494 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        x_reg_168 <= add_ln25_reg_558;
    end else if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        x_reg_168 <= 6'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage3_11001) & (tmp_reg_494 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage3) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
        add_ln25_reg_558 <= add_ln25_fu_391_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((tmp_reg_494_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        psum_0_01_reg_264 <= grp_fu_305_p2;
        psum_1_02_reg_252 <= grp_fu_311_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((tmp_reg_494_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage2_11001) & (1'b1 == ap_CS_fsm_pp0_stage2) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        psum_2_03_reg_240 <= grp_fu_305_p2;
        psum_3_04_reg_228 <= grp_fu_311_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((tmp_reg_494_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage3_11001) & (1'b1 == ap_CS_fsm_pp0_stage3) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        psum_4_05_reg_216 <= grp_fu_305_p2;
        psum_5_06_reg_204 <= grp_fu_311_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((tmp_reg_494_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        psum_6_07_reg_192 <= grp_fu_305_p2;
        psum_7_08_reg_180 <= grp_fu_311_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_reg_494 <= ap_phi_mux_x_phi_fu_172_p4[32'd5];
        tmp_reg_494_pp0_iter1_reg <= tmp_reg_494;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (tmp_fu_323_p3 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        trunc_ln25_reg_498 <= trunc_ln25_fu_336_p1;
    end
end

always @ (*) begin
    if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
        if (((1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            accum_in_0_address0 = zext_ln29_18_fu_412_p1;
        end else if (((1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            accum_in_0_address0 = zext_ln29_16_fu_386_p1;
        end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            accum_in_0_address0 = zext_ln29_14_fu_366_p1;
        end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            accum_in_0_address0 = zext_ln29_fu_346_p1;
        end else begin
            accum_in_0_address0 = 'bx;
        end
    end else begin
        accum_in_0_address0 = 'bx;
    end
end

always @ (*) begin
    if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
        if (((1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            accum_in_0_address1 = zext_ln29_17_fu_402_p1;
        end else if (((1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            accum_in_0_address1 = zext_ln29_15_fu_376_p1;
        end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            accum_in_0_address1 = zext_ln29_13_fu_356_p1;
        end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            accum_in_0_address1 = zext_ln25_fu_331_p1;
        end else begin
            accum_in_0_address1 = 'bx;
        end
    end else begin
        accum_in_0_address1 = 'bx;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1)) | ((1'b0 == ap_block_pp0_stage3_11001) & (1'b1 == ap_CS_fsm_pp0_stage3) & (ap_enable_reg_pp0_iter0 == 1'b1)) | ((1'b0 == ap_block_pp0_stage2_11001) & (1'b1 == ap_CS_fsm_pp0_stage2) & (ap_enable_reg_pp0_iter0 == 1'b1)) | ((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1)))) begin
        accum_in_0_ce0 = 1'b1;
    end else begin
        accum_in_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1)) | ((1'b0 == ap_block_pp0_stage3_11001) & (1'b1 == ap_CS_fsm_pp0_stage3) & (ap_enable_reg_pp0_iter0 == 1'b1)) | ((1'b0 == ap_block_pp0_stage2_11001) & (1'b1 == ap_CS_fsm_pp0_stage2) & (ap_enable_reg_pp0_iter0 == 1'b1)) | ((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1)))) begin
        accum_in_0_ce1 = 1'b1;
    end else begin
        accum_in_0_ce1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state12)) begin
        accum_out_ce0 = 1'b1;
    end else begin
        accum_out_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state12)) begin
        accum_out_ce1 = 1'b1;
    end else begin
        accum_out_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((tmp_36_fu_417_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state12))) begin
        accum_out_we0 = 1'b1;
    end else begin
        accum_out_we0 = 1'b0;
    end
end

always @ (*) begin
    if (((tmp_36_fu_417_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state12))) begin
        accum_out_we1 = 1'b1;
    end else begin
        accum_out_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((tmp_reg_494 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state3 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state3 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state13)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((tmp_36_fu_417_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state12))) begin
        if ((trunc_ln33_fu_430_p1 == 3'd0)) begin
            ap_phi_mux_phi_ln45_phi_fu_290_p8 = psum_0_01_reg_264;
        end else if ((1'b1 == ap_condition_499)) begin
            ap_phi_mux_phi_ln45_phi_fu_290_p8 = psum_6_07_reg_192;
        end else if ((trunc_ln33_fu_430_p1 == 3'd4)) begin
            ap_phi_mux_phi_ln45_phi_fu_290_p8 = psum_4_05_reg_216;
        end else if ((trunc_ln33_fu_430_p1 == 3'd2)) begin
            ap_phi_mux_phi_ln45_phi_fu_290_p8 = psum_2_03_reg_240;
        end else begin
            ap_phi_mux_phi_ln45_phi_fu_290_p8 = 'bx;
        end
    end else begin
        ap_phi_mux_phi_ln45_phi_fu_290_p8 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0) & (tmp_reg_494 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_x_phi_fu_172_p4 = add_ln25_reg_558;
    end else begin
        ap_phi_mux_x_phi_fu_172_p4 = x_reg_168;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state13)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_305_p0 = ap_phi_mux_psum_6_07_phi_fu_196_p4;
    end else if (((1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
        grp_fu_305_p0 = ap_phi_mux_psum_4_05_phi_fu_220_p4;
    end else if (((1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
        grp_fu_305_p0 = ap_phi_mux_psum_2_03_phi_fu_244_p4;
    end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
        grp_fu_305_p0 = grp_fu_305_p2;
    end else begin
        grp_fu_305_p0 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_311_p0 = ap_phi_mux_psum_7_08_phi_fu_184_p4;
    end else if (((1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
        grp_fu_311_p0 = ap_phi_mux_psum_5_06_phi_fu_208_p4;
    end else if (((1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
        grp_fu_311_p0 = ap_phi_mux_psum_3_04_phi_fu_232_p4;
    end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
        grp_fu_311_p0 = grp_fu_311_p2;
    end else begin
        grp_fu_311_p0 = 'bx;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((~((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0)) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end else if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
                ap_NS_fsm = ap_ST_fsm_state11;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_pp0_stage1 : begin
            if ((~((1'b0 == ap_block_pp0_stage1_subdone) & (tmp_reg_494 == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1)) & (1'b0 == ap_block_pp0_stage1_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage2;
            end else if (((1'b0 == ap_block_pp0_stage1_subdone) & (tmp_reg_494 == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
                ap_NS_fsm = ap_ST_fsm_state11;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end
        end
        ap_ST_fsm_pp0_stage2 : begin
            if ((1'b0 == ap_block_pp0_stage2_subdone)) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage3;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage2;
            end
        end
        ap_ST_fsm_pp0_stage3 : begin
            if ((1'b0 == ap_block_pp0_stage3_subdone)) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage3;
            end
        end
        ap_ST_fsm_state11 : begin
            ap_NS_fsm = ap_ST_fsm_state12;
        end
        ap_ST_fsm_state12 : begin
            if (((tmp_36_fu_417_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state12))) begin
                ap_NS_fsm = ap_ST_fsm_state12;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state13;
            end
        end
        ap_ST_fsm_state13 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign accum_out_address0 = zext_ln33_3_fu_446_p1;

assign accum_out_address1 = zext_ln33_fu_425_p1;

assign accum_out_d0 = ((icmp_ln45_6_fu_479_p2[0:0] == 1'b1) ? psum_5_06_reg_204 : select_ln45_5_fu_471_p3);

assign accum_out_d1 = ap_phi_mux_phi_ln45_phi_fu_290_p8;

assign add_ln25_fu_391_p2 = (x_reg_168 + 6'd8);

assign add_ln33_fu_434_p2 = (q_reg_276 + 4'd2);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_pp0_stage1 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_pp0_stage2 = ap_CS_fsm[32'd3];

assign ap_CS_fsm_pp0_stage3 = ap_CS_fsm[32'd4];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state11 = ap_CS_fsm[32'd5];

assign ap_CS_fsm_state12 = ap_CS_fsm[32'd6];

assign ap_CS_fsm_state13 = ap_CS_fsm[32'd7];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1_subdone = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage2 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage2_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage2_subdone = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage3 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage3_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage3_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((ap_done_reg == 1'b1) | (ap_start == 1'b0));
end

assign ap_block_state10_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage1_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage2_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage3_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage1_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage2_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state9_pp0_stage3_iter1 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_condition_499 = (~(trunc_ln33_fu_430_p1 == 3'd0) & ~(trunc_ln33_fu_430_p1 == 3'd4) & ~(trunc_ln33_fu_430_p1 == 3'd2));
end

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign ap_phi_mux_psum_2_03_phi_fu_244_p4 = grp_fu_305_p2;

assign ap_phi_mux_psum_3_04_phi_fu_232_p4 = grp_fu_311_p2;

assign ap_phi_mux_psum_4_05_phi_fu_220_p4 = grp_fu_305_p2;

assign ap_phi_mux_psum_5_06_phi_fu_208_p4 = grp_fu_311_p2;

assign ap_phi_mux_psum_6_07_phi_fu_196_p4 = grp_fu_305_p2;

assign ap_phi_mux_psum_7_08_phi_fu_184_p4 = grp_fu_311_p2;

assign icmp_ln45_5_fu_465_p2 = ((or_ln33_fu_440_p2 == 3'd3) ? 1'b1 : 1'b0);

assign icmp_ln45_6_fu_479_p2 = ((or_ln33_fu_440_p2 == 3'd5) ? 1'b1 : 1'b0);

assign icmp_ln45_fu_451_p2 = ((or_ln33_fu_440_p2 == 3'd1) ? 1'b1 : 1'b0);

assign or_ln29_13_fu_351_p2 = (trunc_ln25_reg_498 | 5'd2);

assign or_ln29_14_fu_361_p2 = (trunc_ln25_reg_498 | 5'd3);

assign or_ln29_15_fu_371_p2 = (trunc_ln25_reg_498 | 5'd4);

assign or_ln29_16_fu_381_p2 = (trunc_ln25_reg_498 | 5'd5);

assign or_ln29_17_fu_397_p2 = (trunc_ln25_reg_498 | 5'd6);

assign or_ln29_18_fu_407_p2 = (trunc_ln25_reg_498 | 5'd7);

assign or_ln29_fu_340_p2 = (trunc_ln25_fu_336_p1 | 5'd1);

assign or_ln33_fu_440_p2 = (trunc_ln33_fu_430_p1 | 3'd1);

assign select_ln45_5_fu_471_p3 = ((icmp_ln45_5_fu_465_p2[0:0] == 1'b1) ? psum_3_04_reg_228 : select_ln45_fu_457_p3);

assign select_ln45_fu_457_p3 = ((icmp_ln45_fu_451_p2[0:0] == 1'b1) ? psum_1_02_reg_252 : psum_7_08_reg_180);

assign tmp_36_fu_417_p3 = q_reg_276[32'd3];

assign tmp_fu_323_p3 = ap_phi_mux_x_phi_fu_172_p4[32'd5];

assign trunc_ln25_fu_336_p1 = ap_phi_mux_x_phi_fu_172_p4[4:0];

assign trunc_ln33_fu_430_p1 = q_reg_276[2:0];

assign zext_ln25_fu_331_p1 = ap_phi_mux_x_phi_fu_172_p4;

assign zext_ln29_13_fu_356_p1 = or_ln29_13_fu_351_p2;

assign zext_ln29_14_fu_366_p1 = or_ln29_14_fu_361_p2;

assign zext_ln29_15_fu_376_p1 = or_ln29_15_fu_371_p2;

assign zext_ln29_16_fu_386_p1 = or_ln29_16_fu_381_p2;

assign zext_ln29_17_fu_402_p1 = or_ln29_17_fu_397_p2;

assign zext_ln29_18_fu_412_p1 = or_ln29_18_fu_407_p2;

assign zext_ln29_fu_346_p1 = or_ln29_fu_340_p2;

assign zext_ln33_3_fu_446_p1 = or_ln33_fu_440_p2;

assign zext_ln33_fu_425_p1 = q_reg_276;

endmodule //td_fused_top_tdf3_accum_1
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf3_accum_2 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        accum_in_14,
        accum_in_14_ap_vld,
        accum_in_address0,
        accum_in_ce0,
        accum_in_q0
);

parameter    ap_ST_fsm_state1 = 7'd1;
parameter    ap_ST_fsm_state2 = 7'd2;
parameter    ap_ST_fsm_state3 = 7'd4;
parameter    ap_ST_fsm_state4 = 7'd8;
parameter    ap_ST_fsm_state5 = 7'd16;
parameter    ap_ST_fsm_state6 = 7'd32;
parameter    ap_ST_fsm_state7 = 7'd64;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [15:0] accum_in_14;
output   accum_in_14_ap_vld;
output  [2:0] accum_in_address0;
output   accum_in_ce0;
input  [15:0] accum_in_q0;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg[15:0] accum_in_14;
reg accum_in_14_ap_vld;
reg accum_in_ce0;

reg    ap_done_reg;
  reg   [6:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
wire   [3:0] add_ln57_fu_74_p2;
reg   [3:0] add_ln57_reg_91;
wire    ap_CS_fsm_state2;
wire   [0:0] icmp_ln57_fu_85_p2;
wire    ap_CS_fsm_state3;
wire   [15:0] grp_fu_68_p2;
wire    ap_CS_fsm_state7;
reg   [3:0] i_1_1_reg_44;
reg    ap_block_state1;
reg   [15:0] sum_01_reg_55;
wire   [63:0] zext_ln57_fu_80_p1;
reg   [15:0] accum_in_14_preg;
reg   [6:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 7'd1;
#0 accum_in_14_preg = 16'd0;
end

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U166(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(sum_01_reg_55),
    .din1(accum_in_q0),
    .dout(grp_fu_68_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        accum_in_14_preg <= 16'd0;
    end else begin
        if (((icmp_ln57_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
            accum_in_14_preg <= sum_01_reg_55;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if (((icmp_ln57_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        i_1_1_reg_44 <= 4'd0;
    end else if ((1'b1 == ap_CS_fsm_state7)) begin
        i_1_1_reg_44 <= add_ln57_reg_91;
    end
end

always @ (posedge ap_clk) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        sum_01_reg_55 <= 16'd0;
    end else if ((1'b1 == ap_CS_fsm_state7)) begin
        sum_01_reg_55 <= grp_fu_68_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        add_ln57_reg_91 <= add_ln57_fu_74_p2;
    end
end

always @ (*) begin
    if (((icmp_ln57_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        accum_in_14 = sum_01_reg_55;
    end else begin
        accum_in_14 = accum_in_14_preg;
    end
end

always @ (*) begin
    if (((icmp_ln57_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        accum_in_14_ap_vld = 1'b1;
    end else begin
        accum_in_14_ap_vld = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        accum_in_ce0 = 1'b1;
    end else begin
        accum_in_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln57_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln57_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_state2 : begin
            if (((icmp_ln57_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end
        end
        ap_ST_fsm_state3 : begin
            ap_NS_fsm = ap_ST_fsm_state4;
        end
        ap_ST_fsm_state4 : begin
            ap_NS_fsm = ap_ST_fsm_state5;
        end
        ap_ST_fsm_state5 : begin
            ap_NS_fsm = ap_ST_fsm_state6;
        end
        ap_ST_fsm_state6 : begin
            ap_NS_fsm = ap_ST_fsm_state7;
        end
        ap_ST_fsm_state7 : begin
            ap_NS_fsm = ap_ST_fsm_state2;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign accum_in_address0 = zext_ln57_fu_80_p1;

assign add_ln57_fu_74_p2 = (i_1_1_reg_44 + 4'd1);

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state7 = ap_CS_fsm[32'd6];

always @ (*) begin
    ap_block_state1 = ((ap_done_reg == 1'b1) | (ap_start == 1'b0));
end

assign icmp_ln57_fu_85_p2 = ((i_1_1_reg_44 == 4'd8) ? 1'b1 : 1'b0);

assign zext_ln57_fu_80_p1 = i_1_1_reg_44;

endmodule //td_fused_top_tdf3_accum_2
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf3_adjust (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        sums_read,
        adjustments_address0,
        adjustments_ce0,
        adjustments_q0,
        indices_23_dout,
        indices_23_empty_n,
        indices_23_read,
        ap_return
);

parameter    ap_ST_fsm_state1 = 17'd1;
parameter    ap_ST_fsm_state2 = 17'd2;
parameter    ap_ST_fsm_state3 = 17'd4;
parameter    ap_ST_fsm_state4 = 17'd8;
parameter    ap_ST_fsm_state5 = 17'd16;
parameter    ap_ST_fsm_state6 = 17'd32;
parameter    ap_ST_fsm_state7 = 17'd64;
parameter    ap_ST_fsm_state8 = 17'd128;
parameter    ap_ST_fsm_state9 = 17'd256;
parameter    ap_ST_fsm_state10 = 17'd512;
parameter    ap_ST_fsm_state11 = 17'd1024;
parameter    ap_ST_fsm_state12 = 17'd2048;
parameter    ap_ST_fsm_state13 = 17'd4096;
parameter    ap_ST_fsm_state14 = 17'd8192;
parameter    ap_ST_fsm_state15 = 17'd16384;
parameter    ap_ST_fsm_state16 = 17'd32768;
parameter    ap_ST_fsm_state17 = 17'd65536;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
input  [15:0] sums_read;
output  [3:0] adjustments_address0;
output   adjustments_ce0;
input  [47:0] adjustments_q0;
input  [3:0] indices_23_dout;
input   indices_23_empty_n;
output   indices_23_read;
output  [15:0] ap_return;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg adjustments_ce0;
reg indices_23_read;

reg    ap_done_reg;
  reg   [16:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    indices_23_blk_n;
wire    ap_CS_fsm_state4;
reg   [15:0] tmp_61_i_i_reg_167;
reg   [15:0] tmp_62_i_i_reg_172;
wire   [15:0] grp_fu_81_p2;
reg   [15:0] sub_i_i_i_reg_177;
wire    ap_CS_fsm_state8;
wire    ap_CS_fsm_state9;
wire   [15:0] grp_fu_86_p2;
reg   [15:0] mul_i_i_i_reg_187;
wire    ap_CS_fsm_state12;
wire    ap_CS_fsm_state13;
wire   [63:0] zext_ln220_fu_90_p1;
reg    ap_block_state1;
wire    ap_CS_fsm_state2;
wire    ap_CS_fsm_state3;
wire   [15:0] grp_fu_77_p1;
wire   [15:0] grp_fu_81_p1;
wire   [15:0] grp_fu_86_p1;
wire   [15:0] trunc_ln220_fu_95_p1;
wire   [15:0] grp_fu_77_p2;
wire    ap_CS_fsm_state17;
wire   [15:0] bitcast_ln648_fu_132_p1;
wire   [0:0] tmp_fu_136_p3;
reg   [16:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 17'd1;
end

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U170(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(mul_i_i_i_reg_187),
    .din1(grp_fu_77_p1),
    .dout(grp_fu_77_p2)
);

td_fused_top_hsub_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hsub_16ns_16ns_16_5_full_dsp_1_U171(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(sums_read),
    .din1(grp_fu_81_p1),
    .dout(grp_fu_81_p2)
);

td_fused_top_hmul_16ns_16ns_16_4_max_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hmul_16ns_16ns_16_4_max_dsp_1_U172(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(sub_i_i_i_reg_177),
    .din1(grp_fu_86_p1),
    .dout(grp_fu_86_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state17)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state12)) begin
        mul_i_i_i_reg_187 <= grp_fu_86_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state8)) begin
        sub_i_i_i_reg_177 <= grp_fu_81_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        tmp_61_i_i_reg_167 <= {{adjustments_q0[31:16]}};
        tmp_62_i_i_reg_172 <= {{adjustments_q0[47:32]}};
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state2) | (~((indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1)))) begin
        adjustments_ce0 = 1'b1;
    end else begin
        adjustments_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state17)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state17)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_23_blk_n = indices_23_empty_n;
    end else begin
        indices_23_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_23_read = 1'b1;
    end else begin
        indices_23_read = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_state2 : begin
            ap_NS_fsm = ap_ST_fsm_state3;
        end
        ap_ST_fsm_state3 : begin
            ap_NS_fsm = ap_ST_fsm_state4;
        end
        ap_ST_fsm_state4 : begin
            ap_NS_fsm = ap_ST_fsm_state5;
        end
        ap_ST_fsm_state5 : begin
            ap_NS_fsm = ap_ST_fsm_state6;
        end
        ap_ST_fsm_state6 : begin
            ap_NS_fsm = ap_ST_fsm_state7;
        end
        ap_ST_fsm_state7 : begin
            ap_NS_fsm = ap_ST_fsm_state8;
        end
        ap_ST_fsm_state8 : begin
            ap_NS_fsm = ap_ST_fsm_state9;
        end
        ap_ST_fsm_state9 : begin
            ap_NS_fsm = ap_ST_fsm_state10;
        end
        ap_ST_fsm_state10 : begin
            ap_NS_fsm = ap_ST_fsm_state11;
        end
        ap_ST_fsm_state11 : begin
            ap_NS_fsm = ap_ST_fsm_state12;
        end
        ap_ST_fsm_state12 : begin
            ap_NS_fsm = ap_ST_fsm_state13;
        end
        ap_ST_fsm_state13 : begin
            ap_NS_fsm = ap_ST_fsm_state14;
        end
        ap_ST_fsm_state14 : begin
            ap_NS_fsm = ap_ST_fsm_state15;
        end
        ap_ST_fsm_state15 : begin
            ap_NS_fsm = ap_ST_fsm_state16;
        end
        ap_ST_fsm_state16 : begin
            ap_NS_fsm = ap_ST_fsm_state17;
        end
        ap_ST_fsm_state17 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign adjustments_address0 = zext_ln220_fu_90_p1;

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state12 = ap_CS_fsm[32'd11];

assign ap_CS_fsm_state13 = ap_CS_fsm[32'd12];

assign ap_CS_fsm_state17 = ap_CS_fsm[32'd16];

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

assign ap_CS_fsm_state8 = ap_CS_fsm[32'd7];

assign ap_CS_fsm_state9 = ap_CS_fsm[32'd8];

always @ (*) begin
    ap_block_state1 = ((indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0));
end

assign ap_return = ((tmp_fu_136_p3[0:0] == 1'b1) ? 16'd0 : grp_fu_77_p2);

assign bitcast_ln648_fu_132_p1 = grp_fu_77_p2;

assign grp_fu_77_p1 = tmp_62_i_i_reg_172;

assign grp_fu_81_p1 = trunc_ln220_fu_95_p1;

assign grp_fu_86_p1 = tmp_61_i_i_reg_167;

assign tmp_fu_136_p3 = bitcast_ln648_fu_132_p1[32'd15];

assign trunc_ln220_fu_95_p1 = adjustments_q0[15:0];

assign zext_ln220_fu_90_p1 = indices_23_dout;

endmodule //td_fused_top_tdf3_adjust
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf3_dot_product (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        ifmap_vec_0_0_address0,
        ifmap_vec_0_0_ce0,
        ifmap_vec_0_0_q0,
        weight_vecs_0_0_0_address0,
        weight_vecs_0_0_0_ce0,
        weight_vecs_0_0_0_q0,
        products_0_address0,
        products_0_ce0,
        products_0_we0,
        products_0_d0
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state7 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [4:0] ifmap_vec_0_0_address0;
output   ifmap_vec_0_0_ce0;
input  [15:0] ifmap_vec_0_0_q0;
output  [4:0] weight_vecs_0_0_0_address0;
output   weight_vecs_0_0_0_ce0;
input  [15:0] weight_vecs_0_0_0_q0;
output  [4:0] products_0_address0;
output   products_0_ce0;
output   products_0_we0;
output  [15:0] products_0_d0;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg ifmap_vec_0_0_ce0;
reg weight_vecs_0_0_0_ce0;
reg products_0_ce0;
reg products_0_we0;

reg    ap_done_reg;
  reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg   [5:0] ic_0_0_reg_69;
wire   [5:0] add_ln149_fu_87_p2;
wire    ap_CS_fsm_pp0_stage0;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
wire    ap_block_state4_pp0_stage0_iter2;
wire    ap_block_state5_pp0_stage0_iter3;
wire    ap_block_state6_pp0_stage0_iter4;
wire    ap_block_pp0_stage0_11001;
wire   [0:0] icmp_ln149_fu_93_p2;
reg   [0:0] icmp_ln149_reg_118;
reg   [0:0] icmp_ln149_reg_118_pp0_iter1_reg;
reg   [0:0] icmp_ln149_reg_118_pp0_iter2_reg;
reg   [0:0] icmp_ln149_reg_118_pp0_iter3_reg;
wire   [4:0] trunc_ln150_fu_105_p1;
reg   [4:0] trunc_ln150_reg_122;
reg   [4:0] trunc_ln150_reg_122_pp0_iter1_reg;
reg   [4:0] trunc_ln150_reg_122_pp0_iter2_reg;
reg   [4:0] trunc_ln150_reg_122_pp0_iter3_reg;
reg    ap_block_state1;
wire    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_exit_iter0_state2;
reg    ap_enable_reg_pp0_iter1;
reg    ap_enable_reg_pp0_iter2;
reg    ap_enable_reg_pp0_iter3;
reg    ap_enable_reg_pp0_iter4;
wire   [63:0] zext_ln149_fu_99_p1;
wire    ap_block_pp0_stage0;
wire   [63:0] idxprom30_0_0_fu_109_p1;
wire   [15:0] grp_fu_80_p2;
wire    ap_CS_fsm_state7;
reg   [2:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
#0 ap_enable_reg_pp0_iter4 = 1'b0;
end

td_fused_top_hmul_16ns_16ns_16_4_max_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hmul_16ns_16ns_16_4_max_dsp_1_U158(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(ifmap_vec_0_0_q0),
    .din1(weight_vecs_0_0_0_q0),
    .dout(grp_fu_80_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state7)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b1 == ap_condition_pp0_exit_iter0_state2))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            if ((1'b1 == ap_condition_pp0_exit_iter0_state2)) begin
                ap_enable_reg_pp0_iter1 <= (1'b1 ^ ap_condition_pp0_exit_iter0_state2);
            end else if ((1'b1 == 1'b1)) begin
                ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
            end
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter4 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
        end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter4 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ic_0_0_reg_69 <= 6'd0;
    end else if (((icmp_ln149_fu_93_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ic_0_0_reg_69 <= add_ln149_fu_87_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln149_reg_118 <= icmp_ln149_fu_93_p2;
        icmp_ln149_reg_118_pp0_iter1_reg <= icmp_ln149_reg_118;
        trunc_ln150_reg_122_pp0_iter1_reg <= trunc_ln150_reg_122;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        icmp_ln149_reg_118_pp0_iter2_reg <= icmp_ln149_reg_118_pp0_iter1_reg;
        icmp_ln149_reg_118_pp0_iter3_reg <= icmp_ln149_reg_118_pp0_iter2_reg;
        trunc_ln150_reg_122_pp0_iter2_reg <= trunc_ln150_reg_122_pp0_iter1_reg;
        trunc_ln150_reg_122_pp0_iter3_reg <= trunc_ln150_reg_122_pp0_iter2_reg;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln149_fu_93_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        trunc_ln150_reg_122 <= trunc_ln150_fu_105_p1;
    end
end

always @ (*) begin
    if ((icmp_ln149_fu_93_p2 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state2 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state2 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state7)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state7)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ifmap_vec_0_0_ce0 = 1'b1;
    end else begin
        ifmap_vec_0_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter4 == 1'b1))) begin
        products_0_ce0 = 1'b1;
    end else begin
        products_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln149_reg_118_pp0_iter3_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter4 == 1'b1))) begin
        products_0_we0 = 1'b1;
    end else begin
        products_0_we0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        weight_vecs_0_0_0_ce0 = 1'b1;
    end else begin
        weight_vecs_0_0_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((~((icmp_ln149_fu_93_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0)) & ~((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter4 == 1'b1) & (ap_enable_reg_pp0_iter3 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if ((((icmp_ln149_fu_93_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0)) | ((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter4 == 1'b1) & (ap_enable_reg_pp0_iter3 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_state7;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state7 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln149_fu_87_p2 = (ic_0_0_reg_69 + 6'd1);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state7 = ap_CS_fsm[32'd2];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (ap_done_reg == 1'b1));
end

assign ap_block_state2_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter4 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign icmp_ln149_fu_93_p2 = ((ic_0_0_reg_69 == 6'd32) ? 1'b1 : 1'b0);

assign idxprom30_0_0_fu_109_p1 = trunc_ln150_reg_122_pp0_iter3_reg;

assign ifmap_vec_0_0_address0 = zext_ln149_fu_99_p1;

assign products_0_address0 = idxprom30_0_0_fu_109_p1;

assign products_0_d0 = grp_fu_80_p2;

assign trunc_ln150_fu_105_p1 = ic_0_0_reg_69[4:0];

assign weight_vecs_0_0_0_address0 = zext_ln149_fu_99_p1;

assign zext_ln149_fu_99_p1 = ic_0_0_reg_69;

endmodule //td_fused_top_tdf3_dot_product
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_tdf3_filters_ram (addr0, ce0, q0, addr1, ce1, d1, we1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 9;
parameter MEM_SIZE = 512;

input[AWIDTH-1:0] addr0;
input ce0;
output wire[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
input clk;

 reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];
wire [AWIDTH-1:0] addr0_t0; 
reg [AWIDTH-1:0] addr0_t1; 
reg [DWIDTH-1:0] q0_t0;
reg [DWIDTH-1:0] q0_t1;
wire [AWIDTH-1:0] addr1_t0; 
reg [AWIDTH-1:0] addr1_t1; 
wire [DWIDTH-1:0] d1_t0; 
wire we1_t0; 
reg [DWIDTH-1:0] d1_t1; 
reg we1_t1; 


assign addr0_t0 = addr0;
assign q0 = q0_t1;
assign addr1_t0 = addr1;
assign d1_t0 = d1;
assign we1_t0 = we1;

always @(posedge clk)  
begin
    if (ce0) 
    begin
        addr0_t1 <= addr0_t0; 
        q0_t1 <= q0_t0;
    end
    if (ce1) 
    begin
        addr1_t1 <= addr1_t0; 
        d1_t1 <= d1_t0;
        we1_t1 <= we1_t0;
    end
end


always @(posedge clk)  
begin 
    if (ce0) begin
        q0_t0 <= ram[addr0_t1];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1_t1) 
            ram[addr1_t1] <= d1_t1; 
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_tdf3_filters(
    reset,
    clk,
    address0,
    ce0,
    q0,
    address1,
    ce1,
    we1,
    d1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd512;
parameter AddressWidth = 32'd9;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;



td_fused_top_tdf3_filters_ram td_fused_top_tdf3_filters_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 )
);

endmodule

// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf3_get_next_ijk (
        ap_clk,
        ap_rst,
        ap_start,
        start_full_n,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        start_out,
        start_write,
        indices_0_din,
        indices_0_full_n,
        indices_0_write,
        indices_1_din,
        indices_1_full_n,
        indices_1_write,
        indices_2_out_din,
        indices_2_out_full_n,
        indices_2_out_write,
        indices_2_out1_din,
        indices_2_out1_full_n,
        indices_2_out1_write
);

parameter    ap_ST_fsm_state1 = 1'd1;

input   ap_clk;
input   ap_rst;
input   ap_start;
input   start_full_n;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output   start_out;
output   start_write;
output  [15:0] indices_0_din;
input   indices_0_full_n;
output   indices_0_write;
output  [15:0] indices_1_din;
input   indices_1_full_n;
output   indices_1_write;
output  [3:0] indices_2_out_din;
input   indices_2_out_full_n;
output   indices_2_out_write;
output  [3:0] indices_2_out1_din;
input   indices_2_out1_full_n;
output   indices_2_out1_write;

reg ap_done;
reg ap_idle;
reg start_write;
reg indices_0_write;
reg indices_1_write;
reg indices_2_out_write;
reg indices_2_out1_write;

reg    real_start;
reg    start_once_reg;
reg    ap_done_reg;
  reg   [0:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    internal_ap_ready;
reg   [15:0] i_2;
reg   [15:0] j_2;
reg   [15:0] k_2;
reg    indices_0_blk_n;
reg    indices_1_blk_n;
reg    indices_2_out_blk_n;
reg    indices_2_out1_blk_n;
reg   [0:0] ap_phi_mux_j_14_flag_0_i_phi_fu_77_p6;
reg    ap_block_state1;
wire   [0:0] icmp_ln78_fu_141_p2;
wire   [0:0] icmp_ln81_fu_154_p2;
reg   [15:0] ap_phi_mux_j_14_new_0_i_phi_fu_91_p6;
wire   [15:0] add_ln80_fu_147_p2;
reg   [15:0] ap_phi_mux_k_14_new_0_i_phi_fu_104_p6;
wire   [15:0] add_ln77_fu_134_p2;
wire   [15:0] select_ln84_fu_172_p3;
wire   [3:0] trunc_ln76_fu_128_p1;
wire   [15:0] add_ln83_fu_160_p2;
wire   [0:0] icmp_ln84_fu_166_p2;
reg   [0:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 start_once_reg = 1'b0;
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 1'd1;
#0 i_2 = 16'd0;
#0 j_2 = 16'd0;
#0 k_2 = 16'd0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((~((real_start == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        start_once_reg <= 1'b0;
    end else begin
        if (((real_start == 1'b1) & (internal_ap_ready == 1'b0))) begin
            start_once_reg <= 1'b1;
        end else if ((internal_ap_ready == 1'b1)) begin
            start_once_reg <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((~((real_start == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (icmp_ln81_fu_154_p2 == 1'd1) & (icmp_ln78_fu_141_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1))) begin
        i_2 <= select_ln84_fu_172_p3;
    end
end

always @ (posedge ap_clk) begin
    if ((~((real_start == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (ap_phi_mux_j_14_flag_0_i_phi_fu_77_p6 == 1'd1) & (1'b1 == ap_CS_fsm_state1))) begin
        j_2 <= ap_phi_mux_j_14_new_0_i_phi_fu_91_p6;
    end
end

always @ (posedge ap_clk) begin
    if ((~((real_start == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        k_2 <= ap_phi_mux_k_14_new_0_i_phi_fu_104_p6;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((real_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln78_fu_141_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_phi_mux_j_14_flag_0_i_phi_fu_77_p6 = 1'd0;
    end else if ((((icmp_ln81_fu_154_p2 == 1'd0) & (icmp_ln78_fu_141_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1)) | ((icmp_ln81_fu_154_p2 == 1'd1) & (icmp_ln78_fu_141_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1)))) begin
        ap_phi_mux_j_14_flag_0_i_phi_fu_77_p6 = 1'd1;
    end else begin
        ap_phi_mux_j_14_flag_0_i_phi_fu_77_p6 = 'bx;
    end
end

always @ (*) begin
    if (((icmp_ln78_fu_141_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1))) begin
        if ((icmp_ln81_fu_154_p2 == 1'd0)) begin
            ap_phi_mux_j_14_new_0_i_phi_fu_91_p6 = add_ln80_fu_147_p2;
        end else if ((icmp_ln81_fu_154_p2 == 1'd1)) begin
            ap_phi_mux_j_14_new_0_i_phi_fu_91_p6 = 16'd0;
        end else begin
            ap_phi_mux_j_14_new_0_i_phi_fu_91_p6 = 'bx;
        end
    end else begin
        ap_phi_mux_j_14_new_0_i_phi_fu_91_p6 = 'bx;
    end
end

always @ (*) begin
    if (((icmp_ln78_fu_141_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_phi_mux_k_14_new_0_i_phi_fu_104_p6 = add_ln77_fu_134_p2;
    end else if ((((icmp_ln81_fu_154_p2 == 1'd0) & (icmp_ln78_fu_141_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1)) | ((icmp_ln81_fu_154_p2 == 1'd1) & (icmp_ln78_fu_141_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1)))) begin
        ap_phi_mux_k_14_new_0_i_phi_fu_104_p6 = 16'd0;
    end else begin
        ap_phi_mux_k_14_new_0_i_phi_fu_104_p6 = 'bx;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_0_blk_n = indices_0_full_n;
    end else begin
        indices_0_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_0_write = 1'b1;
    end else begin
        indices_0_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_1_blk_n = indices_1_full_n;
    end else begin
        indices_1_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_1_write = 1'b1;
    end else begin
        indices_1_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_2_out1_blk_n = indices_2_out1_full_n;
    end else begin
        indices_2_out1_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_2_out1_write = 1'b1;
    end else begin
        indices_2_out1_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_2_out_blk_n = indices_2_out_full_n;
    end else begin
        indices_2_out_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_2_out_write = 1'b1;
    end else begin
        indices_2_out_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        internal_ap_ready = 1'b1;
    end else begin
        internal_ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((start_full_n == 1'b0) & (start_once_reg == 1'b0))) begin
        real_start = 1'b0;
    end else begin
        real_start = ap_start;
    end
end

always @ (*) begin
    if (((real_start == 1'b1) & (start_once_reg == 1'b0))) begin
        start_write = 1'b1;
    end else begin
        start_write = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln77_fu_134_p2 = (k_2 + 16'd1);

assign add_ln80_fu_147_p2 = (j_2 + 16'd1);

assign add_ln83_fu_160_p2 = (i_2 + 16'd1);

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

always @ (*) begin
    ap_block_state1 = ((real_start == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1));
end

assign ap_ready = internal_ap_ready;

assign icmp_ln78_fu_141_p2 = ((add_ln77_fu_134_p2 == 16'd16) ? 1'b1 : 1'b0);

assign icmp_ln81_fu_154_p2 = ((add_ln80_fu_147_p2 == 16'd56) ? 1'b1 : 1'b0);

assign icmp_ln84_fu_166_p2 = ((add_ln83_fu_160_p2 == 16'd56) ? 1'b1 : 1'b0);

assign indices_0_din = i_2;

assign indices_1_din = j_2;

assign indices_2_out1_din = trunc_ln76_fu_128_p1;

assign indices_2_out_din = trunc_ln76_fu_128_p1;

assign select_ln84_fu_172_p3 = ((icmp_ln84_fu_166_p2[0:0] == 1'b1) ? 16'd0 : add_ln83_fu_160_p2);

assign start_out = real_start;

assign trunc_ln76_fu_128_p1 = k_2[3:0];

endmodule //td_fused_top_tdf3_get_next_ijk
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf3_readFilters30 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        filter_data_address0,
        filter_data_ce0,
        filter_data_q0,
        indices_23_dout,
        indices_23_empty_n,
        indices_23_read,
        weight_vecs_0_0_0_address0,
        weight_vecs_0_0_0_ce0,
        weight_vecs_0_0_0_we0,
        weight_vecs_0_0_0_d0
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state6 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [8:0] filter_data_address0;
output   filter_data_ce0;
input  [15:0] filter_data_q0;
input  [3:0] indices_23_dout;
input   indices_23_empty_n;
output   indices_23_read;
output  [4:0] weight_vecs_0_0_0_address0;
output   weight_vecs_0_0_0_ce0;
output   weight_vecs_0_0_0_we0;
output  [15:0] weight_vecs_0_0_0_d0;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg filter_data_ce0;
reg indices_23_read;
reg weight_vecs_0_0_0_ce0;
reg weight_vecs_0_0_0_we0;

reg    ap_done_reg;
  reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    indices_23_blk_n;
reg   [5:0] kk_0_0_i_i_reg_93;
reg   [5:0] kk_0_0_i_i_reg_93_pp0_iter1_reg;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
wire    ap_block_state4_pp0_stage0_iter2;
wire    ap_block_state5_pp0_stage0_iter3;
wire    ap_block_pp0_stage0_11001;
reg   [5:0] kk_0_0_i_i_reg_93_pp0_iter2_reg;
wire   [8:0] tmp_fu_105_p3;
reg   [8:0] tmp_reg_144;
wire   [5:0] add_ln49_fu_113_p2;
reg   [5:0] add_ln49_reg_149;
reg    ap_enable_reg_pp0_iter0;
wire   [0:0] icmp_ln49_fu_119_p2;
reg   [0:0] icmp_ln49_reg_154;
reg   [0:0] icmp_ln49_reg_154_pp0_iter1_reg;
reg   [0:0] icmp_ln49_reg_154_pp0_iter2_reg;
reg    ap_block_state1;
wire    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_exit_iter0_state2;
reg    ap_enable_reg_pp0_iter1;
reg    ap_enable_reg_pp0_iter2;
reg    ap_enable_reg_pp0_iter3;
reg   [5:0] ap_phi_mux_kk_0_0_i_i_phi_fu_97_p4;
wire    ap_block_pp0_stage0;
wire   [63:0] zext_ln55_39_fu_134_p1;
wire   [63:0] zext_ln49_fu_139_p1;
wire   [8:0] zext_ln55_fu_125_p1;
wire   [8:0] add_ln55_fu_129_p2;
wire    ap_CS_fsm_state6;
reg   [2:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state6)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_condition_pp0_exit_iter0_state2) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            if ((1'b1 == ap_condition_pp0_exit_iter0_state2)) begin
                ap_enable_reg_pp0_iter1 <= (1'b1 ^ ap_condition_pp0_exit_iter0_state2);
            end else if ((1'b1 == 1'b1)) begin
                ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
            end
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end else if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter3 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln49_reg_154 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        kk_0_0_i_i_reg_93 <= add_ln49_reg_149;
    end else if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        kk_0_0_i_i_reg_93 <= 6'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        add_ln49_reg_149 <= add_ln49_fu_113_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln49_reg_154 <= icmp_ln49_fu_119_p2;
        icmp_ln49_reg_154_pp0_iter1_reg <= icmp_ln49_reg_154;
        kk_0_0_i_i_reg_93_pp0_iter1_reg <= kk_0_0_i_i_reg_93;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        icmp_ln49_reg_154_pp0_iter2_reg <= icmp_ln49_reg_154_pp0_iter1_reg;
        kk_0_0_i_i_reg_93_pp0_iter2_reg <= kk_0_0_i_i_reg_93_pp0_iter1_reg;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state1)) begin
        tmp_reg_144[8 : 5] <= tmp_fu_105_p3[8 : 5];
    end
end

always @ (*) begin
    if ((icmp_ln49_fu_119_p2 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state2 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state2 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state6)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln49_reg_154 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_kk_0_0_i_i_phi_fu_97_p4 = add_ln49_reg_149;
    end else begin
        ap_phi_mux_kk_0_0_i_i_phi_fu_97_p4 = kk_0_0_i_i_reg_93;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state6)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter3 == 1'b1)))) begin
        filter_data_ce0 = 1'b1;
    end else begin
        filter_data_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_23_blk_n = indices_23_empty_n;
    end else begin
        indices_23_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_23_read = 1'b1;
    end else begin
        indices_23_read = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter3 == 1'b1))) begin
        weight_vecs_0_0_0_ce0 = 1'b1;
    end else begin
        weight_vecs_0_0_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln49_reg_154_pp0_iter2_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter3 == 1'b1))) begin
        weight_vecs_0_0_0_we0 = 1'b1;
    end else begin
        weight_vecs_0_0_0_we0 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((~((icmp_ln49_fu_119_p2 == 1'd1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter1 == 1'b0)) & ~((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter3 == 1'b1) & (ap_enable_reg_pp0_iter2 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if ((((icmp_ln49_fu_119_p2 == 1'd1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter1 == 1'b0)) | ((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter3 == 1'b1) & (ap_enable_reg_pp0_iter2 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_state6;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state6 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln49_fu_113_p2 = (ap_phi_mux_kk_0_0_i_i_phi_fu_97_p4 + 6'd1);

assign add_ln55_fu_129_p2 = (tmp_reg_144 + zext_ln55_fu_125_p1);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state6 = ap_CS_fsm[32'd2];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1));
end

assign ap_block_state2_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign filter_data_address0 = zext_ln55_39_fu_134_p1;

assign icmp_ln49_fu_119_p2 = ((ap_phi_mux_kk_0_0_i_i_phi_fu_97_p4 == 6'd32) ? 1'b1 : 1'b0);

assign tmp_fu_105_p3 = {{indices_23_dout}, {5'd0}};

assign weight_vecs_0_0_0_address0 = zext_ln49_fu_139_p1;

assign weight_vecs_0_0_0_d0 = filter_data_q0;

assign zext_ln49_fu_139_p1 = kk_0_0_i_i_reg_93_pp0_iter2_reg;

assign zext_ln55_39_fu_134_p1 = add_ln55_fu_129_p2;

assign zext_ln55_fu_125_p1 = ap_phi_mux_kk_0_0_i_i_phi_fu_97_p4;

always @ (posedge ap_clk) begin
    tmp_reg_144[4:0] <= 5'b00000;
end

endmodule //td_fused_top_tdf3_readFilters30
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf3_readInputs (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        in_data_address0,
        in_data_ce0,
        in_data_q0,
        indices_01_dout,
        indices_01_empty_n,
        indices_01_read,
        indices_12_dout,
        indices_12_empty_n,
        indices_12_read,
        ifmap_vec_0_0_address0,
        ifmap_vec_0_0_ce0,
        ifmap_vec_0_0_we0,
        ifmap_vec_0_0_d0,
        ifmap_vec_0_0_address1,
        ifmap_vec_0_0_ce1,
        ifmap_vec_0_0_we1,
        ifmap_vec_0_0_d1,
        indices_01_out_din,
        indices_01_out_full_n,
        indices_01_out_write,
        indices_12_out_din,
        indices_12_out_full_n,
        indices_12_out_write
);

parameter    ap_ST_fsm_state1 = 5'd1;
parameter    ap_ST_fsm_state2 = 5'd2;
parameter    ap_ST_fsm_pp0_stage0 = 5'd4;
parameter    ap_ST_fsm_pp0_stage1 = 5'd8;
parameter    ap_ST_fsm_state8 = 5'd16;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [14:0] in_data_address0;
output   in_data_ce0;
input  [63:0] in_data_q0;
input  [15:0] indices_01_dout;
input   indices_01_empty_n;
output   indices_01_read;
input  [15:0] indices_12_dout;
input   indices_12_empty_n;
output   indices_12_read;
output  [4:0] ifmap_vec_0_0_address0;
output   ifmap_vec_0_0_ce0;
output   ifmap_vec_0_0_we0;
output  [15:0] ifmap_vec_0_0_d0;
output  [4:0] ifmap_vec_0_0_address1;
output   ifmap_vec_0_0_ce1;
output   ifmap_vec_0_0_we1;
output  [15:0] ifmap_vec_0_0_d1;
output  [5:0] indices_01_out_din;
input   indices_01_out_full_n;
output   indices_01_out_write;
output  [11:0] indices_12_out_din;
input   indices_12_out_full_n;
output   indices_12_out_write;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg in_data_ce0;
reg indices_01_read;
reg indices_12_read;
reg[4:0] ifmap_vec_0_0_address0;
reg ifmap_vec_0_0_ce0;
reg ifmap_vec_0_0_we0;
reg[15:0] ifmap_vec_0_0_d0;
reg[4:0] ifmap_vec_0_0_address1;
reg ifmap_vec_0_0_ce1;
reg ifmap_vec_0_0_we1;
reg[15:0] ifmap_vec_0_0_d1;
reg indices_01_out_write;
reg indices_12_out_write;

reg    ap_done_reg;
  reg   [4:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    indices_01_blk_n;
reg    indices_12_blk_n;
reg    indices_01_out_blk_n;
reg    indices_12_out_blk_n;
reg   [5:0] kk_0_i_i_reg_178;
reg   [5:0] kk_0_i_i_reg_178_pp0_iter1_reg;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_block_state3_pp0_stage0_iter0;
wire    ap_block_state5_pp0_stage0_iter1;
wire    ap_block_state7_pp0_stage0_iter2;
wire    ap_block_pp0_stage0_11001;
wire   [5:0] trunc_ln135_fu_190_p1;
reg   [5:0] trunc_ln135_reg_432;
reg   [15:0] col_coord_reg_437;
wire   [0:0] is_padding_fu_212_p2;
reg   [0:0] is_padding_reg_442;
wire   [13:0] add_ln32_fu_272_p2;
reg   [13:0] add_ln32_reg_452;
wire    ap_CS_fsm_state2;
wire   [0:0] icmp_ln25_fu_278_p2;
reg   [0:0] icmp_ln25_reg_457;
reg   [0:0] icmp_ln25_reg_457_pp0_iter1_reg;
wire   [5:0] add_ln25_fu_306_p2;
reg   [5:0] add_ln25_reg_466;
wire    ap_CS_fsm_pp0_stage1;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_state4_pp0_stage1_iter0;
wire    ap_block_state6_pp0_stage1_iter1;
wire    ap_block_pp0_stage1_11001;
wire   [4:0] empty_104_fu_317_p1;
reg   [4:0] empty_104_reg_471;
wire   [15:0] select_ln33_20_fu_384_p3;
reg   [15:0] select_ln33_20_reg_477;
wire   [15:0] select_ln33_21_fu_405_p3;
reg   [15:0] select_ln33_21_reg_482;
wire    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_exit_iter0_state3;
reg    ap_enable_reg_pp0_iter1;
wire    ap_block_pp0_stage1_subdone;
reg    ap_enable_reg_pp0_iter2;
reg   [5:0] ap_phi_mux_kk_0_i_i_phi_fu_182_p4;
wire    ap_block_pp0_stage0;
wire   [63:0] sext_ln32_fu_301_p1;
wire   [63:0] kk_0_cast4_i_i_fu_312_p1;
wire    ap_block_pp0_stage1;
wire   [63:0] zext_ln32_16_fu_343_p1;
wire   [63:0] zext_ln32_17_fu_417_p1;
wire   [63:0] zext_ln32_18_fu_427_p1;
reg    ap_block_state1;
wire   [15:0] select_ln33_fu_329_p3;
wire   [15:0] select_ln33_19_fu_362_p3;
wire   [0:0] cmp7_i_i_fu_200_p2;
wire   [0:0] icmp_ln24_fu_206_p2;
wire   [5:0] empty_102_fu_218_p1;
wire   [5:0] row_coord_int_fu_221_p3;
wire   [11:0] tmp_fu_234_p3;
wire   [8:0] tmp_s_fu_246_p3;
wire   [12:0] zext_ln32_fu_242_p1;
wire   [12:0] zext_ln32_20_fu_254_p1;
wire   [12:0] sub_ln32_fu_258_p2;
wire   [5:0] col_coord_int_fu_227_p3;
wire   [13:0] sub_ln32_cast_fu_264_p1;
wire   [13:0] zext_ln32_21_fu_268_p1;
wire   [2:0] lshr_ln_fu_284_p4;
wire   [16:0] tmp_35_fu_294_p3;
wire   [15:0] trunc_ln32_fu_321_p1;
wire   [15:0] bitcast_ln32_fu_325_p1;
wire   [4:0] or_ln25_fu_337_p2;
wire   [15:0] tmp_58_i_i_fu_348_p4;
wire   [15:0] bitcast_ln32_19_fu_358_p1;
wire   [15:0] tmp_59_i_i_fu_370_p4;
wire   [15:0] bitcast_ln32_20_fu_380_p1;
wire   [15:0] tmp_60_i_i_fu_391_p4;
wire   [15:0] bitcast_ln32_21_fu_401_p1;
wire   [4:0] or_ln25_13_fu_412_p2;
wire   [4:0] or_ln25_14_fu_422_p2;
wire    ap_CS_fsm_state8;
reg   [4:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 5'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b1 == ap_condition_pp0_exit_iter0_state3))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1)) | ((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b0)))) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            ap_enable_reg_pp0_iter2 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln25_reg_457 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        kk_0_i_i_reg_178 <= add_ln25_reg_466;
    end else if ((1'b1 == ap_CS_fsm_state2)) begin
        kk_0_i_i_reg_178 <= 6'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln25_reg_457 == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
        add_ln25_reg_466 <= add_ln25_fu_306_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        add_ln32_reg_452 <= add_ln32_fu_272_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state1)) begin
        col_coord_reg_437 <= indices_12_dout;
        is_padding_reg_442 <= is_padding_fu_212_p2;
        trunc_ln135_reg_432 <= trunc_ln135_fu_190_p1;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln25_reg_457_pp0_iter1_reg == 1'd0))) begin
        empty_104_reg_471 <= empty_104_fu_317_p1;
        select_ln33_20_reg_477 <= select_ln33_20_fu_384_p3;
        select_ln33_21_reg_482 <= select_ln33_21_fu_405_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln25_reg_457 <= icmp_ln25_fu_278_p2;
        icmp_ln25_reg_457_pp0_iter1_reg <= icmp_ln25_reg_457;
        kk_0_i_i_reg_178_pp0_iter1_reg <= kk_0_i_i_reg_178;
    end
end

always @ (*) begin
    if ((icmp_ln25_fu_278_p2 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state3 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state3 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state8)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln25_reg_457 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_kk_0_i_i_phi_fu_182_p4 = add_ln25_reg_466;
    end else begin
        ap_phi_mux_kk_0_i_i_phi_fu_182_p4 = kk_0_i_i_reg_178;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state8)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        ifmap_vec_0_0_address0 = zext_ln32_18_fu_427_p1;
    end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ifmap_vec_0_0_address0 = zext_ln32_16_fu_343_p1;
    end else begin
        ifmap_vec_0_0_address0 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        ifmap_vec_0_0_address1 = zext_ln32_17_fu_417_p1;
    end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ifmap_vec_0_0_address1 = kk_0_cast4_i_i_fu_312_p1;
    end else begin
        ifmap_vec_0_0_address1 = 'bx;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1)) | ((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1)))) begin
        ifmap_vec_0_0_ce0 = 1'b1;
    end else begin
        ifmap_vec_0_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1)) | ((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1)))) begin
        ifmap_vec_0_0_ce1 = 1'b1;
    end else begin
        ifmap_vec_0_0_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        ifmap_vec_0_0_d0 = select_ln33_21_reg_482;
    end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ifmap_vec_0_0_d0 = select_ln33_19_fu_362_p3;
    end else begin
        ifmap_vec_0_0_d0 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        ifmap_vec_0_0_d1 = select_ln33_20_reg_477;
    end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ifmap_vec_0_0_d1 = select_ln33_fu_329_p3;
    end else begin
        ifmap_vec_0_0_d1 = 'bx;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1) & (icmp_ln25_reg_457_pp0_iter1_reg == 1'd0)) | ((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln25_reg_457_pp0_iter1_reg == 1'd0)))) begin
        ifmap_vec_0_0_we0 = 1'b1;
    end else begin
        ifmap_vec_0_0_we0 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1) & (icmp_ln25_reg_457_pp0_iter1_reg == 1'd0)) | ((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln25_reg_457_pp0_iter1_reg == 1'd0)))) begin
        ifmap_vec_0_0_we1 = 1'b1;
    end else begin
        ifmap_vec_0_0_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1)) | ((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1)) | ((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1)) | ((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1)))) begin
        in_data_ce0 = 1'b1;
    end else begin
        in_data_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_01_blk_n = indices_01_empty_n;
    end else begin
        indices_01_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_01_out_blk_n = indices_01_out_full_n;
    end else begin
        indices_01_out_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((indices_12_out_full_n == 1'b0) | (indices_01_out_full_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_01_out_write = 1'b1;
    end else begin
        indices_01_out_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((indices_12_out_full_n == 1'b0) | (indices_01_out_full_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_01_read = 1'b1;
    end else begin
        indices_01_read = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_12_blk_n = indices_12_empty_n;
    end else begin
        indices_12_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_12_out_blk_n = indices_12_out_full_n;
    end else begin
        indices_12_out_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((indices_12_out_full_n == 1'b0) | (indices_01_out_full_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_12_out_write = 1'b1;
    end else begin
        indices_12_out_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((indices_12_out_full_n == 1'b0) | (indices_01_out_full_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_12_read = 1'b1;
    end else begin
        indices_12_read = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((indices_12_out_full_n == 1'b0) | (indices_01_out_full_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_state2 : begin
            ap_NS_fsm = ap_ST_fsm_pp0_stage0;
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((~((icmp_ln25_fu_278_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1)) & ~((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0)) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end else if ((((icmp_ln25_fu_278_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1)) | ((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_state8;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_pp0_stage1 : begin
            if ((1'b0 == ap_block_pp0_stage1_subdone)) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end
        end
        ap_ST_fsm_state8 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln25_fu_306_p2 = (kk_0_i_i_reg_178 + 6'd4);

assign add_ln32_fu_272_p2 = ((sub_ln32_cast_fu_264_p1) + (zext_ln32_21_fu_268_p1));

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_pp0_stage1 = ap_CS_fsm[32'd3];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state8 = ap_CS_fsm[32'd4];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((indices_12_out_full_n == 1'b0) | (indices_01_out_full_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0));
end

assign ap_block_state3_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage1_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage1_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign bitcast_ln32_19_fu_358_p1 = tmp_58_i_i_fu_348_p4;

assign bitcast_ln32_20_fu_380_p1 = tmp_59_i_i_fu_370_p4;

assign bitcast_ln32_21_fu_401_p1 = tmp_60_i_i_fu_391_p4;

assign bitcast_ln32_fu_325_p1 = trunc_ln32_fu_321_p1;

assign cmp7_i_i_fu_200_p2 = ((indices_01_dout > 16'd55) ? 1'b1 : 1'b0);

assign col_coord_int_fu_227_p3 = ((is_padding_reg_442[0:0] == 1'b1) ? 6'd0 : empty_102_fu_218_p1);

assign empty_102_fu_218_p1 = col_coord_reg_437[5:0];

assign empty_104_fu_317_p1 = kk_0_i_i_reg_178_pp0_iter1_reg[4:0];

assign icmp_ln24_fu_206_p2 = ((indices_12_dout > 16'd55) ? 1'b1 : 1'b0);

assign icmp_ln25_fu_278_p2 = ((ap_phi_mux_kk_0_i_i_phi_fu_182_p4 == 6'd32) ? 1'b1 : 1'b0);

assign in_data_address0 = sext_ln32_fu_301_p1;

assign indices_01_out_din = indices_01_dout[5:0];

assign indices_12_out_din = indices_12_dout[11:0];

assign is_padding_fu_212_p2 = (icmp_ln24_fu_206_p2 | cmp7_i_i_fu_200_p2);

assign kk_0_cast4_i_i_fu_312_p1 = kk_0_i_i_reg_178_pp0_iter1_reg;

assign lshr_ln_fu_284_p4 = {{ap_phi_mux_kk_0_i_i_phi_fu_182_p4[4:2]}};

assign or_ln25_13_fu_412_p2 = (empty_104_reg_471 | 5'd2);

assign or_ln25_14_fu_422_p2 = (empty_104_reg_471 | 5'd3);

assign or_ln25_fu_337_p2 = (empty_104_fu_317_p1 | 5'd1);

assign row_coord_int_fu_221_p3 = ((is_padding_reg_442[0:0] == 1'b1) ? 6'd0 : trunc_ln135_reg_432);

assign select_ln33_19_fu_362_p3 = ((is_padding_reg_442[0:0] == 1'b1) ? 16'd0 : bitcast_ln32_19_fu_358_p1);

assign select_ln33_20_fu_384_p3 = ((is_padding_reg_442[0:0] == 1'b1) ? 16'd0 : bitcast_ln32_20_fu_380_p1);

assign select_ln33_21_fu_405_p3 = ((is_padding_reg_442[0:0] == 1'b1) ? 16'd0 : bitcast_ln32_21_fu_401_p1);

assign select_ln33_fu_329_p3 = ((is_padding_reg_442[0:0] == 1'b1) ? 16'd0 : bitcast_ln32_fu_325_p1);

assign sext_ln32_fu_301_p1 = (tmp_35_fu_294_p3);

assign sub_ln32_cast_fu_264_p1 = (sub_ln32_fu_258_p2);

assign sub_ln32_fu_258_p2 = (zext_ln32_fu_242_p1 - zext_ln32_20_fu_254_p1);

assign tmp_35_fu_294_p3 = {{add_ln32_reg_452}, {lshr_ln_fu_284_p4}};

assign tmp_58_i_i_fu_348_p4 = {{in_data_q0[31:16]}};

assign tmp_59_i_i_fu_370_p4 = {{in_data_q0[47:32]}};

assign tmp_60_i_i_fu_391_p4 = {{in_data_q0[63:48]}};

assign tmp_fu_234_p3 = {{row_coord_int_fu_221_p3}, {6'd0}};

assign tmp_s_fu_246_p3 = {{row_coord_int_fu_221_p3}, {3'd0}};

assign trunc_ln135_fu_190_p1 = indices_01_dout[5:0];

assign trunc_ln32_fu_321_p1 = in_data_q0[15:0];

assign zext_ln32_16_fu_343_p1 = or_ln25_fu_337_p2;

assign zext_ln32_17_fu_417_p1 = or_ln25_13_fu_412_p2;

assign zext_ln32_18_fu_427_p1 = or_ln25_14_fu_422_p2;

assign zext_ln32_20_fu_254_p1 = tmp_s_fu_246_p3;

assign zext_ln32_21_fu_268_p1 = col_coord_int_fu_227_p3;

assign zext_ln32_fu_242_p1 = tmp_fu_234_p3;

endmodule //td_fused_top_tdf3_readInputs
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf3_writeOutputs_unaligned (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        indices_01_dout,
        indices_01_empty_n,
        indices_01_read,
        indices_12_dout,
        indices_12_empty_n,
        indices_12_read,
        p_read,
        out_data_address1,
        out_data_ce1,
        out_data_we1,
        out_data_d1
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_state2 = 3'd2;
parameter    ap_ST_fsm_state3 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
input  [5:0] indices_01_dout;
input   indices_01_empty_n;
output   indices_01_read;
input  [11:0] indices_12_dout;
input   indices_12_empty_n;
output   indices_12_read;
input  [15:0] p_read;
output  [13:0] out_data_address1;
output   out_data_ce1;
output   out_data_we1;
output  [63:0] out_data_d1;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg indices_01_read;
reg indices_12_read;
reg out_data_ce1;
reg out_data_we1;

reg    ap_done_reg;
  reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg   [15:0] outputCount_6;
reg   [15:0] outputChanIdx_6;
reg   [15:0] outputRow_10_0;
reg   [15:0] outputRow_10_1;
reg   [15:0] outputRow_10_2;
reg   [15:0] outputRow_10_3;
reg    indices_01_blk_n;
reg    indices_12_blk_n;
wire   [13:0] shl_ln89_fu_163_p2;
reg   [13:0] shl_ln89_reg_312;
wire   [15:0] add_ln87_fu_201_p2;
wire    ap_CS_fsm_state2;
wire   [0:0] icmp_ln88_fu_207_p2;
reg   [0:0] icmp_ln88_reg_325;
reg   [15:0] ap_phi_mux_empty_phi_fu_112_p4;
reg   [15:0] empty_reg_109;
wire    ap_CS_fsm_state3;
wire   [63:0] zext_ln94_12_fu_234_p1;
wire   [15:0] select_ln97_fu_292_p3;
wire   [1:0] trunc_ln86_fu_173_p1;
reg   [15:0] ap_sig_allocacmp_outputRow_10_0_load;
reg   [15:0] ap_sig_allocacmp_outputRow_10_1_load;
reg   [15:0] ap_sig_allocacmp_outputRow_10_2_load;
reg   [15:0] ap_sig_allocacmp_outputRow_10_3_load;
reg    ap_block_state1;
wire   [11:0] tmp_fu_119_p3;
wire   [8:0] tmp_s_fu_131_p3;
wire   [12:0] zext_ln94_fu_127_p1;
wire   [12:0] zext_ln94_9_fu_139_p1;
wire   [12:0] sub_ln94_fu_143_p2;
wire   [13:0] sub_ln94_cast13_fu_149_p1;
wire   [13:0] zext_ln94_10_fu_153_p1;
wire   [13:0] add_ln94_fu_157_p2;
wire   [3:0] trunc_ln94_fu_221_p1;
wire   [13:0] zext_ln94_11_fu_225_p1;
wire   [13:0] add_ln94_5_fu_229_p2;
wire   [15:0] bitcast_ln94_15_fu_263_p1;
wire   [15:0] bitcast_ln94_14_fu_255_p1;
wire   [15:0] bitcast_ln94_13_fu_247_p1;
wire   [15:0] bitcast_ln94_fu_239_p1;
wire   [15:0] add_ln96_fu_280_p2;
wire   [0:0] icmp_ln97_fu_286_p2;
reg   [2:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 3'd1;
#0 outputCount_6 = 16'd0;
#0 outputChanIdx_6 = 16'd0;
#0 outputRow_10_0 = 16'd0;
#0 outputRow_10_1 = 16'd0;
#0 outputRow_10_2 = 16'd0;
#0 outputRow_10_3 = 16'd0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state3)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln88_reg_325 == 1'd1) & (1'b1 == ap_CS_fsm_state3))) begin
        empty_reg_109 <= 16'd0;
    end else if (((icmp_ln88_fu_207_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state2))) begin
        empty_reg_109 <= add_ln87_fu_201_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        icmp_ln88_reg_325 <= icmp_ln88_fu_207_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln88_fu_207_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        outputChanIdx_6 <= select_ln97_fu_292_p3;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state3)) begin
        outputCount_6 <= ap_phi_mux_empty_phi_fu_112_p4;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln86_fu_173_p1 == 2'd0) & (1'b1 == ap_CS_fsm_state2))) begin
        outputRow_10_0 <= p_read;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln86_fu_173_p1 == 2'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        outputRow_10_1 <= p_read;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln86_fu_173_p1 == 2'd2) & (1'b1 == ap_CS_fsm_state2))) begin
        outputRow_10_2 <= p_read;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln86_fu_173_p1 == 2'd3) & (1'b1 == ap_CS_fsm_state2))) begin
        outputRow_10_3 <= p_read;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state1)) begin
        shl_ln89_reg_312[13 : 2] <= shl_ln89_fu_163_p2[13 : 2];
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state3)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln88_reg_325 == 1'd1) & (1'b1 == ap_CS_fsm_state3))) begin
        ap_phi_mux_empty_phi_fu_112_p4 = 16'd0;
    end else begin
        ap_phi_mux_empty_phi_fu_112_p4 = empty_reg_109;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state3)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((trunc_ln86_fu_173_p1 == 2'd0) & (1'b1 == ap_CS_fsm_state2))) begin
        ap_sig_allocacmp_outputRow_10_0_load = p_read;
    end else begin
        ap_sig_allocacmp_outputRow_10_0_load = outputRow_10_0;
    end
end

always @ (*) begin
    if (((trunc_ln86_fu_173_p1 == 2'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        ap_sig_allocacmp_outputRow_10_1_load = p_read;
    end else begin
        ap_sig_allocacmp_outputRow_10_1_load = outputRow_10_1;
    end
end

always @ (*) begin
    if (((trunc_ln86_fu_173_p1 == 2'd2) & (1'b1 == ap_CS_fsm_state2))) begin
        ap_sig_allocacmp_outputRow_10_2_load = p_read;
    end else begin
        ap_sig_allocacmp_outputRow_10_2_load = outputRow_10_2;
    end
end

always @ (*) begin
    if (((trunc_ln86_fu_173_p1 == 2'd3) & (1'b1 == ap_CS_fsm_state2))) begin
        ap_sig_allocacmp_outputRow_10_3_load = p_read;
    end else begin
        ap_sig_allocacmp_outputRow_10_3_load = outputRow_10_3;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_01_blk_n = indices_01_empty_n;
    end else begin
        indices_01_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_01_read = 1'b1;
    end else begin
        indices_01_read = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_12_blk_n = indices_12_empty_n;
    end else begin
        indices_12_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_12_read = 1'b1;
    end else begin
        indices_12_read = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state2))) begin
        out_data_ce1 = 1'b1;
    end else begin
        out_data_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln88_fu_207_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        out_data_we1 = 1'b1;
    end else begin
        out_data_we1 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_start == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_state2 : begin
            ap_NS_fsm = ap_ST_fsm_state3;
        end
        ap_ST_fsm_state3 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln87_fu_201_p2 = (outputCount_6 + 16'd1);

assign add_ln94_5_fu_229_p2 = (shl_ln89_reg_312 + zext_ln94_11_fu_225_p1);

assign add_ln94_fu_157_p2 = (sub_ln94_cast13_fu_149_p1 + zext_ln94_10_fu_153_p1);

assign add_ln96_fu_280_p2 = (outputChanIdx_6 + 16'd1);

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1));
end

assign bitcast_ln94_13_fu_247_p1 = ap_sig_allocacmp_outputRow_10_1_load;

assign bitcast_ln94_14_fu_255_p1 = ap_sig_allocacmp_outputRow_10_2_load;

assign bitcast_ln94_15_fu_263_p1 = ap_sig_allocacmp_outputRow_10_3_load;

assign bitcast_ln94_fu_239_p1 = ap_sig_allocacmp_outputRow_10_0_load;

assign icmp_ln88_fu_207_p2 = ((add_ln87_fu_201_p2 == 16'd4) ? 1'b1 : 1'b0);

assign icmp_ln97_fu_286_p2 = ((add_ln96_fu_280_p2 == 16'd4) ? 1'b1 : 1'b0);

assign out_data_address1 = zext_ln94_12_fu_234_p1;

assign out_data_d1 = {{{{bitcast_ln94_15_fu_263_p1}, {bitcast_ln94_14_fu_255_p1}}, {bitcast_ln94_13_fu_247_p1}}, {bitcast_ln94_fu_239_p1}};

assign select_ln97_fu_292_p3 = ((icmp_ln97_fu_286_p2[0:0] == 1'b1) ? 16'd0 : add_ln96_fu_280_p2);

assign shl_ln89_fu_163_p2 = add_ln94_fu_157_p2 << 14'd2;

assign sub_ln94_cast13_fu_149_p1 = sub_ln94_fu_143_p2;

assign sub_ln94_fu_143_p2 = (zext_ln94_fu_127_p1 - zext_ln94_9_fu_139_p1);

assign tmp_fu_119_p3 = {{indices_01_dout}, {6'd0}};

assign tmp_s_fu_131_p3 = {{indices_01_dout}, {3'd0}};

assign trunc_ln86_fu_173_p1 = outputCount_6[1:0];

assign trunc_ln94_fu_221_p1 = outputChanIdx_6[3:0];

assign zext_ln94_10_fu_153_p1 = indices_12_dout;

assign zext_ln94_11_fu_225_p1 = trunc_ln94_fu_221_p1;

assign zext_ln94_12_fu_234_p1 = add_ln94_5_fu_229_p2;

assign zext_ln94_9_fu_139_p1 = tmp_s_fu_131_p3;

assign zext_ln94_fu_127_p1 = tmp_fu_119_p3;

always @ (posedge ap_clk) begin
    shl_ln89_reg_312[1:0] <= 2'b00;
end

endmodule //td_fused_top_tdf3_writeOutputs_unaligned
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf4_111 (
        in_data_address0,
        in_data_ce0,
        in_data_d0,
        in_data_q0,
        in_data_we0,
        in_data_address1,
        in_data_ce1,
        in_data_d1,
        in_data_q1,
        in_data_we1,
        out_data_address0,
        out_data_ce0,
        out_data_d0,
        out_data_q0,
        out_data_we0,
        out_data_address1,
        out_data_ce1,
        out_data_d1,
        out_data_q1,
        out_data_we1,
        l1_filter_data_address0,
        l1_filter_data_ce0,
        l1_filter_data_d0,
        l1_filter_data_q0,
        l1_filter_data_we0,
        l1_filter_data_address1,
        l1_filter_data_ce1,
        l1_filter_data_d1,
        l1_filter_data_q1,
        l1_filter_data_we1,
        l2_filter_data_address0,
        l2_filter_data_ce0,
        l2_filter_data_d0,
        l2_filter_data_q0,
        l2_filter_data_we0,
        l2_filter_data_address1,
        l2_filter_data_ce1,
        l2_filter_data_d1,
        l2_filter_data_q1,
        l2_filter_data_we1,
        l1_adjustments_address0,
        l1_adjustments_ce0,
        l1_adjustments_d0,
        l1_adjustments_q0,
        l1_adjustments_we0,
        l1_adjustments_address1,
        l1_adjustments_ce1,
        l1_adjustments_d1,
        l1_adjustments_q1,
        l1_adjustments_we1,
        l2_adjustments_address0,
        l2_adjustments_ce0,
        l2_adjustments_d0,
        l2_adjustments_q0,
        l2_adjustments_we0,
        l2_adjustments_address1,
        l2_adjustments_ce1,
        l2_adjustments_d1,
        l2_adjustments_q1,
        l2_adjustments_we1,
        ap_clk,
        ap_rst,
        in_data_empty_n,
        in_data_read,
        out_data_full_n,
        out_data_write,
        ap_start,
        ap_done,
        ap_ready,
        ap_idle,
        ap_continue
);


output  [13:0] in_data_address0;
output   in_data_ce0;
output  [63:0] in_data_d0;
input  [63:0] in_data_q0;
output   in_data_we0;
output  [13:0] in_data_address1;
output   in_data_ce1;
output  [63:0] in_data_d1;
input  [63:0] in_data_q1;
output   in_data_we1;
output  [13:0] out_data_address0;
output   out_data_ce0;
output  [63:0] out_data_d0;
input  [63:0] out_data_q0;
output   out_data_we0;
output  [13:0] out_data_address1;
output   out_data_ce1;
output  [63:0] out_data_d1;
input  [63:0] out_data_q1;
output   out_data_we1;
output  [14:0] l1_filter_data_address0;
output   l1_filter_data_ce0;
output  [15:0] l1_filter_data_d0;
input  [15:0] l1_filter_data_q0;
output   l1_filter_data_we0;
output  [14:0] l1_filter_data_address1;
output   l1_filter_data_ce1;
output  [15:0] l1_filter_data_d1;
input  [15:0] l1_filter_data_q1;
output   l1_filter_data_we1;
output  [10:0] l2_filter_data_address0;
output   l2_filter_data_ce0;
output  [15:0] l2_filter_data_d0;
input  [15:0] l2_filter_data_q0;
output   l2_filter_data_we0;
output  [10:0] l2_filter_data_address1;
output   l2_filter_data_ce1;
output  [15:0] l2_filter_data_d1;
input  [15:0] l2_filter_data_q1;
output   l2_filter_data_we1;
output  [6:0] l1_adjustments_address0;
output   l1_adjustments_ce0;
output  [47:0] l1_adjustments_d0;
input  [47:0] l1_adjustments_q0;
output   l1_adjustments_we0;
output  [6:0] l1_adjustments_address1;
output   l1_adjustments_ce1;
output  [47:0] l1_adjustments_d1;
input  [47:0] l1_adjustments_q1;
output   l1_adjustments_we1;
output  [3:0] l2_adjustments_address0;
output   l2_adjustments_ce0;
output  [47:0] l2_adjustments_d0;
input  [47:0] l2_adjustments_q0;
output   l2_adjustments_we0;
output  [3:0] l2_adjustments_address1;
output   l2_adjustments_ce1;
output  [47:0] l2_adjustments_d1;
input  [47:0] l2_adjustments_q1;
output   l2_adjustments_we1;
input   ap_clk;
input   ap_rst;
input   in_data_empty_n;
output   in_data_read;
input   out_data_full_n;
output   out_data_write;
input   ap_start;
output   ap_done;
output   ap_ready;
output   ap_idle;
input   ap_continue;

reg ap_done;
reg ap_ready;
reg ap_idle;

wire   [13:0] dataflow_in_loop_TOP_LOOP37832_U0_in_data_address0;
wire    dataflow_in_loop_TOP_LOOP37832_U0_in_data_ce0;
wire   [63:0] dataflow_in_loop_TOP_LOOP37832_U0_in_data_d0;
wire    dataflow_in_loop_TOP_LOOP37832_U0_in_data_we0;
wire   [13:0] dataflow_in_loop_TOP_LOOP37832_U0_in_data_address1;
wire    dataflow_in_loop_TOP_LOOP37832_U0_in_data_ce1;
wire   [63:0] dataflow_in_loop_TOP_LOOP37832_U0_in_data_d1;
wire    dataflow_in_loop_TOP_LOOP37832_U0_in_data_we1;
wire   [14:0] dataflow_in_loop_TOP_LOOP37832_U0_l1_filter_data_address0;
wire    dataflow_in_loop_TOP_LOOP37832_U0_l1_filter_data_ce0;
wire   [15:0] dataflow_in_loop_TOP_LOOP37832_U0_l1_filter_data_d0;
wire    dataflow_in_loop_TOP_LOOP37832_U0_l1_filter_data_we0;
wire   [14:0] dataflow_in_loop_TOP_LOOP37832_U0_l1_filter_data_address1;
wire    dataflow_in_loop_TOP_LOOP37832_U0_l1_filter_data_ce1;
wire   [15:0] dataflow_in_loop_TOP_LOOP37832_U0_l1_filter_data_d1;
wire    dataflow_in_loop_TOP_LOOP37832_U0_l1_filter_data_we1;
wire   [6:0] dataflow_in_loop_TOP_LOOP37832_U0_l1_adjustments_address0;
wire    dataflow_in_loop_TOP_LOOP37832_U0_l1_adjustments_ce0;
wire   [47:0] dataflow_in_loop_TOP_LOOP37832_U0_l1_adjustments_d0;
wire    dataflow_in_loop_TOP_LOOP37832_U0_l1_adjustments_we0;
wire   [6:0] dataflow_in_loop_TOP_LOOP37832_U0_l1_adjustments_address1;
wire    dataflow_in_loop_TOP_LOOP37832_U0_l1_adjustments_ce1;
wire   [47:0] dataflow_in_loop_TOP_LOOP37832_U0_l1_adjustments_d1;
wire    dataflow_in_loop_TOP_LOOP37832_U0_l1_adjustments_we1;
wire   [10:0] dataflow_in_loop_TOP_LOOP37832_U0_l2_filter_data_address0;
wire    dataflow_in_loop_TOP_LOOP37832_U0_l2_filter_data_ce0;
wire   [15:0] dataflow_in_loop_TOP_LOOP37832_U0_l2_filter_data_d0;
wire    dataflow_in_loop_TOP_LOOP37832_U0_l2_filter_data_we0;
wire   [10:0] dataflow_in_loop_TOP_LOOP37832_U0_l2_filter_data_address1;
wire    dataflow_in_loop_TOP_LOOP37832_U0_l2_filter_data_ce1;
wire   [15:0] dataflow_in_loop_TOP_LOOP37832_U0_l2_filter_data_d1;
wire    dataflow_in_loop_TOP_LOOP37832_U0_l2_filter_data_we1;
wire   [13:0] dataflow_in_loop_TOP_LOOP37832_U0_out_data_address0;
wire    dataflow_in_loop_TOP_LOOP37832_U0_out_data_ce0;
wire   [63:0] dataflow_in_loop_TOP_LOOP37832_U0_out_data_d0;
wire    dataflow_in_loop_TOP_LOOP37832_U0_out_data_we0;
wire   [13:0] dataflow_in_loop_TOP_LOOP37832_U0_out_data_address1;
wire    dataflow_in_loop_TOP_LOOP37832_U0_out_data_ce1;
wire   [63:0] dataflow_in_loop_TOP_LOOP37832_U0_out_data_d1;
wire    dataflow_in_loop_TOP_LOOP37832_U0_out_data_we1;
wire   [3:0] dataflow_in_loop_TOP_LOOP37832_U0_l2_adjustments_address0;
wire    dataflow_in_loop_TOP_LOOP37832_U0_l2_adjustments_ce0;
wire   [47:0] dataflow_in_loop_TOP_LOOP37832_U0_l2_adjustments_d0;
wire    dataflow_in_loop_TOP_LOOP37832_U0_l2_adjustments_we0;
wire   [3:0] dataflow_in_loop_TOP_LOOP37832_U0_l2_adjustments_address1;
wire    dataflow_in_loop_TOP_LOOP37832_U0_l2_adjustments_ce1;
wire   [47:0] dataflow_in_loop_TOP_LOOP37832_U0_l2_adjustments_d1;
wire    dataflow_in_loop_TOP_LOOP37832_U0_l2_adjustments_we1;
wire    dataflow_in_loop_TOP_LOOP37832_U0_ap_start;
wire    dataflow_in_loop_TOP_LOOP37832_U0_in_data_read;
wire    dataflow_in_loop_TOP_LOOP37832_U0_out_data_write;
wire    dataflow_in_loop_TOP_LOOP37832_U0_ap_done;
wire    dataflow_in_loop_TOP_LOOP37832_U0_ap_ready;
wire    dataflow_in_loop_TOP_LOOP37832_U0_ap_idle;
reg    dataflow_in_loop_TOP_LOOP37832_U0_ap_continue;
wire    dataflow_in_loop_TOP_LOOP37832_U0_in_data_full_n;
wire    dataflow_in_loop_TOP_LOOP37832_U0_in_data_write;
wire    ap_sync_continue;
wire    ap_sync_done;
wire    ap_sync_ready;
reg   [18:0] loop_dataflow_input_count;
reg   [18:0] loop_dataflow_output_count;
wire   [18:0] bound_minus_1;
wire    dataflow_in_loop_TOP_LOOP37832_U0_start_full_n;
wire    dataflow_in_loop_TOP_LOOP37832_U0_start_write;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 loop_dataflow_input_count = 19'd0;
#0 loop_dataflow_output_count = 19'd0;
end

td_fused_top_dataflow_in_loop_TOP_LOOP37832 dataflow_in_loop_TOP_LOOP37832_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .in_data_address0(dataflow_in_loop_TOP_LOOP37832_U0_in_data_address0),
    .in_data_ce0(dataflow_in_loop_TOP_LOOP37832_U0_in_data_ce0),
    .in_data_d0(dataflow_in_loop_TOP_LOOP37832_U0_in_data_d0),
    .in_data_q0(in_data_q0),
    .in_data_we0(dataflow_in_loop_TOP_LOOP37832_U0_in_data_we0),
    .in_data_address1(dataflow_in_loop_TOP_LOOP37832_U0_in_data_address1),
    .in_data_ce1(dataflow_in_loop_TOP_LOOP37832_U0_in_data_ce1),
    .in_data_d1(dataflow_in_loop_TOP_LOOP37832_U0_in_data_d1),
    .in_data_q1(64'd0),
    .in_data_we1(dataflow_in_loop_TOP_LOOP37832_U0_in_data_we1),
    .l1_filter_data_address0(dataflow_in_loop_TOP_LOOP37832_U0_l1_filter_data_address0),
    .l1_filter_data_ce0(dataflow_in_loop_TOP_LOOP37832_U0_l1_filter_data_ce0),
    .l1_filter_data_d0(dataflow_in_loop_TOP_LOOP37832_U0_l1_filter_data_d0),
    .l1_filter_data_q0(l1_filter_data_q0),
    .l1_filter_data_we0(dataflow_in_loop_TOP_LOOP37832_U0_l1_filter_data_we0),
    .l1_filter_data_address1(dataflow_in_loop_TOP_LOOP37832_U0_l1_filter_data_address1),
    .l1_filter_data_ce1(dataflow_in_loop_TOP_LOOP37832_U0_l1_filter_data_ce1),
    .l1_filter_data_d1(dataflow_in_loop_TOP_LOOP37832_U0_l1_filter_data_d1),
    .l1_filter_data_q1(16'd0),
    .l1_filter_data_we1(dataflow_in_loop_TOP_LOOP37832_U0_l1_filter_data_we1),
    .l1_adjustments_address0(dataflow_in_loop_TOP_LOOP37832_U0_l1_adjustments_address0),
    .l1_adjustments_ce0(dataflow_in_loop_TOP_LOOP37832_U0_l1_adjustments_ce0),
    .l1_adjustments_d0(dataflow_in_loop_TOP_LOOP37832_U0_l1_adjustments_d0),
    .l1_adjustments_q0(l1_adjustments_q0),
    .l1_adjustments_we0(dataflow_in_loop_TOP_LOOP37832_U0_l1_adjustments_we0),
    .l1_adjustments_address1(dataflow_in_loop_TOP_LOOP37832_U0_l1_adjustments_address1),
    .l1_adjustments_ce1(dataflow_in_loop_TOP_LOOP37832_U0_l1_adjustments_ce1),
    .l1_adjustments_d1(dataflow_in_loop_TOP_LOOP37832_U0_l1_adjustments_d1),
    .l1_adjustments_q1(48'd0),
    .l1_adjustments_we1(dataflow_in_loop_TOP_LOOP37832_U0_l1_adjustments_we1),
    .l2_filter_data_address0(dataflow_in_loop_TOP_LOOP37832_U0_l2_filter_data_address0),
    .l2_filter_data_ce0(dataflow_in_loop_TOP_LOOP37832_U0_l2_filter_data_ce0),
    .l2_filter_data_d0(dataflow_in_loop_TOP_LOOP37832_U0_l2_filter_data_d0),
    .l2_filter_data_q0(l2_filter_data_q0),
    .l2_filter_data_we0(dataflow_in_loop_TOP_LOOP37832_U0_l2_filter_data_we0),
    .l2_filter_data_address1(dataflow_in_loop_TOP_LOOP37832_U0_l2_filter_data_address1),
    .l2_filter_data_ce1(dataflow_in_loop_TOP_LOOP37832_U0_l2_filter_data_ce1),
    .l2_filter_data_d1(dataflow_in_loop_TOP_LOOP37832_U0_l2_filter_data_d1),
    .l2_filter_data_q1(16'd0),
    .l2_filter_data_we1(dataflow_in_loop_TOP_LOOP37832_U0_l2_filter_data_we1),
    .out_data_address0(dataflow_in_loop_TOP_LOOP37832_U0_out_data_address0),
    .out_data_ce0(dataflow_in_loop_TOP_LOOP37832_U0_out_data_ce0),
    .out_data_d0(dataflow_in_loop_TOP_LOOP37832_U0_out_data_d0),
    .out_data_q0(64'd0),
    .out_data_we0(dataflow_in_loop_TOP_LOOP37832_U0_out_data_we0),
    .out_data_address1(dataflow_in_loop_TOP_LOOP37832_U0_out_data_address1),
    .out_data_ce1(dataflow_in_loop_TOP_LOOP37832_U0_out_data_ce1),
    .out_data_d1(dataflow_in_loop_TOP_LOOP37832_U0_out_data_d1),
    .out_data_q1(64'd0),
    .out_data_we1(dataflow_in_loop_TOP_LOOP37832_U0_out_data_we1),
    .l2_adjustments_address0(dataflow_in_loop_TOP_LOOP37832_U0_l2_adjustments_address0),
    .l2_adjustments_ce0(dataflow_in_loop_TOP_LOOP37832_U0_l2_adjustments_ce0),
    .l2_adjustments_d0(dataflow_in_loop_TOP_LOOP37832_U0_l2_adjustments_d0),
    .l2_adjustments_q0(l2_adjustments_q0),
    .l2_adjustments_we0(dataflow_in_loop_TOP_LOOP37832_U0_l2_adjustments_we0),
    .l2_adjustments_address1(dataflow_in_loop_TOP_LOOP37832_U0_l2_adjustments_address1),
    .l2_adjustments_ce1(dataflow_in_loop_TOP_LOOP37832_U0_l2_adjustments_ce1),
    .l2_adjustments_d1(dataflow_in_loop_TOP_LOOP37832_U0_l2_adjustments_d1),
    .l2_adjustments_q1(48'd0),
    .l2_adjustments_we1(dataflow_in_loop_TOP_LOOP37832_U0_l2_adjustments_we1),
    .ap_start(dataflow_in_loop_TOP_LOOP37832_U0_ap_start),
    .in_data_empty_n(1'b0),
    .in_data_read(dataflow_in_loop_TOP_LOOP37832_U0_in_data_read),
    .out_data_full_n(out_data_full_n),
    .out_data_write(dataflow_in_loop_TOP_LOOP37832_U0_out_data_write),
    .ap_done(dataflow_in_loop_TOP_LOOP37832_U0_ap_done),
    .ap_ready(dataflow_in_loop_TOP_LOOP37832_U0_ap_ready),
    .ap_idle(dataflow_in_loop_TOP_LOOP37832_U0_ap_idle),
    .ap_continue(dataflow_in_loop_TOP_LOOP37832_U0_ap_continue)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        loop_dataflow_input_count <= 19'd0;
    end else begin
        if ((~(loop_dataflow_input_count == bound_minus_1) & (ap_start == 1'b1) & (dataflow_in_loop_TOP_LOOP37832_U0_ap_ready == 1'b1))) begin
            loop_dataflow_input_count <= (loop_dataflow_input_count + 19'd1);
        end else if (((loop_dataflow_input_count == bound_minus_1) & (ap_start == 1'b1) & (dataflow_in_loop_TOP_LOOP37832_U0_ap_ready == 1'b1))) begin
            loop_dataflow_input_count <= 19'd0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        loop_dataflow_output_count <= 19'd0;
    end else begin
        if ((~(loop_dataflow_output_count == bound_minus_1) & (dataflow_in_loop_TOP_LOOP37832_U0_ap_continue == 1'b1) & (dataflow_in_loop_TOP_LOOP37832_U0_ap_done == 1'b1))) begin
            loop_dataflow_output_count <= (loop_dataflow_output_count + 19'd1);
        end else if (((loop_dataflow_output_count == bound_minus_1) & (dataflow_in_loop_TOP_LOOP37832_U0_ap_continue == 1'b1) & (dataflow_in_loop_TOP_LOOP37832_U0_ap_done == 1'b1))) begin
            loop_dataflow_output_count <= 19'd0;
        end
    end
end

always @ (*) begin
    if (((loop_dataflow_output_count == bound_minus_1) & (dataflow_in_loop_TOP_LOOP37832_U0_ap_done == 1'b1))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = 1'b0;
    end
end

always @ (*) begin
    if (((loop_dataflow_output_count == 19'd0) & (ap_start == 1'b0) & (dataflow_in_loop_TOP_LOOP37832_U0_ap_idle == 1'b1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((loop_dataflow_input_count == bound_minus_1) & (ap_start == 1'b1) & (dataflow_in_loop_TOP_LOOP37832_U0_ap_ready == 1'b1))) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((~(loop_dataflow_output_count == bound_minus_1) | (ap_continue == 1'b1))) begin
        dataflow_in_loop_TOP_LOOP37832_U0_ap_continue = 1'b1;
    end else begin
        dataflow_in_loop_TOP_LOOP37832_U0_ap_continue = 1'b0;
    end
end

assign ap_sync_continue = ap_continue;

assign ap_sync_done = dataflow_in_loop_TOP_LOOP37832_U0_ap_done;

assign ap_sync_ready = dataflow_in_loop_TOP_LOOP37832_U0_ap_ready;

assign bound_minus_1 = (19'd401408 - 19'd1);

assign dataflow_in_loop_TOP_LOOP37832_U0_ap_start = ap_start;

assign dataflow_in_loop_TOP_LOOP37832_U0_in_data_full_n = in_data_empty_n;

assign dataflow_in_loop_TOP_LOOP37832_U0_in_data_write = 1'b0;

assign dataflow_in_loop_TOP_LOOP37832_U0_start_full_n = 1'b1;

assign dataflow_in_loop_TOP_LOOP37832_U0_start_write = 1'b0;

assign in_data_address0 = dataflow_in_loop_TOP_LOOP37832_U0_in_data_address0;

assign in_data_address1 = 14'd0;

assign in_data_ce0 = dataflow_in_loop_TOP_LOOP37832_U0_in_data_ce0;

assign in_data_ce1 = 1'b0;

assign in_data_d0 = 64'd0;

assign in_data_d1 = 64'd0;

assign in_data_read = dataflow_in_loop_TOP_LOOP37832_U0_in_data_write;

assign in_data_we0 = 1'b0;

assign in_data_we1 = 1'b0;

assign l1_adjustments_address0 = dataflow_in_loop_TOP_LOOP37832_U0_l1_adjustments_address0;

assign l1_adjustments_address1 = 7'd0;

assign l1_adjustments_ce0 = dataflow_in_loop_TOP_LOOP37832_U0_l1_adjustments_ce0;

assign l1_adjustments_ce1 = 1'b0;

assign l1_adjustments_d0 = 48'd0;

assign l1_adjustments_d1 = 48'd0;

assign l1_adjustments_we0 = 1'b0;

assign l1_adjustments_we1 = 1'b0;

assign l1_filter_data_address0 = dataflow_in_loop_TOP_LOOP37832_U0_l1_filter_data_address0;

assign l1_filter_data_address1 = 15'd0;

assign l1_filter_data_ce0 = dataflow_in_loop_TOP_LOOP37832_U0_l1_filter_data_ce0;

assign l1_filter_data_ce1 = 1'b0;

assign l1_filter_data_d0 = 16'd0;

assign l1_filter_data_d1 = 16'd0;

assign l1_filter_data_we0 = 1'b0;

assign l1_filter_data_we1 = 1'b0;

assign l2_adjustments_address0 = dataflow_in_loop_TOP_LOOP37832_U0_l2_adjustments_address0;

assign l2_adjustments_address1 = 4'd0;

assign l2_adjustments_ce0 = dataflow_in_loop_TOP_LOOP37832_U0_l2_adjustments_ce0;

assign l2_adjustments_ce1 = 1'b0;

assign l2_adjustments_d0 = 48'd0;

assign l2_adjustments_d1 = 48'd0;

assign l2_adjustments_we0 = 1'b0;

assign l2_adjustments_we1 = 1'b0;

assign l2_filter_data_address0 = dataflow_in_loop_TOP_LOOP37832_U0_l2_filter_data_address0;

assign l2_filter_data_address1 = 11'd0;

assign l2_filter_data_ce0 = dataflow_in_loop_TOP_LOOP37832_U0_l2_filter_data_ce0;

assign l2_filter_data_ce1 = 1'b0;

assign l2_filter_data_d0 = 16'd0;

assign l2_filter_data_d1 = 16'd0;

assign l2_filter_data_we0 = 1'b0;

assign l2_filter_data_we1 = 1'b0;

assign out_data_address0 = 14'd0;

assign out_data_address1 = dataflow_in_loop_TOP_LOOP37832_U0_out_data_address1;

assign out_data_ce0 = 1'b0;

assign out_data_ce1 = dataflow_in_loop_TOP_LOOP37832_U0_out_data_ce1;

assign out_data_d0 = 64'd0;

assign out_data_d1 = dataflow_in_loop_TOP_LOOP37832_U0_out_data_d1;

assign out_data_we0 = 1'b0;

assign out_data_we1 = dataflow_in_loop_TOP_LOOP37832_U0_out_data_we1;

assign out_data_write = dataflow_in_loop_TOP_LOOP37832_U0_out_data_write;

endmodule //td_fused_top_tdf4_111
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf4_accum_1 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        accum_in_0_address0,
        accum_in_0_ce0,
        accum_in_0_q0,
        accum_in_0_address1,
        accum_in_0_ce1,
        accum_in_0_q1,
        accum_out_address0,
        accum_out_ce0,
        accum_out_we0,
        accum_out_d0,
        accum_out_address1,
        accum_out_ce1,
        accum_out_we1,
        accum_out_d1
);

parameter    ap_ST_fsm_state1 = 8'd1;
parameter    ap_ST_fsm_pp0_stage0 = 8'd2;
parameter    ap_ST_fsm_pp0_stage1 = 8'd4;
parameter    ap_ST_fsm_pp0_stage2 = 8'd8;
parameter    ap_ST_fsm_pp0_stage3 = 8'd16;
parameter    ap_ST_fsm_state12 = 8'd32;
parameter    ap_ST_fsm_state13 = 8'd64;
parameter    ap_ST_fsm_state14 = 8'd128;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [7:0] accum_in_0_address0;
output   accum_in_0_ce0;
input  [15:0] accum_in_0_q0;
output  [7:0] accum_in_0_address1;
output   accum_in_0_ce1;
input  [15:0] accum_in_0_q1;
output  [2:0] accum_out_address0;
output   accum_out_ce0;
output   accum_out_we0;
output  [15:0] accum_out_d0;
output  [2:0] accum_out_address1;
output   accum_out_ce1;
output   accum_out_we1;
output  [15:0] accum_out_d1;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg[7:0] accum_in_0_address0;
reg accum_in_0_ce0;
reg[7:0] accum_in_0_address1;
reg accum_in_0_ce1;
reg accum_out_ce0;
reg accum_out_we0;
reg accum_out_ce1;
reg accum_out_we1;

reg    ap_done_reg;
  reg   [7:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg   [7:0] x_reg_168;
reg   [15:0] psum_7_08_reg_180;
reg   [15:0] psum_6_07_reg_192;
reg   [15:0] psum_5_06_reg_204;
reg   [15:0] psum_4_05_reg_216;
reg   [15:0] psum_3_04_reg_228;
reg   [15:0] psum_2_03_reg_240;
reg   [15:0] psum_1_02_reg_252;
reg   [15:0] psum_0_01_reg_264;
wire   [0:0] icmp_ln132_fu_321_p2;
reg   [0:0] icmp_ln132_reg_492;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state6_pp0_stage0_iter1;
wire    ap_block_state10_pp0_stage0_iter2;
wire    ap_block_pp0_stage0_11001;
reg   [0:0] icmp_ln132_reg_492_pp0_iter1_reg;
reg   [0:0] icmp_ln132_reg_492_pp0_iter2_reg;
reg   [15:0] accum_in_0_load_reg_506;
wire    ap_CS_fsm_pp0_stage1;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_state3_pp0_stage1_iter0;
wire    ap_block_state7_pp0_stage1_iter1;
wire    ap_block_state11_pp0_stage1_iter2;
wire    ap_block_pp0_stage1_11001;
reg   [15:0] accum_in_0_load_36_reg_511;
reg   [15:0] accum_in_0_load_37_reg_526;
wire    ap_CS_fsm_pp0_stage2;
wire    ap_block_state4_pp0_stage2_iter0;
wire    ap_block_state8_pp0_stage2_iter1;
wire    ap_block_pp0_stage2_11001;
reg   [15:0] accum_in_0_load_38_reg_531;
wire   [7:0] add_ln132_fu_387_p2;
reg   [7:0] add_ln132_reg_546;
wire    ap_CS_fsm_pp0_stage3;
wire    ap_block_state5_pp0_stage3_iter0;
wire    ap_block_state9_pp0_stage3_iter1;
wire    ap_block_pp0_stage3_11001;
reg   [15:0] accum_in_0_load_39_reg_551;
reg   [15:0] accum_in_0_load_40_reg_556;
reg   [15:0] accum_in_0_load_41_reg_571;
reg    ap_enable_reg_pp0_iter1;
reg   [15:0] accum_in_0_load_42_reg_576;
wire   [15:0] grp_fu_305_p2;
wire   [15:0] grp_fu_310_p2;
reg    ap_enable_reg_pp0_iter2;
wire   [3:0] add_ln140_fu_432_p2;
wire    ap_CS_fsm_state13;
wire   [0:0] tmp_fu_415_p3;
reg    ap_block_state1;
wire    ap_block_pp0_stage2_subdone;
reg    ap_condition_pp0_exit_iter0_state4;
wire    ap_block_pp0_stage3_subdone;
wire    ap_block_pp0_stage1_subdone;
reg   [7:0] ap_phi_mux_x_phi_fu_172_p4;
wire    ap_block_pp0_stage0;
wire   [15:0] ap_phi_mux_psum_7_08_phi_fu_184_p4;
wire    ap_block_pp0_stage1;
wire   [15:0] ap_phi_mux_psum_6_07_phi_fu_196_p4;
wire   [15:0] ap_phi_mux_psum_5_06_phi_fu_208_p4;
wire   [15:0] ap_phi_mux_psum_4_05_phi_fu_220_p4;
wire   [15:0] ap_phi_mux_psum_3_04_phi_fu_232_p4;
wire    ap_block_pp0_stage3;
wire   [15:0] ap_phi_mux_psum_2_03_phi_fu_244_p4;
wire    ap_block_pp0_stage2;
reg   [3:0] q_reg_276;
wire    ap_CS_fsm_state12;
reg   [15:0] ap_phi_mux_phi_ln152_phi_fu_290_p8;
wire   [2:0] trunc_ln140_fu_428_p1;
wire   [63:0] zext_ln132_fu_327_p1;
wire   [63:0] zext_ln136_fu_338_p1;
wire   [63:0] zext_ln136_7_fu_349_p1;
wire   [63:0] zext_ln136_8_fu_360_p1;
wire   [63:0] zext_ln136_9_fu_371_p1;
wire   [63:0] zext_ln136_10_fu_382_p1;
wire   [63:0] zext_ln136_11_fu_399_p1;
wire   [63:0] zext_ln136_12_fu_410_p1;
wire   [63:0] zext_ln140_fu_423_p1;
wire   [63:0] zext_ln140_2_fu_444_p1;
reg   [15:0] grp_fu_305_p0;
reg   [15:0] grp_fu_305_p1;
reg   [15:0] grp_fu_310_p0;
reg   [15:0] grp_fu_310_p1;
wire   [7:0] or_ln136_fu_332_p2;
wire   [7:0] or_ln136_7_fu_343_p2;
wire   [7:0] or_ln136_8_fu_354_p2;
wire   [7:0] or_ln136_9_fu_365_p2;
wire   [7:0] or_ln136_10_fu_376_p2;
wire   [7:0] or_ln136_11_fu_393_p2;
wire   [7:0] or_ln136_12_fu_404_p2;
wire   [2:0] or_ln140_fu_438_p2;
wire   [0:0] icmp_ln152_fu_449_p2;
wire   [0:0] icmp_ln152_3_fu_463_p2;
wire   [15:0] select_ln152_fu_455_p3;
wire   [0:0] icmp_ln152_4_fu_477_p2;
wire   [15:0] select_ln152_3_fu_469_p3;
wire    ap_CS_fsm_state14;
reg   [7:0] ap_NS_fsm;
wire    ap_block_pp0_stage0_subdone;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
reg    ap_condition_514;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 8'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
end

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U220(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(grp_fu_305_p0),
    .din1(grp_fu_305_p1),
    .dout(grp_fu_305_p2)
);

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U221(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(grp_fu_310_p0),
    .din1(grp_fu_310_p1),
    .dout(grp_fu_310_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state14)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage2_subdone) & (1'b1 == ap_condition_pp0_exit_iter0_state4) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage3_subdone) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b0)) | ((1'b0 == ap_block_pp0_stage3_subdone) & (1'b1 == ap_CS_fsm_pp0_stage3)))) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end else if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter2 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state12)) begin
        q_reg_276 <= 4'd0;
    end else if (((tmp_fu_415_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state13))) begin
        q_reg_276 <= add_ln140_fu_432_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln132_reg_492 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        x_reg_168 <= add_ln132_reg_546;
    end else if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        x_reg_168 <= 8'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage1_11001) & (icmp_ln132_reg_492 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
        accum_in_0_load_36_reg_511 <= accum_in_0_q0;
        accum_in_0_load_reg_506 <= accum_in_0_q1;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2_11001) & (icmp_ln132_reg_492 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
        accum_in_0_load_37_reg_526 <= accum_in_0_q1;
        accum_in_0_load_38_reg_531 <= accum_in_0_q0;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage3_11001) & (icmp_ln132_reg_492 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
        accum_in_0_load_39_reg_551 <= accum_in_0_q1;
        accum_in_0_load_40_reg_556 <= accum_in_0_q0;
        add_ln132_reg_546 <= add_ln132_fu_387_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln132_reg_492 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        accum_in_0_load_41_reg_571 <= accum_in_0_q1;
        accum_in_0_load_42_reg_576 <= accum_in_0_q0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln132_reg_492 <= icmp_ln132_fu_321_p2;
        icmp_ln132_reg_492_pp0_iter1_reg <= icmp_ln132_reg_492;
        icmp_ln132_reg_492_pp0_iter2_reg <= icmp_ln132_reg_492_pp0_iter1_reg;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln132_reg_492_pp0_iter1_reg == 1'd1) & (1'b0 == ap_block_pp0_stage2_11001) & (1'b1 == ap_CS_fsm_pp0_stage2) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        psum_0_01_reg_264 <= grp_fu_305_p2;
        psum_1_02_reg_252 <= grp_fu_310_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln132_reg_492_pp0_iter1_reg == 1'd1) & (1'b0 == ap_block_pp0_stage3_11001) & (1'b1 == ap_CS_fsm_pp0_stage3) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        psum_2_03_reg_240 <= grp_fu_305_p2;
        psum_3_04_reg_228 <= grp_fu_310_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln132_reg_492_pp0_iter1_reg == 1'd1) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        psum_4_05_reg_216 <= grp_fu_305_p2;
        psum_5_06_reg_204 <= grp_fu_310_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln132_reg_492_pp0_iter2_reg == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        psum_6_07_reg_192 <= grp_fu_305_p2;
        psum_7_08_reg_180 <= grp_fu_310_p2;
    end
end

always @ (*) begin
    if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
        if (((1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            accum_in_0_address0 = zext_ln136_12_fu_410_p1;
        end else if (((1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            accum_in_0_address0 = zext_ln136_10_fu_382_p1;
        end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            accum_in_0_address0 = zext_ln136_8_fu_360_p1;
        end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            accum_in_0_address0 = zext_ln136_fu_338_p1;
        end else begin
            accum_in_0_address0 = 'bx;
        end
    end else begin
        accum_in_0_address0 = 'bx;
    end
end

always @ (*) begin
    if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
        if (((1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            accum_in_0_address1 = zext_ln136_11_fu_399_p1;
        end else if (((1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            accum_in_0_address1 = zext_ln136_9_fu_371_p1;
        end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            accum_in_0_address1 = zext_ln136_7_fu_349_p1;
        end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            accum_in_0_address1 = zext_ln132_fu_327_p1;
        end else begin
            accum_in_0_address1 = 'bx;
        end
    end else begin
        accum_in_0_address1 = 'bx;
    end
end

always @ (*) begin
    if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage3_11001) & (1'b1 == ap_CS_fsm_pp0_stage3)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2_11001) & (1'b1 == ap_CS_fsm_pp0_stage2)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1)))) begin
        accum_in_0_ce0 = 1'b1;
    end else begin
        accum_in_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage3_11001) & (1'b1 == ap_CS_fsm_pp0_stage3)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2_11001) & (1'b1 == ap_CS_fsm_pp0_stage2)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1)))) begin
        accum_in_0_ce1 = 1'b1;
    end else begin
        accum_in_0_ce1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state13)) begin
        accum_out_ce0 = 1'b1;
    end else begin
        accum_out_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state13)) begin
        accum_out_ce1 = 1'b1;
    end else begin
        accum_out_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((tmp_fu_415_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state13))) begin
        accum_out_we0 = 1'b1;
    end else begin
        accum_out_we0 = 1'b0;
    end
end

always @ (*) begin
    if (((tmp_fu_415_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state13))) begin
        accum_out_we1 = 1'b1;
    end else begin
        accum_out_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((icmp_ln132_reg_492 == 1'd0)) begin
        ap_condition_pp0_exit_iter0_state4 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state4 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state14)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((tmp_fu_415_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state13))) begin
        if ((trunc_ln140_fu_428_p1 == 3'd0)) begin
            ap_phi_mux_phi_ln152_phi_fu_290_p8 = psum_0_01_reg_264;
        end else if ((1'b1 == ap_condition_514)) begin
            ap_phi_mux_phi_ln152_phi_fu_290_p8 = psum_6_07_reg_192;
        end else if ((trunc_ln140_fu_428_p1 == 3'd4)) begin
            ap_phi_mux_phi_ln152_phi_fu_290_p8 = psum_4_05_reg_216;
        end else if ((trunc_ln140_fu_428_p1 == 3'd2)) begin
            ap_phi_mux_phi_ln152_phi_fu_290_p8 = psum_2_03_reg_240;
        end else begin
            ap_phi_mux_phi_ln152_phi_fu_290_p8 = 'bx;
        end
    end else begin
        ap_phi_mux_phi_ln152_phi_fu_290_p8 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0) & (icmp_ln132_reg_492 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_x_phi_fu_172_p4 = add_ln132_reg_546;
    end else begin
        ap_phi_mux_x_phi_fu_172_p4 = x_reg_168;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state14)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_305_p0 = ap_phi_mux_psum_6_07_phi_fu_196_p4;
    end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_305_p0 = ap_phi_mux_psum_4_05_phi_fu_220_p4;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
        grp_fu_305_p0 = ap_phi_mux_psum_2_03_phi_fu_244_p4;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
        grp_fu_305_p0 = grp_fu_305_p2;
    end else begin
        grp_fu_305_p0 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_305_p1 = accum_in_0_load_41_reg_571;
    end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_305_p1 = accum_in_0_load_39_reg_551;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
        grp_fu_305_p1 = accum_in_0_load_37_reg_526;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
        grp_fu_305_p1 = accum_in_0_load_reg_506;
    end else begin
        grp_fu_305_p1 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_310_p0 = ap_phi_mux_psum_7_08_phi_fu_184_p4;
    end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_310_p0 = ap_phi_mux_psum_5_06_phi_fu_208_p4;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
        grp_fu_310_p0 = ap_phi_mux_psum_3_04_phi_fu_232_p4;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
        grp_fu_310_p0 = grp_fu_310_p2;
    end else begin
        grp_fu_310_p0 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_310_p1 = accum_in_0_load_42_reg_576;
    end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_310_p1 = accum_in_0_load_40_reg_556;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
        grp_fu_310_p1 = accum_in_0_load_38_reg_531;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
        grp_fu_310_p1 = accum_in_0_load_36_reg_511;
    end else begin
        grp_fu_310_p1 = 'bx;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_pp0_stage1 : begin
            if ((~((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter2 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0)) & (1'b0 == ap_block_pp0_stage1_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage2;
            end else if (((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter2 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
                ap_NS_fsm = ap_ST_fsm_state12;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end
        end
        ap_ST_fsm_pp0_stage2 : begin
            if ((~((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2_subdone) & (icmp_ln132_reg_492 == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b0)) & (1'b0 == ap_block_pp0_stage2_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage3;
            end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2_subdone) & (icmp_ln132_reg_492 == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
                ap_NS_fsm = ap_ST_fsm_state12;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage2;
            end
        end
        ap_ST_fsm_pp0_stage3 : begin
            if ((1'b0 == ap_block_pp0_stage3_subdone)) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage3;
            end
        end
        ap_ST_fsm_state12 : begin
            ap_NS_fsm = ap_ST_fsm_state13;
        end
        ap_ST_fsm_state13 : begin
            if (((tmp_fu_415_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state13))) begin
                ap_NS_fsm = ap_ST_fsm_state13;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state14;
            end
        end
        ap_ST_fsm_state14 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign accum_out_address0 = zext_ln140_2_fu_444_p1;

assign accum_out_address1 = zext_ln140_fu_423_p1;

assign accum_out_d0 = ((icmp_ln152_4_fu_477_p2[0:0] == 1'b1) ? psum_5_06_reg_204 : select_ln152_3_fu_469_p3);

assign accum_out_d1 = ap_phi_mux_phi_ln152_phi_fu_290_p8;

assign add_ln132_fu_387_p2 = (x_reg_168 + 8'd8);

assign add_ln140_fu_432_p2 = (q_reg_276 + 4'd2);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_pp0_stage1 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_pp0_stage2 = ap_CS_fsm[32'd3];

assign ap_CS_fsm_pp0_stage3 = ap_CS_fsm[32'd4];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state12 = ap_CS_fsm[32'd5];

assign ap_CS_fsm_state13 = ap_CS_fsm[32'd6];

assign ap_CS_fsm_state14 = ap_CS_fsm[32'd7];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1_subdone = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage2 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage2_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage2_subdone = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage3 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage3_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage3_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((ap_done_reg == 1'b1) | (ap_start == 1'b0));
end

assign ap_block_state10_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state11_pp0_stage1_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage1_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage2_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage3_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage1_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage2_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state9_pp0_stage3_iter1 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_condition_514 = (~(trunc_ln140_fu_428_p1 == 3'd0) & ~(trunc_ln140_fu_428_p1 == 3'd4) & ~(trunc_ln140_fu_428_p1 == 3'd2));
end

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign ap_phi_mux_psum_2_03_phi_fu_244_p4 = grp_fu_305_p2;

assign ap_phi_mux_psum_3_04_phi_fu_232_p4 = grp_fu_310_p2;

assign ap_phi_mux_psum_4_05_phi_fu_220_p4 = grp_fu_305_p2;

assign ap_phi_mux_psum_5_06_phi_fu_208_p4 = grp_fu_310_p2;

assign ap_phi_mux_psum_6_07_phi_fu_196_p4 = grp_fu_305_p2;

assign ap_phi_mux_psum_7_08_phi_fu_184_p4 = grp_fu_310_p2;

assign icmp_ln132_fu_321_p2 = ((ap_phi_mux_x_phi_fu_172_p4 < 8'd144) ? 1'b1 : 1'b0);

assign icmp_ln152_3_fu_463_p2 = ((or_ln140_fu_438_p2 == 3'd3) ? 1'b1 : 1'b0);

assign icmp_ln152_4_fu_477_p2 = ((or_ln140_fu_438_p2 == 3'd5) ? 1'b1 : 1'b0);

assign icmp_ln152_fu_449_p2 = ((or_ln140_fu_438_p2 == 3'd1) ? 1'b1 : 1'b0);

assign or_ln136_10_fu_376_p2 = (x_reg_168 | 8'd5);

assign or_ln136_11_fu_393_p2 = (x_reg_168 | 8'd6);

assign or_ln136_12_fu_404_p2 = (x_reg_168 | 8'd7);

assign or_ln136_7_fu_343_p2 = (x_reg_168 | 8'd2);

assign or_ln136_8_fu_354_p2 = (x_reg_168 | 8'd3);

assign or_ln136_9_fu_365_p2 = (x_reg_168 | 8'd4);

assign or_ln136_fu_332_p2 = (ap_phi_mux_x_phi_fu_172_p4 | 8'd1);

assign or_ln140_fu_438_p2 = (trunc_ln140_fu_428_p1 | 3'd1);

assign select_ln152_3_fu_469_p3 = ((icmp_ln152_3_fu_463_p2[0:0] == 1'b1) ? psum_3_04_reg_228 : select_ln152_fu_455_p3);

assign select_ln152_fu_455_p3 = ((icmp_ln152_fu_449_p2[0:0] == 1'b1) ? psum_1_02_reg_252 : psum_7_08_reg_180);

assign tmp_fu_415_p3 = q_reg_276[32'd3];

assign trunc_ln140_fu_428_p1 = q_reg_276[2:0];

assign zext_ln132_fu_327_p1 = ap_phi_mux_x_phi_fu_172_p4;

assign zext_ln136_10_fu_382_p1 = or_ln136_10_fu_376_p2;

assign zext_ln136_11_fu_399_p1 = or_ln136_11_fu_393_p2;

assign zext_ln136_12_fu_410_p1 = or_ln136_12_fu_404_p2;

assign zext_ln136_7_fu_349_p1 = or_ln136_7_fu_343_p2;

assign zext_ln136_8_fu_360_p1 = or_ln136_8_fu_354_p2;

assign zext_ln136_9_fu_371_p1 = or_ln136_9_fu_365_p2;

assign zext_ln136_fu_338_p1 = or_ln136_fu_332_p2;

assign zext_ln140_2_fu_444_p1 = or_ln140_fu_438_p2;

assign zext_ln140_fu_423_p1 = q_reg_276;

endmodule //td_fused_top_tdf4_accum_1
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf4_accum_2 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        accum_in_12,
        accum_in_12_ap_vld,
        accum_in_address0,
        accum_in_ce0,
        accum_in_q0
);

parameter    ap_ST_fsm_state1 = 7'd1;
parameter    ap_ST_fsm_state2 = 7'd2;
parameter    ap_ST_fsm_state3 = 7'd4;
parameter    ap_ST_fsm_state4 = 7'd8;
parameter    ap_ST_fsm_state5 = 7'd16;
parameter    ap_ST_fsm_state6 = 7'd32;
parameter    ap_ST_fsm_state7 = 7'd64;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [15:0] accum_in_12;
output   accum_in_12_ap_vld;
output  [2:0] accum_in_address0;
output   accum_in_ce0;
input  [15:0] accum_in_q0;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg[15:0] accum_in_12;
reg accum_in_12_ap_vld;
reg accum_in_ce0;

reg    ap_done_reg;
  reg   [6:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
wire   [3:0] add_ln164_fu_74_p2;
reg   [3:0] add_ln164_reg_91;
wire    ap_CS_fsm_state2;
wire   [0:0] icmp_ln164_fu_85_p2;
wire    ap_CS_fsm_state3;
wire   [15:0] grp_fu_68_p2;
wire    ap_CS_fsm_state7;
reg   [3:0] i_1_1_reg_44;
reg    ap_block_state1;
reg   [15:0] sum_01_reg_55;
wire   [63:0] zext_ln164_fu_80_p1;
reg   [15:0] accum_in_12_preg;
reg   [6:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 7'd1;
#0 accum_in_12_preg = 16'd0;
end

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U224(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(sum_01_reg_55),
    .din1(accum_in_q0),
    .dout(grp_fu_68_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        accum_in_12_preg <= 16'd0;
    end else begin
        if (((icmp_ln164_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
            accum_in_12_preg <= sum_01_reg_55;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if (((icmp_ln164_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        i_1_1_reg_44 <= 4'd0;
    end else if ((1'b1 == ap_CS_fsm_state7)) begin
        i_1_1_reg_44 <= add_ln164_reg_91;
    end
end

always @ (posedge ap_clk) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        sum_01_reg_55 <= 16'd0;
    end else if ((1'b1 == ap_CS_fsm_state7)) begin
        sum_01_reg_55 <= grp_fu_68_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        add_ln164_reg_91 <= add_ln164_fu_74_p2;
    end
end

always @ (*) begin
    if (((icmp_ln164_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        accum_in_12 = sum_01_reg_55;
    end else begin
        accum_in_12 = accum_in_12_preg;
    end
end

always @ (*) begin
    if (((icmp_ln164_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        accum_in_12_ap_vld = 1'b1;
    end else begin
        accum_in_12_ap_vld = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        accum_in_ce0 = 1'b1;
    end else begin
        accum_in_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln164_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln164_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_state2 : begin
            if (((icmp_ln164_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end
        end
        ap_ST_fsm_state3 : begin
            ap_NS_fsm = ap_ST_fsm_state4;
        end
        ap_ST_fsm_state4 : begin
            ap_NS_fsm = ap_ST_fsm_state5;
        end
        ap_ST_fsm_state5 : begin
            ap_NS_fsm = ap_ST_fsm_state6;
        end
        ap_ST_fsm_state6 : begin
            ap_NS_fsm = ap_ST_fsm_state7;
        end
        ap_ST_fsm_state7 : begin
            ap_NS_fsm = ap_ST_fsm_state2;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign accum_in_address0 = zext_ln164_fu_80_p1;

assign add_ln164_fu_74_p2 = (i_1_1_reg_44 + 4'd1);

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state7 = ap_CS_fsm[32'd6];

always @ (*) begin
    ap_block_state1 = ((ap_done_reg == 1'b1) | (ap_start == 1'b0));
end

assign icmp_ln164_fu_85_p2 = ((i_1_1_reg_44 == 4'd8) ? 1'b1 : 1'b0);

assign zext_ln164_fu_80_p1 = i_1_1_reg_44;

endmodule //td_fused_top_tdf4_accum_2
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_tdf4_adjustments_ram (addr0, ce0, q0, addr1, ce1, d1, we1,  clk);

parameter DWIDTH = 48;
parameter AWIDTH = 7;
parameter MEM_SIZE = 128;

input[AWIDTH-1:0] addr0;
input ce0;
output wire[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
input clk;

 reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];
wire [AWIDTH-1:0] addr0_t0; 
reg [AWIDTH-1:0] addr0_t1; 
reg [DWIDTH-1:0] q0_t0;
reg [DWIDTH-1:0] q0_t1;
wire [AWIDTH-1:0] addr1_t0; 
reg [AWIDTH-1:0] addr1_t1; 
wire [DWIDTH-1:0] d1_t0; 
wire we1_t0; 
reg [DWIDTH-1:0] d1_t1; 
reg we1_t1; 


assign addr0_t0 = addr0;
assign q0 = q0_t1;
assign addr1_t0 = addr1;
assign d1_t0 = d1;
assign we1_t0 = we1;

always @(posedge clk)  
begin
    if (ce0) 
    begin
        addr0_t1 <= addr0_t0; 
        q0_t1 <= q0_t0;
    end
    if (ce1) 
    begin
        addr1_t1 <= addr1_t0; 
        d1_t1 <= d1_t0;
        we1_t1 <= we1_t0;
    end
end


always @(posedge clk)  
begin 
    if (ce0) begin
        q0_t0 <= ram[addr0_t1];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1_t1) 
            ram[addr1_t1] <= d1_t1; 
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_tdf4_adjustments(
    reset,
    clk,
    address0,
    ce0,
    q0,
    address1,
    ce1,
    we1,
    d1);

parameter DataWidth = 32'd48;
parameter AddressRange = 32'd128;
parameter AddressWidth = 32'd7;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;



td_fused_top_tdf4_adjustments_ram td_fused_top_tdf4_adjustments_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 )
);

endmodule

// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf4_adjust (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        sums_read,
        adjustments_address0,
        adjustments_ce0,
        adjustments_q0,
        indices_23_dout,
        indices_23_empty_n,
        indices_23_read,
        indices_23_out_din,
        indices_23_out_full_n,
        indices_23_out_write,
        ap_return
);

parameter    ap_ST_fsm_state1 = 17'd1;
parameter    ap_ST_fsm_state2 = 17'd2;
parameter    ap_ST_fsm_state3 = 17'd4;
parameter    ap_ST_fsm_state4 = 17'd8;
parameter    ap_ST_fsm_state5 = 17'd16;
parameter    ap_ST_fsm_state6 = 17'd32;
parameter    ap_ST_fsm_state7 = 17'd64;
parameter    ap_ST_fsm_state8 = 17'd128;
parameter    ap_ST_fsm_state9 = 17'd256;
parameter    ap_ST_fsm_state10 = 17'd512;
parameter    ap_ST_fsm_state11 = 17'd1024;
parameter    ap_ST_fsm_state12 = 17'd2048;
parameter    ap_ST_fsm_state13 = 17'd4096;
parameter    ap_ST_fsm_state14 = 17'd8192;
parameter    ap_ST_fsm_state15 = 17'd16384;
parameter    ap_ST_fsm_state16 = 17'd32768;
parameter    ap_ST_fsm_state17 = 17'd65536;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
input  [15:0] sums_read;
output  [6:0] adjustments_address0;
output   adjustments_ce0;
input  [47:0] adjustments_q0;
input  [10:0] indices_23_dout;
input   indices_23_empty_n;
output   indices_23_read;
output  [10:0] indices_23_out_din;
input   indices_23_out_full_n;
output   indices_23_out_write;
output  [15:0] ap_return;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg adjustments_ce0;
reg indices_23_read;
reg indices_23_out_write;

reg    ap_done_reg;
  reg   [16:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    indices_23_blk_n;
reg    indices_23_out_blk_n;
wire    ap_CS_fsm_state4;
reg   [15:0] tmp_53_i_i_reg_183;
reg   [15:0] tmp_54_i_i_reg_188;
wire   [15:0] grp_fu_93_p2;
reg   [15:0] sub_i_i_i_reg_193;
wire    ap_CS_fsm_state8;
wire    ap_CS_fsm_state9;
wire   [15:0] grp_fu_98_p2;
reg   [15:0] mul_i_i_i_reg_203;
wire    ap_CS_fsm_state12;
wire    ap_CS_fsm_state13;
wire   [63:0] zext_ln220_fu_106_p1;
reg    ap_block_state1;
wire    ap_CS_fsm_state2;
wire    ap_CS_fsm_state3;
wire   [15:0] grp_fu_89_p1;
wire   [15:0] grp_fu_93_p1;
wire   [15:0] grp_fu_98_p1;
wire   [6:0] trunc_ln251_fu_102_p1;
wire   [15:0] trunc_ln220_fu_111_p1;
wire   [15:0] grp_fu_89_p2;
wire    ap_CS_fsm_state17;
wire   [15:0] bitcast_ln648_fu_148_p1;
wire   [0:0] tmp_fu_152_p3;
reg   [16:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 17'd1;
end

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U228(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(mul_i_i_i_reg_203),
    .din1(grp_fu_89_p1),
    .dout(grp_fu_89_p2)
);

td_fused_top_hsub_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hsub_16ns_16ns_16_5_full_dsp_1_U229(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(sums_read),
    .din1(grp_fu_93_p1),
    .dout(grp_fu_93_p2)
);

td_fused_top_hmul_16ns_16ns_16_4_max_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hmul_16ns_16ns_16_4_max_dsp_1_U230(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(sub_i_i_i_reg_193),
    .din1(grp_fu_98_p1),
    .dout(grp_fu_98_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state17)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state12)) begin
        mul_i_i_i_reg_203 <= grp_fu_98_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state8)) begin
        sub_i_i_i_reg_193 <= grp_fu_93_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        tmp_53_i_i_reg_183 <= {{adjustments_q0[31:16]}};
        tmp_54_i_i_reg_188 <= {{adjustments_q0[47:32]}};
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state2) | (~((indices_23_out_full_n == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1)))) begin
        adjustments_ce0 = 1'b1;
    end else begin
        adjustments_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state17)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state17)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_23_blk_n = indices_23_empty_n;
    end else begin
        indices_23_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_23_out_blk_n = indices_23_out_full_n;
    end else begin
        indices_23_out_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((indices_23_out_full_n == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_23_out_write = 1'b1;
    end else begin
        indices_23_out_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((indices_23_out_full_n == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_23_read = 1'b1;
    end else begin
        indices_23_read = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((indices_23_out_full_n == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_state2 : begin
            ap_NS_fsm = ap_ST_fsm_state3;
        end
        ap_ST_fsm_state3 : begin
            ap_NS_fsm = ap_ST_fsm_state4;
        end
        ap_ST_fsm_state4 : begin
            ap_NS_fsm = ap_ST_fsm_state5;
        end
        ap_ST_fsm_state5 : begin
            ap_NS_fsm = ap_ST_fsm_state6;
        end
        ap_ST_fsm_state6 : begin
            ap_NS_fsm = ap_ST_fsm_state7;
        end
        ap_ST_fsm_state7 : begin
            ap_NS_fsm = ap_ST_fsm_state8;
        end
        ap_ST_fsm_state8 : begin
            ap_NS_fsm = ap_ST_fsm_state9;
        end
        ap_ST_fsm_state9 : begin
            ap_NS_fsm = ap_ST_fsm_state10;
        end
        ap_ST_fsm_state10 : begin
            ap_NS_fsm = ap_ST_fsm_state11;
        end
        ap_ST_fsm_state11 : begin
            ap_NS_fsm = ap_ST_fsm_state12;
        end
        ap_ST_fsm_state12 : begin
            ap_NS_fsm = ap_ST_fsm_state13;
        end
        ap_ST_fsm_state13 : begin
            ap_NS_fsm = ap_ST_fsm_state14;
        end
        ap_ST_fsm_state14 : begin
            ap_NS_fsm = ap_ST_fsm_state15;
        end
        ap_ST_fsm_state15 : begin
            ap_NS_fsm = ap_ST_fsm_state16;
        end
        ap_ST_fsm_state16 : begin
            ap_NS_fsm = ap_ST_fsm_state17;
        end
        ap_ST_fsm_state17 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign adjustments_address0 = zext_ln220_fu_106_p1;

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state12 = ap_CS_fsm[32'd11];

assign ap_CS_fsm_state13 = ap_CS_fsm[32'd12];

assign ap_CS_fsm_state17 = ap_CS_fsm[32'd16];

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

assign ap_CS_fsm_state8 = ap_CS_fsm[32'd7];

assign ap_CS_fsm_state9 = ap_CS_fsm[32'd8];

always @ (*) begin
    ap_block_state1 = ((indices_23_out_full_n == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0));
end

assign ap_return = ((tmp_fu_152_p3[0:0] == 1'b1) ? 16'd0 : grp_fu_89_p2);

assign bitcast_ln648_fu_148_p1 = grp_fu_89_p2;

assign grp_fu_89_p1 = tmp_54_i_i_reg_188;

assign grp_fu_93_p1 = trunc_ln220_fu_111_p1;

assign grp_fu_98_p1 = tmp_53_i_i_reg_183;

assign indices_23_out_din = indices_23_dout;

assign tmp_fu_152_p3 = bitcast_ln648_fu_148_p1[32'd15];

assign trunc_ln220_fu_111_p1 = adjustments_q0[15:0];

assign trunc_ln251_fu_102_p1 = indices_23_dout[6:0];

assign zext_ln220_fu_106_p1 = trunc_ln251_fu_102_p1;

endmodule //td_fused_top_tdf4_adjust
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf4_dot_product (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        ifmap_vec_address0,
        ifmap_vec_ce0,
        ifmap_vec_q0,
        weight_vecs_0_address0,
        weight_vecs_0_ce0,
        weight_vecs_0_q0,
        products_0_address0,
        products_0_ce0,
        products_0_we0,
        products_0_d0
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state10 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [7:0] ifmap_vec_address0;
output   ifmap_vec_ce0;
input  [15:0] ifmap_vec_q0;
output  [7:0] weight_vecs_0_address0;
output   weight_vecs_0_ce0;
input  [15:0] weight_vecs_0_q0;
output  [7:0] products_0_address0;
output   products_0_ce0;
output   products_0_we0;
output  [15:0] products_0_d0;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg ifmap_vec_ce0;
reg weight_vecs_0_ce0;
reg products_0_ce0;
reg products_0_we0;

reg    ap_done_reg;
  reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg   [7:0] indvar_flatten17_reg_97;
reg   [6:0] indvar_flatten_reg_108;
reg   [1:0] jj_reg_119;
reg   [4:0] ic_reg_131;
reg   [1:0] ii_reg_142;
wire   [7:0] add_ln147_4_fu_157_p2;
wire    ap_CS_fsm_pp0_stage0;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
wire    ap_block_state4_pp0_stage0_iter2;
wire    ap_block_state5_pp0_stage0_iter3;
wire    ap_block_state6_pp0_stage0_iter4;
wire    ap_block_state7_pp0_stage0_iter5;
wire    ap_block_state8_pp0_stage0_iter6;
wire    ap_block_state9_pp0_stage0_iter7;
wire    ap_block_pp0_stage0_11001;
wire   [0:0] icmp_ln147_fu_163_p2;
reg   [0:0] icmp_ln147_reg_408;
reg   [0:0] icmp_ln147_reg_408_pp0_iter1_reg;
reg   [0:0] icmp_ln147_reg_408_pp0_iter2_reg;
reg   [0:0] icmp_ln147_reg_408_pp0_iter3_reg;
reg   [0:0] icmp_ln147_reg_408_pp0_iter4_reg;
reg   [0:0] icmp_ln147_reg_408_pp0_iter5_reg;
reg   [0:0] icmp_ln147_reg_408_pp0_iter6_reg;
wire   [0:0] icmp_ln148_fu_169_p2;
reg   [0:0] icmp_ln148_reg_412;
wire   [0:0] and_ln147_fu_195_p2;
reg   [0:0] and_ln147_reg_419;
wire   [1:0] add_ln148_fu_201_p2;
reg   [1:0] add_ln148_reg_424;
wire   [4:0] select_ln148_fu_213_p3;
reg   [4:0] select_ln148_reg_429;
wire   [1:0] select_ln148_10_fu_221_p3;
reg   [1:0] select_ln148_10_reg_434;
wire   [3:0] trunc_ln150_fu_229_p1;
reg   [3:0] trunc_ln150_reg_440;
reg   [3:0] trunc_ln150_reg_440_pp0_iter1_reg;
reg   [3:0] trunc_ln150_reg_440_pp0_iter2_reg;
reg   [3:0] trunc_ln150_reg_440_pp0_iter3_reg;
reg   [3:0] trunc_ln150_reg_440_pp0_iter4_reg;
reg   [3:0] trunc_ln150_reg_440_pp0_iter5_reg;
reg   [3:0] trunc_ln150_reg_440_pp0_iter6_reg;
wire   [4:0] add_ln149_fu_233_p2;
wire   [6:0] select_ln148_12_fu_245_p3;
wire   [1:0] select_ln147_11_fu_287_p3;
reg   [1:0] select_ln147_11_reg_455;
reg    ap_enable_reg_pp0_iter1;
wire   [3:0] select_ln148_11_fu_370_p3;
reg   [3:0] select_ln148_11_reg_460;
reg   [3:0] select_ln148_11_reg_460_pp0_iter2_reg;
reg   [3:0] select_ln148_11_reg_460_pp0_iter3_reg;
reg   [3:0] select_ln148_11_reg_460_pp0_iter4_reg;
reg   [3:0] select_ln148_11_reg_460_pp0_iter5_reg;
reg   [3:0] select_ln148_11_reg_460_pp0_iter6_reg;
reg   [15:0] ifmap_vec_load_reg_475;
reg   [15:0] weight_vecs_0_load_reg_480;
wire   [15:0] grp_fu_153_p2;
reg   [15:0] mul_reg_485;
reg    ap_block_state1;
wire    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_flush_enable;
reg    ap_enable_reg_pp0_iter2;
reg    ap_condition_pp0_exit_iter1_state3;
reg    ap_enable_reg_pp0_iter3;
reg    ap_enable_reg_pp0_iter4;
reg    ap_enable_reg_pp0_iter5;
reg    ap_enable_reg_pp0_iter6;
reg    ap_enable_reg_pp0_iter7;
reg   [1:0] ap_phi_mux_jj_phi_fu_123_p4;
wire    ap_block_pp0_stage0;
reg   [1:0] ap_phi_mux_ii_phi_fu_146_p4;
wire   [63:0] p_cast25_fu_386_p1;
wire   [63:0] idxprom30_fu_398_p1;
wire   [0:0] icmp_ln149_fu_189_p2;
wire   [0:0] xor_ln147_fu_183_p2;
wire   [1:0] select_ln147_fu_175_p3;
wire   [0:0] or_ln148_fu_207_p2;
wire   [6:0] add_ln148_4_fu_239_p2;
wire   [3:0] shl_ln_fu_257_p3;
wire   [3:0] zext_ln150_fu_253_p1;
wire   [3:0] sub_ln150_fu_265_p2;
wire   [3:0] zext_ln150_4_fu_271_p1;
wire   [1:0] add_ln147_fu_281_p2;
wire   [3:0] tmp_fu_298_p3;
wire   [3:0] select_ln147_14_cast_fu_294_p1;
wire   [3:0] shl_ln150_mid1_fu_316_p3;
wire   [3:0] zext_ln150_8_fu_312_p1;
wire   [3:0] sub_ln150_4_fu_324_p2;
wire   [3:0] add_ln150_fu_275_p2;
wire   [3:0] empty_98_fu_306_p2;
wire   [3:0] select_ln148_13_cast_fu_344_p1;
wire   [3:0] empty_99_fu_347_p2;
wire   [3:0] select_ln147_12_fu_330_p3;
wire   [3:0] zext_ln150_9_fu_361_p1;
wire   [3:0] add_ln150_4_fu_364_p2;
wire   [3:0] select_ln147_13_fu_337_p3;
wire   [7:0] tmp_100_cast_fu_353_p3;
wire   [7:0] select_ln148_cast_fu_377_p1;
wire   [7:0] empty_100_fu_380_p2;
wire   [7:0] p_fu_392_p3;
wire    ap_CS_fsm_state10;
reg   [2:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
#0 ap_enable_reg_pp0_iter4 = 1'b0;
#0 ap_enable_reg_pp0_iter5 = 1'b0;
#0 ap_enable_reg_pp0_iter6 = 1'b0;
#0 ap_enable_reg_pp0_iter7 = 1'b0;
end

td_fused_top_hmul_16ns_16ns_16_4_max_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hmul_16ns_16ns_16_4_max_dsp_1_U216(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(ifmap_vec_load_reg_475),
    .din1(weight_vecs_0_load_reg_480),
    .dout(grp_fu_153_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state10)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if ((1'b1 == ap_condition_pp0_flush_enable)) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            if ((1'b1 == ap_condition_pp0_exit_iter1_state3)) begin
                ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter0;
            end else if ((1'b1 == 1'b1)) begin
                ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
            end
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter4 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter5 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter5 <= ap_enable_reg_pp0_iter4;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter6 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter6 <= ap_enable_reg_pp0_iter5;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter7 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter7 <= ap_enable_reg_pp0_iter6;
        end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter7 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_fu_163_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ic_reg_131 <= add_ln149_fu_233_p2;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ic_reg_131 <= 5'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_reg_408_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        ii_reg_142 <= select_ln147_11_reg_455;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ii_reg_142 <= 2'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_fu_163_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        indvar_flatten17_reg_97 <= add_ln147_4_fu_157_p2;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indvar_flatten17_reg_97 <= 8'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_fu_163_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        indvar_flatten_reg_108 <= select_ln148_12_fu_245_p3;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indvar_flatten_reg_108 <= 7'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_reg_408 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        jj_reg_119 <= select_ln148_10_reg_434;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        jj_reg_119 <= 2'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_fu_163_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        add_ln148_reg_424 <= add_ln148_fu_201_p2;
        and_ln147_reg_419 <= and_ln147_fu_195_p2;
        icmp_ln148_reg_412 <= icmp_ln148_fu_169_p2;
        select_ln148_reg_429 <= select_ln148_fu_213_p3;
        trunc_ln150_reg_440 <= trunc_ln150_fu_229_p1;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln147_reg_408 <= icmp_ln147_fu_163_p2;
        icmp_ln147_reg_408_pp0_iter1_reg <= icmp_ln147_reg_408;
        trunc_ln150_reg_440_pp0_iter1_reg <= trunc_ln150_reg_440;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        icmp_ln147_reg_408_pp0_iter2_reg <= icmp_ln147_reg_408_pp0_iter1_reg;
        icmp_ln147_reg_408_pp0_iter3_reg <= icmp_ln147_reg_408_pp0_iter2_reg;
        icmp_ln147_reg_408_pp0_iter4_reg <= icmp_ln147_reg_408_pp0_iter3_reg;
        icmp_ln147_reg_408_pp0_iter5_reg <= icmp_ln147_reg_408_pp0_iter4_reg;
        icmp_ln147_reg_408_pp0_iter6_reg <= icmp_ln147_reg_408_pp0_iter5_reg;
        select_ln148_11_reg_460_pp0_iter2_reg <= select_ln148_11_reg_460;
        select_ln148_11_reg_460_pp0_iter3_reg <= select_ln148_11_reg_460_pp0_iter2_reg;
        select_ln148_11_reg_460_pp0_iter4_reg <= select_ln148_11_reg_460_pp0_iter3_reg;
        select_ln148_11_reg_460_pp0_iter5_reg <= select_ln148_11_reg_460_pp0_iter4_reg;
        select_ln148_11_reg_460_pp0_iter6_reg <= select_ln148_11_reg_460_pp0_iter5_reg;
        trunc_ln150_reg_440_pp0_iter2_reg <= trunc_ln150_reg_440_pp0_iter1_reg;
        trunc_ln150_reg_440_pp0_iter3_reg <= trunc_ln150_reg_440_pp0_iter2_reg;
        trunc_ln150_reg_440_pp0_iter4_reg <= trunc_ln150_reg_440_pp0_iter3_reg;
        trunc_ln150_reg_440_pp0_iter5_reg <= trunc_ln150_reg_440_pp0_iter4_reg;
        trunc_ln150_reg_440_pp0_iter6_reg <= trunc_ln150_reg_440_pp0_iter5_reg;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_reg_408_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        ifmap_vec_load_reg_475 <= ifmap_vec_q0;
        weight_vecs_0_load_reg_480 <= weight_vecs_0_q0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_reg_408_pp0_iter5_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        mul_reg_485 <= grp_fu_153_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_reg_408 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        select_ln147_11_reg_455 <= select_ln147_11_fu_287_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_fu_163_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        select_ln148_10_reg_434 <= select_ln148_10_fu_221_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_reg_408 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        select_ln148_11_reg_460 <= select_ln148_11_fu_370_p3;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_condition_pp0_exit_iter1_state3 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter1_state3 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln147_fu_163_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_condition_pp0_flush_enable = 1'b1;
    end else begin
        ap_condition_pp0_flush_enable = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state10)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter7 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln147_reg_408_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        ap_phi_mux_ii_phi_fu_146_p4 = select_ln147_11_reg_455;
    end else begin
        ap_phi_mux_ii_phi_fu_146_p4 = ii_reg_142;
    end
end

always @ (*) begin
    if (((icmp_ln147_reg_408 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_jj_phi_fu_123_p4 = select_ln148_10_reg_434;
    end else begin
        ap_phi_mux_jj_phi_fu_123_p4 = jj_reg_119;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state10)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ifmap_vec_ce0 = 1'b1;
    end else begin
        ifmap_vec_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter7 == 1'b1))) begin
        products_0_ce0 = 1'b1;
    end else begin
        products_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln147_reg_408_pp0_iter6_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter7 == 1'b1))) begin
        products_0_we0 = 1'b1;
    end else begin
        products_0_we0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        weight_vecs_0_ce0 = 1'b1;
    end else begin
        weight_vecs_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((~((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b1)) & ~((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter7 == 1'b1) & (ap_enable_reg_pp0_iter6 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if ((((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter7 == 1'b1) & (ap_enable_reg_pp0_iter6 == 1'b0)) | ((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b1)))) begin
                ap_NS_fsm = ap_ST_fsm_state10;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state10 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln147_4_fu_157_p2 = (indvar_flatten17_reg_97 + 8'd1);

assign add_ln147_fu_281_p2 = (ap_phi_mux_ii_phi_fu_146_p4 + 2'd1);

assign add_ln148_4_fu_239_p2 = (indvar_flatten_reg_108 + 7'd1);

assign add_ln148_fu_201_p2 = (select_ln147_fu_175_p3 + 2'd1);

assign add_ln149_fu_233_p2 = (select_ln148_fu_213_p3 + 5'd1);

assign add_ln150_4_fu_364_p2 = (select_ln147_12_fu_330_p3 + zext_ln150_9_fu_361_p1);

assign add_ln150_fu_275_p2 = (sub_ln150_fu_265_p2 + zext_ln150_4_fu_271_p1);

assign and_ln147_fu_195_p2 = (xor_ln147_fu_183_p2 & icmp_ln149_fu_189_p2);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state10 = ap_CS_fsm[32'd2];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (ap_done_reg == 1'b1));
end

assign ap_block_state2_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter4 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage0_iter5 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage0_iter6 = ~(1'b1 == 1'b1);

assign ap_block_state9_pp0_stage0_iter7 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign empty_100_fu_380_p2 = (tmp_100_cast_fu_353_p3 + select_ln148_cast_fu_377_p1);

assign empty_98_fu_306_p2 = (tmp_fu_298_p3 - select_ln147_14_cast_fu_294_p1);

assign empty_99_fu_347_p2 = (empty_98_fu_306_p2 + select_ln148_13_cast_fu_344_p1);

assign icmp_ln147_fu_163_p2 = ((indvar_flatten17_reg_97 == 8'd144) ? 1'b1 : 1'b0);

assign icmp_ln148_fu_169_p2 = ((indvar_flatten_reg_108 == 7'd48) ? 1'b1 : 1'b0);

assign icmp_ln149_fu_189_p2 = ((ic_reg_131 == 5'd16) ? 1'b1 : 1'b0);

assign idxprom30_fu_398_p1 = p_fu_392_p3;

assign ifmap_vec_address0 = p_cast25_fu_386_p1;

assign or_ln148_fu_207_p2 = (icmp_ln148_fu_169_p2 | and_ln147_fu_195_p2);

assign p_cast25_fu_386_p1 = empty_100_fu_380_p2;

assign p_fu_392_p3 = {{select_ln148_11_reg_460_pp0_iter6_reg}, {trunc_ln150_reg_440_pp0_iter6_reg}};

assign products_0_address0 = idxprom30_fu_398_p1;

assign products_0_d0 = mul_reg_485;

assign select_ln147_11_fu_287_p3 = ((icmp_ln148_reg_412[0:0] == 1'b1) ? add_ln147_fu_281_p2 : ap_phi_mux_ii_phi_fu_146_p4);

assign select_ln147_12_fu_330_p3 = ((icmp_ln148_reg_412[0:0] == 1'b1) ? sub_ln150_4_fu_324_p2 : sub_ln150_fu_265_p2);

assign select_ln147_13_fu_337_p3 = ((icmp_ln148_reg_412[0:0] == 1'b1) ? sub_ln150_4_fu_324_p2 : add_ln150_fu_275_p2);

assign select_ln147_14_cast_fu_294_p1 = select_ln147_11_fu_287_p3;

assign select_ln147_fu_175_p3 = ((icmp_ln148_fu_169_p2[0:0] == 1'b1) ? 2'd0 : ap_phi_mux_jj_phi_fu_123_p4);

assign select_ln148_10_fu_221_p3 = ((and_ln147_fu_195_p2[0:0] == 1'b1) ? add_ln148_fu_201_p2 : select_ln147_fu_175_p3);

assign select_ln148_11_fu_370_p3 = ((and_ln147_reg_419[0:0] == 1'b1) ? add_ln150_4_fu_364_p2 : select_ln147_13_fu_337_p3);

assign select_ln148_12_fu_245_p3 = ((icmp_ln148_fu_169_p2[0:0] == 1'b1) ? 7'd1 : add_ln148_4_fu_239_p2);

assign select_ln148_13_cast_fu_344_p1 = select_ln148_10_reg_434;

assign select_ln148_cast_fu_377_p1 = select_ln148_reg_429;

assign select_ln148_fu_213_p3 = ((or_ln148_fu_207_p2[0:0] == 1'b1) ? 5'd0 : ic_reg_131);

assign shl_ln150_mid1_fu_316_p3 = {{add_ln147_fu_281_p2}, {2'd0}};

assign shl_ln_fu_257_p3 = {{ap_phi_mux_ii_phi_fu_146_p4}, {2'd0}};

assign sub_ln150_4_fu_324_p2 = (shl_ln150_mid1_fu_316_p3 - zext_ln150_8_fu_312_p1);

assign sub_ln150_fu_265_p2 = (shl_ln_fu_257_p3 - zext_ln150_fu_253_p1);

assign tmp_100_cast_fu_353_p3 = {{empty_99_fu_347_p2}, {4'd0}};

assign tmp_fu_298_p3 = {{select_ln147_11_fu_287_p3}, {2'd0}};

assign trunc_ln150_fu_229_p1 = select_ln148_fu_213_p3[3:0];

assign weight_vecs_0_address0 = p_cast25_fu_386_p1;

assign xor_ln147_fu_183_p2 = (icmp_ln148_fu_169_p2 ^ 1'd1);

assign zext_ln150_4_fu_271_p1 = jj_reg_119;

assign zext_ln150_8_fu_312_p1 = add_ln147_fu_281_p2;

assign zext_ln150_9_fu_361_p1 = add_ln148_reg_424;

assign zext_ln150_fu_253_p1 = ap_phi_mux_ii_phi_fu_146_p4;

endmodule //td_fused_top_tdf4_dot_product
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_tdf4_filters_ram (addr0, ce0, q0, addr1, ce1, d1, we1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 15;
parameter MEM_SIZE = 18432;

input[AWIDTH-1:0] addr0;
input ce0;
output wire[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
input clk;

 reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];
wire [AWIDTH-1:0] addr0_t0; 
reg [AWIDTH-1:0] addr0_t1; 
reg [DWIDTH-1:0] q0_t0;
reg [DWIDTH-1:0] q0_t1;
wire [AWIDTH-1:0] addr1_t0; 
reg [AWIDTH-1:0] addr1_t1; 
wire [DWIDTH-1:0] d1_t0; 
wire we1_t0; 
reg [DWIDTH-1:0] d1_t1; 
reg we1_t1; 


assign addr0_t0 = addr0;
assign q0 = q0_t1;
assign addr1_t0 = addr1;
assign d1_t0 = d1;
assign we1_t0 = we1;

always @(posedge clk)  
begin
    if (ce0) 
    begin
        addr0_t1 <= addr0_t0; 
        q0_t1 <= q0_t0;
    end
    if (ce1) 
    begin
        addr1_t1 <= addr1_t0; 
        d1_t1 <= d1_t0;
        we1_t1 <= we1_t0;
    end
end


always @(posedge clk)  
begin 
    if (ce0) begin
        q0_t0 <= ram[addr0_t1];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1_t1) 
            ram[addr1_t1] <= d1_t1; 
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_tdf4_filters(
    reset,
    clk,
    address0,
    ce0,
    q0,
    address1,
    ce1,
    we1,
    d1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd18432;
parameter AddressWidth = 32'd15;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;



td_fused_top_tdf4_filters_ram td_fused_top_tdf4_filters_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 )
);

endmodule

// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf4_get_next_ijk (
        ap_clk,
        ap_rst,
        ap_start,
        start_full_n,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        start_out,
        start_write,
        indices_0_din,
        indices_0_full_n,
        indices_0_write,
        indices_1_din,
        indices_1_full_n,
        indices_1_write,
        indices_2_out_din,
        indices_2_out_full_n,
        indices_2_out_write,
        indices_2_out1_din,
        indices_2_out1_full_n,
        indices_2_out1_write,
        write_r_din,
        write_r_full_n,
        write_r_write
);

parameter    ap_ST_fsm_state1 = 1'd1;

input   ap_clk;
input   ap_rst;
input   ap_start;
input   start_full_n;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output   start_out;
output   start_write;
output  [15:0] indices_0_din;
input   indices_0_full_n;
output   indices_0_write;
output  [15:0] indices_1_din;
input   indices_1_full_n;
output   indices_1_write;
output  [6:0] indices_2_out_din;
input   indices_2_out_full_n;
output   indices_2_out_write;
output  [10:0] indices_2_out1_din;
input   indices_2_out1_full_n;
output   indices_2_out1_write;
output   write_r_din;
input   write_r_full_n;
output   write_r_write;

reg ap_done;
reg ap_idle;
reg start_write;
reg indices_0_write;
reg indices_1_write;
reg indices_2_out_write;
reg indices_2_out1_write;
reg write_r_write;

reg    real_start;
reg    start_once_reg;
reg    ap_done_reg;
  reg   [0:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    internal_ap_ready;
reg   [15:0] i_4;
reg   [15:0] j_4;
reg   [15:0] k_4;
reg    indices_0_blk_n;
reg    indices_1_blk_n;
reg    indices_2_out_blk_n;
reg    indices_2_out1_blk_n;
reg    write_r_blk_n;
reg   [0:0] ap_phi_mux_j_15_flag_0_i_phi_fu_92_p6;
reg    ap_block_state1;
wire   [0:0] icmp_ln188_fu_167_p2;
wire   [0:0] icmp_ln191_fu_180_p2;
reg   [15:0] ap_phi_mux_j_15_new_0_i_phi_fu_106_p6;
wire   [15:0] add_ln190_fu_173_p2;
reg   [15:0] ap_phi_mux_k_15_new_0_i_phi_fu_119_p6;
wire   [15:0] add_ln187_fu_160_p2;
wire   [15:0] select_ln194_fu_198_p3;
wire   [15:0] add_ln193_fu_186_p2;
wire   [0:0] icmp_ln194_fu_192_p2;
reg   [0:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 start_once_reg = 1'b0;
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 1'd1;
#0 i_4 = 16'd0;
#0 j_4 = 16'd0;
#0 k_4 = 16'd0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((~((real_start == 1'b0) | (write_r_full_n == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        start_once_reg <= 1'b0;
    end else begin
        if (((real_start == 1'b1) & (internal_ap_ready == 1'b0))) begin
            start_once_reg <= 1'b1;
        end else if ((internal_ap_ready == 1'b1)) begin
            start_once_reg <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((~((real_start == 1'b0) | (write_r_full_n == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (icmp_ln191_fu_180_p2 == 1'd1) & (icmp_ln188_fu_167_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1))) begin
        i_4 <= select_ln194_fu_198_p3;
    end
end

always @ (posedge ap_clk) begin
    if ((~((real_start == 1'b0) | (write_r_full_n == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (ap_phi_mux_j_15_flag_0_i_phi_fu_92_p6 == 1'd1) & (1'b1 == ap_CS_fsm_state1))) begin
        j_4 <= ap_phi_mux_j_15_new_0_i_phi_fu_106_p6;
    end
end

always @ (posedge ap_clk) begin
    if ((~((real_start == 1'b0) | (write_r_full_n == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        k_4 <= ap_phi_mux_k_15_new_0_i_phi_fu_119_p6;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (write_r_full_n == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((real_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln188_fu_167_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_phi_mux_j_15_flag_0_i_phi_fu_92_p6 = 1'd0;
    end else if ((((icmp_ln191_fu_180_p2 == 1'd0) & (icmp_ln188_fu_167_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1)) | ((icmp_ln191_fu_180_p2 == 1'd1) & (icmp_ln188_fu_167_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1)))) begin
        ap_phi_mux_j_15_flag_0_i_phi_fu_92_p6 = 1'd1;
    end else begin
        ap_phi_mux_j_15_flag_0_i_phi_fu_92_p6 = 'bx;
    end
end

always @ (*) begin
    if (((icmp_ln188_fu_167_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1))) begin
        if ((icmp_ln191_fu_180_p2 == 1'd0)) begin
            ap_phi_mux_j_15_new_0_i_phi_fu_106_p6 = add_ln190_fu_173_p2;
        end else if ((icmp_ln191_fu_180_p2 == 1'd1)) begin
            ap_phi_mux_j_15_new_0_i_phi_fu_106_p6 = 16'd0;
        end else begin
            ap_phi_mux_j_15_new_0_i_phi_fu_106_p6 = 'bx;
        end
    end else begin
        ap_phi_mux_j_15_new_0_i_phi_fu_106_p6 = 'bx;
    end
end

always @ (*) begin
    if (((icmp_ln188_fu_167_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_phi_mux_k_15_new_0_i_phi_fu_119_p6 = add_ln187_fu_160_p2;
    end else if ((((icmp_ln191_fu_180_p2 == 1'd0) & (icmp_ln188_fu_167_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1)) | ((icmp_ln191_fu_180_p2 == 1'd1) & (icmp_ln188_fu_167_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1)))) begin
        ap_phi_mux_k_15_new_0_i_phi_fu_119_p6 = 16'd0;
    end else begin
        ap_phi_mux_k_15_new_0_i_phi_fu_119_p6 = 'bx;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_0_blk_n = indices_0_full_n;
    end else begin
        indices_0_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (write_r_full_n == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_0_write = 1'b1;
    end else begin
        indices_0_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_1_blk_n = indices_1_full_n;
    end else begin
        indices_1_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (write_r_full_n == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_1_write = 1'b1;
    end else begin
        indices_1_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_2_out1_blk_n = indices_2_out1_full_n;
    end else begin
        indices_2_out1_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (write_r_full_n == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_2_out1_write = 1'b1;
    end else begin
        indices_2_out1_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_2_out_blk_n = indices_2_out_full_n;
    end else begin
        indices_2_out_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (write_r_full_n == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_2_out_write = 1'b1;
    end else begin
        indices_2_out_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (write_r_full_n == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        internal_ap_ready = 1'b1;
    end else begin
        internal_ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((start_full_n == 1'b0) & (start_once_reg == 1'b0))) begin
        real_start = 1'b0;
    end else begin
        real_start = ap_start;
    end
end

always @ (*) begin
    if (((real_start == 1'b1) & (start_once_reg == 1'b0))) begin
        start_write = 1'b1;
    end else begin
        start_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        write_r_blk_n = write_r_full_n;
    end else begin
        write_r_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (write_r_full_n == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        write_r_write = 1'b1;
    end else begin
        write_r_write = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln187_fu_160_p2 = (k_4 + 16'd1);

assign add_ln190_fu_173_p2 = (j_4 + 16'd1);

assign add_ln193_fu_186_p2 = (i_4 + 16'd1);

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

always @ (*) begin
    ap_block_state1 = ((real_start == 1'b0) | (write_r_full_n == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1));
end

assign ap_ready = internal_ap_ready;

assign icmp_ln188_fu_167_p2 = ((add_ln187_fu_160_p2 == 16'd128) ? 1'b1 : 1'b0);

assign icmp_ln191_fu_180_p2 = ((add_ln190_fu_173_p2 == 16'd56) ? 1'b1 : 1'b0);

assign icmp_ln194_fu_192_p2 = ((add_ln193_fu_186_p2 == 16'd56) ? 1'b1 : 1'b0);

assign indices_0_din = i_4;

assign indices_1_din = j_4;

assign indices_2_out1_din = k_4[10:0];

assign indices_2_out_din = k_4[6:0];

assign select_ln194_fu_198_p3 = ((icmp_ln194_fu_192_p2[0:0] == 1'b1) ? 16'd0 : add_ln193_fu_186_p2);

assign start_out = real_start;

assign write_r_din = ((k_4 == 16'd127) ? 1'b1 : 1'b0);

endmodule //td_fused_top_tdf4_get_next_ijk
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_tdf4_l2_filters_ram (addr0, ce0, q0, addr1, ce1, d1, we1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 11;
parameter MEM_SIZE = 2048;

input[AWIDTH-1:0] addr0;
input ce0;
output wire[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
input clk;

 reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];
wire [AWIDTH-1:0] addr0_t0; 
reg [AWIDTH-1:0] addr0_t1; 
reg [DWIDTH-1:0] q0_t0;
reg [DWIDTH-1:0] q0_t1;
wire [AWIDTH-1:0] addr1_t0; 
reg [AWIDTH-1:0] addr1_t1; 
wire [DWIDTH-1:0] d1_t0; 
wire we1_t0; 
reg [DWIDTH-1:0] d1_t1; 
reg we1_t1; 


assign addr0_t0 = addr0;
assign q0 = q0_t1;
assign addr1_t0 = addr1;
assign d1_t0 = d1;
assign we1_t0 = we1;

always @(posedge clk)  
begin
    if (ce0) 
    begin
        addr0_t1 <= addr0_t0; 
        q0_t1 <= q0_t0;
    end
    if (ce1) 
    begin
        addr1_t1 <= addr1_t0; 
        d1_t1 <= d1_t0;
        we1_t1 <= we1_t0;
    end
end


always @(posedge clk)  
begin 
    if (ce0) begin
        q0_t0 <= ram[addr0_t1];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1_t1) 
            ram[addr1_t1] <= d1_t1; 
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_tdf4_l2_filters(
    reset,
    clk,
    address0,
    ce0,
    q0,
    address1,
    ce1,
    we1,
    d1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd2048;
parameter AddressWidth = 32'd11;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;



td_fused_top_tdf4_l2_filters_ram td_fused_top_tdf4_l2_filters_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 )
);

endmodule

// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf4_l2_multiply34 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        intermediate_fmaps_read,
        l2_filter_data_address0,
        l2_filter_data_ce0,
        l2_filter_data_q0,
        l2_products_address0,
        l2_products_ce0,
        l2_products_we0,
        l2_products_d0,
        indices_23_dout,
        indices_23_empty_n,
        indices_23_read
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state10 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
input  [15:0] intermediate_fmaps_read;
output  [10:0] l2_filter_data_address0;
output   l2_filter_data_ce0;
input  [15:0] l2_filter_data_q0;
output  [3:0] l2_products_address0;
output   l2_products_ce0;
output   l2_products_we0;
output  [15:0] l2_products_d0;
input  [10:0] indices_23_dout;
input   indices_23_empty_n;
output   indices_23_read;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg l2_filter_data_ce0;
reg l2_products_ce0;
reg l2_products_we0;
reg indices_23_read;

reg    ap_done_reg;
  reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    indices_23_blk_n;
reg   [4:0] i_1_1_reg_106;
reg   [10:0] l2_ichan_reg_165;
wire   [4:0] add_ln20_fu_122_p2;
wire    ap_CS_fsm_pp0_stage0;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
wire    ap_block_state4_pp0_stage0_iter2;
wire    ap_block_state5_pp0_stage0_iter3;
wire    ap_block_state6_pp0_stage0_iter4;
wire    ap_block_state7_pp0_stage0_iter5;
wire    ap_block_state8_pp0_stage0_iter6;
wire    ap_block_state9_pp0_stage0_iter7;
wire    ap_block_pp0_stage0_11001;
wire   [0:0] icmp_ln20_fu_128_p2;
reg   [0:0] icmp_ln20_reg_175;
reg   [0:0] icmp_ln20_reg_175_pp0_iter1_reg;
reg   [0:0] icmp_ln20_reg_175_pp0_iter2_reg;
reg   [0:0] icmp_ln20_reg_175_pp0_iter3_reg;
reg   [0:0] icmp_ln20_reg_175_pp0_iter4_reg;
reg   [0:0] icmp_ln20_reg_175_pp0_iter5_reg;
reg   [0:0] icmp_ln20_reg_175_pp0_iter6_reg;
wire   [3:0] l2_o_fu_134_p1;
reg   [3:0] l2_o_reg_179;
reg   [3:0] l2_o_reg_179_pp0_iter1_reg;
reg   [3:0] l2_o_reg_179_pp0_iter2_reg;
reg   [3:0] l2_o_reg_179_pp0_iter3_reg;
reg   [3:0] l2_o_reg_179_pp0_iter4_reg;
reg   [3:0] l2_o_reg_179_pp0_iter5_reg;
reg   [3:0] l2_o_reg_179_pp0_iter6_reg;
wire   [15:0] grp_fu_117_p2;
reg   [15:0] mul_i_i_reg_194;
reg    ap_block_state1;
wire    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_exit_iter0_state2;
reg    ap_enable_reg_pp0_iter1;
reg    ap_enable_reg_pp0_iter2;
reg    ap_enable_reg_pp0_iter3;
reg    ap_enable_reg_pp0_iter4;
reg    ap_enable_reg_pp0_iter5;
reg    ap_enable_reg_pp0_iter6;
reg    ap_enable_reg_pp0_iter7;
wire   [63:0] zext_ln29_13_fu_151_p1;
wire    ap_block_pp0_stage0;
wire   [63:0] zext_ln29_fu_156_p1;
wire   [10:0] tmp_s_fu_138_p3;
wire   [10:0] add_ln29_fu_146_p2;
wire    ap_CS_fsm_state10;
reg   [2:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
#0 ap_enable_reg_pp0_iter4 = 1'b0;
#0 ap_enable_reg_pp0_iter5 = 1'b0;
#0 ap_enable_reg_pp0_iter6 = 1'b0;
#0 ap_enable_reg_pp0_iter7 = 1'b0;
end

td_fused_top_hmul_16ns_16ns_16_4_max_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hmul_16ns_16ns_16_4_max_dsp_1_U235(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(l2_filter_data_q0),
    .din1(intermediate_fmaps_read),
    .dout(grp_fu_117_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state10)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b1 == ap_condition_pp0_exit_iter0_state2))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            if ((1'b1 == ap_condition_pp0_exit_iter0_state2)) begin
                ap_enable_reg_pp0_iter1 <= (1'b1 ^ ap_condition_pp0_exit_iter0_state2);
            end else if ((1'b1 == 1'b1)) begin
                ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
            end
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter4 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter5 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter5 <= ap_enable_reg_pp0_iter4;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter6 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter6 <= ap_enable_reg_pp0_iter5;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter7 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter7 <= ap_enable_reg_pp0_iter6;
        end else if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter7 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        i_1_1_reg_106 <= 5'd0;
    end else if (((icmp_ln20_fu_128_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        i_1_1_reg_106 <= add_ln20_fu_122_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln20_reg_175 <= icmp_ln20_fu_128_p2;
        icmp_ln20_reg_175_pp0_iter1_reg <= icmp_ln20_reg_175;
        l2_o_reg_179_pp0_iter1_reg <= l2_o_reg_179;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        icmp_ln20_reg_175_pp0_iter2_reg <= icmp_ln20_reg_175_pp0_iter1_reg;
        icmp_ln20_reg_175_pp0_iter3_reg <= icmp_ln20_reg_175_pp0_iter2_reg;
        icmp_ln20_reg_175_pp0_iter4_reg <= icmp_ln20_reg_175_pp0_iter3_reg;
        icmp_ln20_reg_175_pp0_iter5_reg <= icmp_ln20_reg_175_pp0_iter4_reg;
        icmp_ln20_reg_175_pp0_iter6_reg <= icmp_ln20_reg_175_pp0_iter5_reg;
        l2_o_reg_179_pp0_iter2_reg <= l2_o_reg_179_pp0_iter1_reg;
        l2_o_reg_179_pp0_iter3_reg <= l2_o_reg_179_pp0_iter2_reg;
        l2_o_reg_179_pp0_iter4_reg <= l2_o_reg_179_pp0_iter3_reg;
        l2_o_reg_179_pp0_iter5_reg <= l2_o_reg_179_pp0_iter4_reg;
        l2_o_reg_179_pp0_iter6_reg <= l2_o_reg_179_pp0_iter5_reg;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state1)) begin
        l2_ichan_reg_165 <= indices_23_dout;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln20_fu_128_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        l2_o_reg_179 <= l2_o_fu_134_p1;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln20_reg_175_pp0_iter5_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        mul_i_i_reg_194 <= grp_fu_117_p2;
    end
end

always @ (*) begin
    if ((icmp_ln20_fu_128_p2 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state2 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state2 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state10)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter7 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state10)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_23_blk_n = indices_23_empty_n;
    end else begin
        indices_23_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_23_read = 1'b1;
    end else begin
        indices_23_read = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter3 == 1'b1)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1)))) begin
        l2_filter_data_ce0 = 1'b1;
    end else begin
        l2_filter_data_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter7 == 1'b1))) begin
        l2_products_ce0 = 1'b1;
    end else begin
        l2_products_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln20_reg_175_pp0_iter6_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter7 == 1'b1))) begin
        l2_products_we0 = 1'b1;
    end else begin
        l2_products_we0 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((~((icmp_ln20_fu_128_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0)) & ~((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter7 == 1'b1) & (ap_enable_reg_pp0_iter6 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if ((((icmp_ln20_fu_128_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0)) | ((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter7 == 1'b1) & (ap_enable_reg_pp0_iter6 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_state10;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state10 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln20_fu_122_p2 = (i_1_1_reg_106 + 5'd1);

assign add_ln29_fu_146_p2 = (tmp_s_fu_138_p3 + l2_ichan_reg_165);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state10 = ap_CS_fsm[32'd2];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1));
end

assign ap_block_state2_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter4 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage0_iter5 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage0_iter6 = ~(1'b1 == 1'b1);

assign ap_block_state9_pp0_stage0_iter7 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign icmp_ln20_fu_128_p2 = ((i_1_1_reg_106 == 5'd16) ? 1'b1 : 1'b0);

assign l2_filter_data_address0 = zext_ln29_13_fu_151_p1;

assign l2_o_fu_134_p1 = i_1_1_reg_106[3:0];

assign l2_products_address0 = zext_ln29_fu_156_p1;

assign l2_products_d0 = mul_i_i_reg_194;

assign tmp_s_fu_138_p3 = {{l2_o_fu_134_p1}, {7'd0}};

assign zext_ln29_13_fu_151_p1 = add_ln29_fu_146_p2;

assign zext_ln29_fu_156_p1 = l2_o_reg_179_pp0_iter6_reg;

endmodule //td_fused_top_tdf4_l2_multiply34
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_tdf4_l2_writeOutputs_133_running_sums_1_ram (addr0, ce0, d0, we0, addr1, ce1, q1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 4;
parameter MEM_SIZE = 16;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
input[AWIDTH-1:0] addr1;
input ce1;
output reg[DWIDTH-1:0] q1;
input clk;

 reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];

//initial begin
//    $readmemh("./td_fused_top_tdf4_l2_writeOutputs_133_running_sums_1_ram.dat", ram);
//end



always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        q1 <= ram[addr1];
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_tdf4_l2_writeOutputs_133_running_sums_1(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    address1,
    ce1,
    q1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16;
parameter AddressWidth = 32'd4;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
input[AddressWidth - 1:0] address1;
input ce1;
output[DataWidth - 1:0] q1;



td_fused_top_tdf4_l2_writeOutputs_133_running_sums_1_ram td_fused_top_tdf4_l2_writeOutputs_133_running_sums_1_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .q1( q1 )
);

endmodule

// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf4_l2_writeOutputs_133 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        indices_01_dout,
        indices_01_empty_n,
        indices_01_read,
        indices_12_dout,
        indices_12_empty_n,
        indices_12_read,
        write4_dout,
        write4_empty_n,
        write4_read,
        l2_partial_sums_address0,
        l2_partial_sums_ce0,
        l2_partial_sums_q0,
        out_data_address1,
        out_data_ce1,
        out_data_we1,
        out_data_d1,
        l2_adjustments_address0,
        l2_adjustments_ce0,
        l2_adjustments_q0
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state25 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
input  [5:0] indices_01_dout;
input   indices_01_empty_n;
output   indices_01_read;
input  [11:0] indices_12_dout;
input   indices_12_empty_n;
output   indices_12_read;
input  [0:0] write4_dout;
input   write4_empty_n;
output   write4_read;
output  [3:0] l2_partial_sums_address0;
output   l2_partial_sums_ce0;
input  [15:0] l2_partial_sums_q0;
output  [13:0] out_data_address1;
output   out_data_ce1;
output   out_data_we1;
output  [63:0] out_data_d1;
output  [3:0] l2_adjustments_address0;
output   l2_adjustments_ce0;
input  [47:0] l2_adjustments_q0;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg indices_01_read;
reg indices_12_read;
reg write4_read;
reg l2_partial_sums_ce0;
reg out_data_ce1;
reg out_data_we1;
reg l2_adjustments_ce0;

reg    ap_done_reg;
  reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    running_sums_1_ce0;
reg    running_sums_1_we0;
wire   [15:0] running_sums_1_d0;
wire   [3:0] running_sums_1_address1;
reg    running_sums_1_ce1;
wire   [15:0] running_sums_1_q1;
reg    indices_01_blk_n;
reg    indices_12_blk_n;
reg    write4_blk_n;
reg   [4:0] ochan_reg_208;
reg   [0:0] write4_read_reg_567;
wire   [13:0] add_ln109_fu_273_p2;
reg   [13:0] add_ln109_reg_573;
wire   [4:0] add_ln86_fu_279_p2;
wire    ap_CS_fsm_pp0_stage0;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
wire    ap_block_state4_pp0_stage0_iter2;
wire    ap_block_state5_pp0_stage0_iter3;
wire    ap_block_state6_pp0_stage0_iter4;
wire    ap_block_state7_pp0_stage0_iter5;
wire    ap_block_state8_pp0_stage0_iter6;
wire    ap_block_state9_pp0_stage0_iter7;
wire    ap_block_state10_pp0_stage0_iter8;
wire    ap_block_state11_pp0_stage0_iter9;
wire    ap_block_state12_pp0_stage0_iter10;
wire    ap_block_state13_pp0_stage0_iter11;
wire    ap_block_state14_pp0_stage0_iter12;
wire    ap_block_state15_pp0_stage0_iter13;
wire    ap_block_state16_pp0_stage0_iter14;
wire    ap_block_state17_pp0_stage0_iter15;
wire    ap_block_state18_pp0_stage0_iter16;
wire    ap_block_state19_pp0_stage0_iter17;
wire    ap_block_state20_pp0_stage0_iter18;
wire    ap_block_state21_pp0_stage0_iter19;
wire    ap_block_state22_pp0_stage0_iter20;
wire    ap_block_state23_pp0_stage0_iter21;
wire    ap_block_state24_pp0_stage0_iter22;
wire    ap_block_pp0_stage0_11001;
wire   [0:0] icmp_ln86_fu_285_p2;
wire   [63:0] zext_ln86_fu_291_p1;
reg   [63:0] zext_ln86_reg_587;
reg   [63:0] zext_ln86_reg_587_pp0_iter1_reg;
reg   [63:0] zext_ln86_reg_587_pp0_iter2_reg;
reg   [63:0] zext_ln86_reg_587_pp0_iter3_reg;
reg   [3:0] running_sums_1_addr_reg_597;
reg   [3:0] running_sums_1_addr_reg_597_pp0_iter1_reg;
reg   [3:0] running_sums_1_addr_reg_597_pp0_iter2_reg;
reg   [3:0] running_sums_1_addr_reg_597_pp0_iter3_reg;
reg   [3:0] running_sums_1_addr_reg_597_pp0_iter4_reg;
reg   [3:0] running_sums_1_addr_reg_597_pp0_iter5_reg;
reg   [3:0] running_sums_1_addr_reg_597_pp0_iter6_reg;
wire   [1:0] trunc_ln99_fu_297_p1;
reg   [1:0] trunc_ln99_reg_603;
reg   [1:0] trunc_ln99_reg_603_pp0_iter1_reg;
reg   [1:0] trunc_ln99_reg_603_pp0_iter2_reg;
reg   [1:0] trunc_ln99_reg_603_pp0_iter3_reg;
reg   [1:0] trunc_ln99_reg_603_pp0_iter4_reg;
reg   [1:0] trunc_ln99_reg_603_pp0_iter5_reg;
reg   [1:0] trunc_ln99_reg_603_pp0_iter6_reg;
reg   [1:0] trunc_ln99_reg_603_pp0_iter7_reg;
reg   [1:0] trunc_ln99_reg_603_pp0_iter8_reg;
reg   [1:0] trunc_ln99_reg_603_pp0_iter9_reg;
reg   [1:0] trunc_ln99_reg_603_pp0_iter10_reg;
reg   [1:0] trunc_ln99_reg_603_pp0_iter11_reg;
reg   [1:0] trunc_ln99_reg_603_pp0_iter12_reg;
reg   [1:0] trunc_ln99_reg_603_pp0_iter13_reg;
reg   [1:0] trunc_ln99_reg_603_pp0_iter14_reg;
reg   [1:0] trunc_ln99_reg_603_pp0_iter15_reg;
reg   [1:0] trunc_ln99_reg_603_pp0_iter16_reg;
reg   [1:0] trunc_ln99_reg_603_pp0_iter17_reg;
reg   [1:0] trunc_ln99_reg_603_pp0_iter18_reg;
reg   [1:0] trunc_ln99_reg_603_pp0_iter19_reg;
reg   [1:0] trunc_ln99_reg_603_pp0_iter20_reg;
wire   [0:0] and_ln103_fu_307_p2;
reg   [0:0] and_ln103_reg_610;
reg   [0:0] and_ln103_reg_610_pp0_iter1_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter2_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter3_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter4_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter5_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter6_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter7_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter8_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter9_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter10_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter11_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter12_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter13_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter14_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter15_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter16_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter17_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter18_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter19_reg;
reg   [0:0] and_ln103_reg_610_pp0_iter20_reg;
reg   [1:0] lshr_ln_reg_614;
reg   [1:0] lshr_ln_reg_614_pp0_iter1_reg;
reg   [1:0] lshr_ln_reg_614_pp0_iter2_reg;
reg   [1:0] lshr_ln_reg_614_pp0_iter3_reg;
reg   [1:0] lshr_ln_reg_614_pp0_iter4_reg;
reg   [1:0] lshr_ln_reg_614_pp0_iter5_reg;
reg   [1:0] lshr_ln_reg_614_pp0_iter6_reg;
reg   [1:0] lshr_ln_reg_614_pp0_iter7_reg;
reg   [1:0] lshr_ln_reg_614_pp0_iter8_reg;
reg   [1:0] lshr_ln_reg_614_pp0_iter9_reg;
reg   [1:0] lshr_ln_reg_614_pp0_iter10_reg;
reg   [1:0] lshr_ln_reg_614_pp0_iter11_reg;
reg   [1:0] lshr_ln_reg_614_pp0_iter12_reg;
reg   [1:0] lshr_ln_reg_614_pp0_iter13_reg;
reg   [1:0] lshr_ln_reg_614_pp0_iter14_reg;
reg   [1:0] lshr_ln_reg_614_pp0_iter15_reg;
reg   [1:0] lshr_ln_reg_614_pp0_iter16_reg;
reg   [1:0] lshr_ln_reg_614_pp0_iter17_reg;
reg   [1:0] lshr_ln_reg_614_pp0_iter18_reg;
reg   [1:0] lshr_ln_reg_614_pp0_iter19_reg;
reg   [1:0] lshr_ln_reg_614_pp0_iter20_reg;
reg   [15:0] val_reg_619;
reg   [15:0] running_sums_1_load_reg_624;
reg    ap_enable_reg_pp0_iter1;
wire   [15:0] grp_fu_219_p2;
reg   [15:0] sum_reg_634;
reg   [15:0] tmp_47_i_i_reg_645;
reg   [15:0] tmp_47_i_i_reg_645_pp0_iter8_reg;
reg   [15:0] tmp_47_i_i_reg_645_pp0_iter9_reg;
reg   [15:0] tmp_47_i_i_reg_645_pp0_iter10_reg;
reg   [15:0] tmp_47_i_i_reg_645_pp0_iter11_reg;
reg   [15:0] tmp_48_i_i_reg_650;
reg   [15:0] tmp_48_i_i_reg_650_pp0_iter8_reg;
reg   [15:0] tmp_48_i_i_reg_650_pp0_iter9_reg;
reg   [15:0] tmp_48_i_i_reg_650_pp0_iter10_reg;
reg   [15:0] tmp_48_i_i_reg_650_pp0_iter11_reg;
reg   [15:0] tmp_48_i_i_reg_650_pp0_iter12_reg;
reg   [15:0] tmp_48_i_i_reg_650_pp0_iter13_reg;
reg   [15:0] tmp_48_i_i_reg_650_pp0_iter14_reg;
reg   [15:0] tmp_48_i_i_reg_650_pp0_iter15_reg;
wire   [15:0] grp_fu_227_p2;
reg   [15:0] sub_i_i_i_reg_655;
wire   [15:0] grp_fu_231_p2;
reg   [15:0] normalized_reg_665;
wire   [15:0] grp_fu_223_p2;
reg   [15:0] biased_reg_675;
reg    ap_block_state1;
wire    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_exit_iter0_state2;
reg    ap_enable_reg_pp0_iter2;
reg    ap_enable_reg_pp0_iter3;
reg    ap_enable_reg_pp0_iter4;
reg    ap_enable_reg_pp0_iter5;
reg    ap_enable_reg_pp0_iter6;
reg    ap_enable_reg_pp0_iter7;
reg    ap_enable_reg_pp0_iter8;
reg    ap_enable_reg_pp0_iter9;
reg    ap_enable_reg_pp0_iter10;
reg    ap_enable_reg_pp0_iter11;
reg    ap_enable_reg_pp0_iter12;
reg    ap_enable_reg_pp0_iter13;
reg    ap_enable_reg_pp0_iter14;
reg    ap_enable_reg_pp0_iter15;
reg    ap_enable_reg_pp0_iter16;
reg    ap_enable_reg_pp0_iter17;
reg    ap_enable_reg_pp0_iter18;
reg    ap_enable_reg_pp0_iter19;
reg    ap_enable_reg_pp0_iter20;
reg    ap_enable_reg_pp0_iter21;
reg    ap_enable_reg_pp0_iter22;
wire    ap_block_pp0_stage0;
wire   [63:0] sext_ln109_fu_509_p1;
reg   [15:0] quad_3_14_fu_114;
wire   [15:0] quad_3_26_fu_475_p3;
reg   [15:0] quad_3_15_fu_118;
wire   [15:0] quad_3_25_fu_467_p3;
reg   [15:0] quad_3_16_fu_122;
wire   [15:0] quad_3_23_fu_451_p3;
reg   [15:0] quad_3_17_fu_126;
wire   [15:0] quad_3_20_fu_427_p3;
wire   [15:0] grp_fu_223_p1;
wire   [15:0] grp_fu_227_p1;
wire   [15:0] grp_fu_231_p1;
wire   [11:0] tmp_fu_235_p3;
wire   [8:0] tmp_s_fu_247_p3;
wire   [12:0] zext_ln109_fu_243_p1;
wire   [12:0] zext_ln109_3_fu_255_p1;
wire   [12:0] sub_ln109_fu_259_p2;
wire   [13:0] sub_ln109_cast_fu_265_p1;
wire   [13:0] zext_ln109_4_fu_269_p1;
wire   [0:0] icmp_ln103_fu_301_p2;
wire   [15:0] trunc_ln95_fu_329_p1;
wire   [15:0] data_V_fu_378_p1;
wire   [0:0] p_Result_s_fu_381_p3;
wire   [0:0] icmp_ln99_fu_396_p2;
wire   [15:0] quad_0_fu_389_p3;
wire   [0:0] icmp_ln99_3_fu_409_p2;
wire   [15:0] quad_3_fu_401_p3;
wire   [0:0] icmp_ln99_4_fu_422_p2;
wire   [15:0] quad_3_19_fu_414_p3;
wire   [15:0] quad_3_21_fu_435_p3;
wire   [15:0] quad_3_22_fu_443_p3;
wire   [15:0] quad_3_24_fu_459_p3;
wire   [15:0] tmp_34_fu_503_p3;
wire   [15:0] bitcast_ln109_6_fu_526_p1;
wire   [15:0] bitcast_ln109_5_fu_522_p1;
wire   [15:0] bitcast_ln109_4_fu_518_p1;
wire   [15:0] bitcast_ln109_fu_514_p1;
wire    ap_CS_fsm_state25;
reg   [2:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
#0 ap_enable_reg_pp0_iter4 = 1'b0;
#0 ap_enable_reg_pp0_iter5 = 1'b0;
#0 ap_enable_reg_pp0_iter6 = 1'b0;
#0 ap_enable_reg_pp0_iter7 = 1'b0;
#0 ap_enable_reg_pp0_iter8 = 1'b0;
#0 ap_enable_reg_pp0_iter9 = 1'b0;
#0 ap_enable_reg_pp0_iter10 = 1'b0;
#0 ap_enable_reg_pp0_iter11 = 1'b0;
#0 ap_enable_reg_pp0_iter12 = 1'b0;
#0 ap_enable_reg_pp0_iter13 = 1'b0;
#0 ap_enable_reg_pp0_iter14 = 1'b0;
#0 ap_enable_reg_pp0_iter15 = 1'b0;
#0 ap_enable_reg_pp0_iter16 = 1'b0;
#0 ap_enable_reg_pp0_iter17 = 1'b0;
#0 ap_enable_reg_pp0_iter18 = 1'b0;
#0 ap_enable_reg_pp0_iter19 = 1'b0;
#0 ap_enable_reg_pp0_iter20 = 1'b0;
#0 ap_enable_reg_pp0_iter21 = 1'b0;
#0 ap_enable_reg_pp0_iter22 = 1'b0;
end

td_fused_top_tdf4_l2_writeOutputs_133_running_sums_1 #(
    .DataWidth( 16 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
running_sums_1_U(
    .reset(ap_rst),
    .clk(ap_clk),
    .address0(running_sums_1_addr_reg_597_pp0_iter6_reg),
    .ce0(running_sums_1_ce0),
    .we0(running_sums_1_we0),
    .d0(running_sums_1_d0),
    .address1(running_sums_1_address1),
    .ce1(running_sums_1_ce1),
    .q1(running_sums_1_q1)
);

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U240(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(running_sums_1_load_reg_624),
    .din1(val_reg_619),
    .dout(grp_fu_219_p2)
);

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U241(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(normalized_reg_665),
    .din1(grp_fu_223_p1),
    .dout(grp_fu_223_p2)
);

td_fused_top_hsub_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hsub_16ns_16ns_16_5_full_dsp_1_U242(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(sum_reg_634),
    .din1(grp_fu_227_p1),
    .dout(grp_fu_227_p2)
);

td_fused_top_hmul_16ns_16ns_16_4_max_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hmul_16ns_16ns_16_4_max_dsp_1_U243(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(sub_i_i_i_reg_655),
    .din1(grp_fu_231_p1),
    .dout(grp_fu_231_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state25)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b1 == ap_condition_pp0_exit_iter0_state2) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((~((ap_start == 1'b0) | (write4_empty_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            if ((1'b1 == ap_condition_pp0_exit_iter0_state2)) begin
                ap_enable_reg_pp0_iter1 <= (1'b1 ^ ap_condition_pp0_exit_iter0_state2);
            end else if ((1'b1 == 1'b1)) begin
                ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
            end
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter10 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter10 <= ap_enable_reg_pp0_iter9;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter11 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter11 <= ap_enable_reg_pp0_iter10;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter12 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter12 <= ap_enable_reg_pp0_iter11;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter13 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter13 <= ap_enable_reg_pp0_iter12;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter14 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter14 <= ap_enable_reg_pp0_iter13;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter15 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter15 <= ap_enable_reg_pp0_iter14;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter16 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter16 <= ap_enable_reg_pp0_iter15;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter17 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter17 <= ap_enable_reg_pp0_iter16;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter18 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter18 <= ap_enable_reg_pp0_iter17;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter19 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter19 <= ap_enable_reg_pp0_iter18;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter20 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter20 <= ap_enable_reg_pp0_iter19;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter21 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter21 <= ap_enable_reg_pp0_iter20;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter22 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter22 <= ap_enable_reg_pp0_iter21;
        end else if ((~((ap_start == 1'b0) | (write4_empty_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter22 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter4 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter5 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter5 <= ap_enable_reg_pp0_iter4;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter6 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter6 <= ap_enable_reg_pp0_iter5;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter7 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter7 <= ap_enable_reg_pp0_iter6;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter8 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter8 <= ap_enable_reg_pp0_iter7;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter9 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter9 <= ap_enable_reg_pp0_iter8;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (icmp_ln86_fu_285_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        ochan_reg_208 <= add_ln86_fu_279_p2;
    end else if ((~((ap_start == 1'b0) | (write4_empty_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ochan_reg_208 <= 5'd0;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state1)) begin
        add_ln109_reg_573 <= add_ln109_fu_273_p2;
        write4_read_reg_567 <= write4_dout;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (icmp_ln86_fu_285_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        and_ln103_reg_610 <= and_ln103_fu_307_p2;
        running_sums_1_addr_reg_597 <= zext_ln86_fu_291_p1;
        trunc_ln99_reg_603 <= trunc_ln99_fu_297_p1;
        zext_ln86_reg_587[4 : 0] <= zext_ln86_fu_291_p1[4 : 0];
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        and_ln103_reg_610_pp0_iter10_reg <= and_ln103_reg_610_pp0_iter9_reg;
        and_ln103_reg_610_pp0_iter11_reg <= and_ln103_reg_610_pp0_iter10_reg;
        and_ln103_reg_610_pp0_iter12_reg <= and_ln103_reg_610_pp0_iter11_reg;
        and_ln103_reg_610_pp0_iter13_reg <= and_ln103_reg_610_pp0_iter12_reg;
        and_ln103_reg_610_pp0_iter14_reg <= and_ln103_reg_610_pp0_iter13_reg;
        and_ln103_reg_610_pp0_iter15_reg <= and_ln103_reg_610_pp0_iter14_reg;
        and_ln103_reg_610_pp0_iter16_reg <= and_ln103_reg_610_pp0_iter15_reg;
        and_ln103_reg_610_pp0_iter17_reg <= and_ln103_reg_610_pp0_iter16_reg;
        and_ln103_reg_610_pp0_iter18_reg <= and_ln103_reg_610_pp0_iter17_reg;
        and_ln103_reg_610_pp0_iter19_reg <= and_ln103_reg_610_pp0_iter18_reg;
        and_ln103_reg_610_pp0_iter20_reg <= and_ln103_reg_610_pp0_iter19_reg;
        and_ln103_reg_610_pp0_iter2_reg <= and_ln103_reg_610_pp0_iter1_reg;
        and_ln103_reg_610_pp0_iter3_reg <= and_ln103_reg_610_pp0_iter2_reg;
        and_ln103_reg_610_pp0_iter4_reg <= and_ln103_reg_610_pp0_iter3_reg;
        and_ln103_reg_610_pp0_iter5_reg <= and_ln103_reg_610_pp0_iter4_reg;
        and_ln103_reg_610_pp0_iter6_reg <= and_ln103_reg_610_pp0_iter5_reg;
        and_ln103_reg_610_pp0_iter7_reg <= and_ln103_reg_610_pp0_iter6_reg;
        and_ln103_reg_610_pp0_iter8_reg <= and_ln103_reg_610_pp0_iter7_reg;
        and_ln103_reg_610_pp0_iter9_reg <= and_ln103_reg_610_pp0_iter8_reg;
        biased_reg_675 <= grp_fu_223_p2;
        lshr_ln_reg_614_pp0_iter10_reg <= lshr_ln_reg_614_pp0_iter9_reg;
        lshr_ln_reg_614_pp0_iter11_reg <= lshr_ln_reg_614_pp0_iter10_reg;
        lshr_ln_reg_614_pp0_iter12_reg <= lshr_ln_reg_614_pp0_iter11_reg;
        lshr_ln_reg_614_pp0_iter13_reg <= lshr_ln_reg_614_pp0_iter12_reg;
        lshr_ln_reg_614_pp0_iter14_reg <= lshr_ln_reg_614_pp0_iter13_reg;
        lshr_ln_reg_614_pp0_iter15_reg <= lshr_ln_reg_614_pp0_iter14_reg;
        lshr_ln_reg_614_pp0_iter16_reg <= lshr_ln_reg_614_pp0_iter15_reg;
        lshr_ln_reg_614_pp0_iter17_reg <= lshr_ln_reg_614_pp0_iter16_reg;
        lshr_ln_reg_614_pp0_iter18_reg <= lshr_ln_reg_614_pp0_iter17_reg;
        lshr_ln_reg_614_pp0_iter19_reg <= lshr_ln_reg_614_pp0_iter18_reg;
        lshr_ln_reg_614_pp0_iter20_reg <= lshr_ln_reg_614_pp0_iter19_reg;
        lshr_ln_reg_614_pp0_iter2_reg <= lshr_ln_reg_614_pp0_iter1_reg;
        lshr_ln_reg_614_pp0_iter3_reg <= lshr_ln_reg_614_pp0_iter2_reg;
        lshr_ln_reg_614_pp0_iter4_reg <= lshr_ln_reg_614_pp0_iter3_reg;
        lshr_ln_reg_614_pp0_iter5_reg <= lshr_ln_reg_614_pp0_iter4_reg;
        lshr_ln_reg_614_pp0_iter6_reg <= lshr_ln_reg_614_pp0_iter5_reg;
        lshr_ln_reg_614_pp0_iter7_reg <= lshr_ln_reg_614_pp0_iter6_reg;
        lshr_ln_reg_614_pp0_iter8_reg <= lshr_ln_reg_614_pp0_iter7_reg;
        lshr_ln_reg_614_pp0_iter9_reg <= lshr_ln_reg_614_pp0_iter8_reg;
        normalized_reg_665 <= grp_fu_231_p2;
        running_sums_1_addr_reg_597_pp0_iter2_reg <= running_sums_1_addr_reg_597_pp0_iter1_reg;
        running_sums_1_addr_reg_597_pp0_iter3_reg <= running_sums_1_addr_reg_597_pp0_iter2_reg;
        running_sums_1_addr_reg_597_pp0_iter4_reg <= running_sums_1_addr_reg_597_pp0_iter3_reg;
        running_sums_1_addr_reg_597_pp0_iter5_reg <= running_sums_1_addr_reg_597_pp0_iter4_reg;
        running_sums_1_addr_reg_597_pp0_iter6_reg <= running_sums_1_addr_reg_597_pp0_iter5_reg;
        sub_i_i_i_reg_655 <= grp_fu_227_p2;
        sum_reg_634 <= grp_fu_219_p2;
        tmp_47_i_i_reg_645 <= {{l2_adjustments_q0[31:16]}};
        tmp_47_i_i_reg_645_pp0_iter10_reg <= tmp_47_i_i_reg_645_pp0_iter9_reg;
        tmp_47_i_i_reg_645_pp0_iter11_reg <= tmp_47_i_i_reg_645_pp0_iter10_reg;
        tmp_47_i_i_reg_645_pp0_iter8_reg <= tmp_47_i_i_reg_645;
        tmp_47_i_i_reg_645_pp0_iter9_reg <= tmp_47_i_i_reg_645_pp0_iter8_reg;
        tmp_48_i_i_reg_650 <= {{l2_adjustments_q0[47:32]}};
        tmp_48_i_i_reg_650_pp0_iter10_reg <= tmp_48_i_i_reg_650_pp0_iter9_reg;
        tmp_48_i_i_reg_650_pp0_iter11_reg <= tmp_48_i_i_reg_650_pp0_iter10_reg;
        tmp_48_i_i_reg_650_pp0_iter12_reg <= tmp_48_i_i_reg_650_pp0_iter11_reg;
        tmp_48_i_i_reg_650_pp0_iter13_reg <= tmp_48_i_i_reg_650_pp0_iter12_reg;
        tmp_48_i_i_reg_650_pp0_iter14_reg <= tmp_48_i_i_reg_650_pp0_iter13_reg;
        tmp_48_i_i_reg_650_pp0_iter15_reg <= tmp_48_i_i_reg_650_pp0_iter14_reg;
        tmp_48_i_i_reg_650_pp0_iter8_reg <= tmp_48_i_i_reg_650;
        tmp_48_i_i_reg_650_pp0_iter9_reg <= tmp_48_i_i_reg_650_pp0_iter8_reg;
        trunc_ln99_reg_603_pp0_iter10_reg <= trunc_ln99_reg_603_pp0_iter9_reg;
        trunc_ln99_reg_603_pp0_iter11_reg <= trunc_ln99_reg_603_pp0_iter10_reg;
        trunc_ln99_reg_603_pp0_iter12_reg <= trunc_ln99_reg_603_pp0_iter11_reg;
        trunc_ln99_reg_603_pp0_iter13_reg <= trunc_ln99_reg_603_pp0_iter12_reg;
        trunc_ln99_reg_603_pp0_iter14_reg <= trunc_ln99_reg_603_pp0_iter13_reg;
        trunc_ln99_reg_603_pp0_iter15_reg <= trunc_ln99_reg_603_pp0_iter14_reg;
        trunc_ln99_reg_603_pp0_iter16_reg <= trunc_ln99_reg_603_pp0_iter15_reg;
        trunc_ln99_reg_603_pp0_iter17_reg <= trunc_ln99_reg_603_pp0_iter16_reg;
        trunc_ln99_reg_603_pp0_iter18_reg <= trunc_ln99_reg_603_pp0_iter17_reg;
        trunc_ln99_reg_603_pp0_iter19_reg <= trunc_ln99_reg_603_pp0_iter18_reg;
        trunc_ln99_reg_603_pp0_iter20_reg <= trunc_ln99_reg_603_pp0_iter19_reg;
        trunc_ln99_reg_603_pp0_iter2_reg <= trunc_ln99_reg_603_pp0_iter1_reg;
        trunc_ln99_reg_603_pp0_iter3_reg <= trunc_ln99_reg_603_pp0_iter2_reg;
        trunc_ln99_reg_603_pp0_iter4_reg <= trunc_ln99_reg_603_pp0_iter3_reg;
        trunc_ln99_reg_603_pp0_iter5_reg <= trunc_ln99_reg_603_pp0_iter4_reg;
        trunc_ln99_reg_603_pp0_iter6_reg <= trunc_ln99_reg_603_pp0_iter5_reg;
        trunc_ln99_reg_603_pp0_iter7_reg <= trunc_ln99_reg_603_pp0_iter6_reg;
        trunc_ln99_reg_603_pp0_iter8_reg <= trunc_ln99_reg_603_pp0_iter7_reg;
        trunc_ln99_reg_603_pp0_iter9_reg <= trunc_ln99_reg_603_pp0_iter8_reg;
        zext_ln86_reg_587_pp0_iter2_reg[4 : 0] <= zext_ln86_reg_587_pp0_iter1_reg[4 : 0];
        zext_ln86_reg_587_pp0_iter3_reg[4 : 0] <= zext_ln86_reg_587_pp0_iter2_reg[4 : 0];
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        and_ln103_reg_610_pp0_iter1_reg <= and_ln103_reg_610;
        lshr_ln_reg_614_pp0_iter1_reg <= lshr_ln_reg_614;
        running_sums_1_addr_reg_597_pp0_iter1_reg <= running_sums_1_addr_reg_597;
        trunc_ln99_reg_603_pp0_iter1_reg <= trunc_ln99_reg_603;
        val_reg_619 <= l2_partial_sums_q0;
        zext_ln86_reg_587_pp0_iter1_reg[4 : 0] <= zext_ln86_reg_587[4 : 0];
    end
end

always @ (posedge ap_clk) begin
    if (((1'd1 == and_ln103_fu_307_p2) & (1'b1 == ap_CS_fsm_pp0_stage0) & (icmp_ln86_fu_285_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        lshr_ln_reg_614 <= {{ochan_reg_208[3:2]}};
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        quad_3_14_fu_114 <= quad_3_26_fu_475_p3;
        quad_3_15_fu_118 <= quad_3_25_fu_467_p3;
        quad_3_16_fu_122 <= quad_3_23_fu_451_p3;
        quad_3_17_fu_126 <= quad_3_20_fu_427_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        running_sums_1_load_reg_624 <= running_sums_1_q1;
    end
end

always @ (*) begin
    if ((icmp_ln86_fu_285_p2 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state2 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state2 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state25)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter22 == 1'b0) & (ap_enable_reg_pp0_iter21 == 1'b0) & (ap_enable_reg_pp0_iter20 == 1'b0) & (ap_enable_reg_pp0_iter19 == 1'b0) & (ap_enable_reg_pp0_iter18 == 1'b0) & (ap_enable_reg_pp0_iter17 == 1'b0) & (ap_enable_reg_pp0_iter16 == 1'b0) & (ap_enable_reg_pp0_iter15 == 1'b0) & (ap_enable_reg_pp0_iter14 == 1'b0) & (ap_enable_reg_pp0_iter13 == 1'b0) & (ap_enable_reg_pp0_iter12 == 1'b0) & (ap_enable_reg_pp0_iter11 == 1'b0) & (ap_enable_reg_pp0_iter10 == 1'b0) & (ap_enable_reg_pp0_iter9 == 1'b0) & (ap_enable_reg_pp0_iter8 == 1'b0) & (ap_enable_reg_pp0_iter7 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state25)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_01_blk_n = indices_01_empty_n;
    end else begin
        indices_01_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (write4_empty_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_01_read = 1'b1;
    end else begin
        indices_01_read = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_12_blk_n = indices_12_empty_n;
    end else begin
        indices_12_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (write4_empty_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_12_read = 1'b1;
    end else begin
        indices_12_read = 1'b0;
    end
end

always @ (*) begin
    if ((((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001)) | ((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001)) | ((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001)) | ((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
        l2_adjustments_ce0 = 1'b1;
    end else begin
        l2_adjustments_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        l2_partial_sums_ce0 = 1'b1;
    end else begin
        l2_partial_sums_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001)) | ((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
        out_data_ce1 = 1'b1;
    end else begin
        out_data_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'd1 == and_ln103_reg_610_pp0_iter20_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        out_data_we1 = 1'b1;
    end else begin
        out_data_we1 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        running_sums_1_ce0 = 1'b1;
    end else begin
        running_sums_1_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        running_sums_1_ce1 = 1'b1;
    end else begin
        running_sums_1_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        running_sums_1_we0 = 1'b1;
    end else begin
        running_sums_1_we0 = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        write4_blk_n = write4_empty_n;
    end else begin
        write4_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (write4_empty_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        write4_read = 1'b1;
    end else begin
        write4_read = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_start == 1'b0) | (write4_empty_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((~((ap_enable_reg_pp0_iter0 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0) & (icmp_ln86_fu_285_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone)) & ~((ap_enable_reg_pp0_iter22 == 1'b1) & (ap_enable_reg_pp0_iter21 == 1'b0) & (1'b0 == ap_block_pp0_stage0_subdone)))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0) & (icmp_ln86_fu_285_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone)) | ((ap_enable_reg_pp0_iter22 == 1'b1) & (ap_enable_reg_pp0_iter21 == 1'b0) & (1'b0 == ap_block_pp0_stage0_subdone)))) begin
                ap_NS_fsm = ap_ST_fsm_state25;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state25 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln109_fu_273_p2 = ((sub_ln109_cast_fu_265_p1) + (zext_ln109_4_fu_269_p1));

assign add_ln86_fu_279_p2 = (ochan_reg_208 + 5'd1);

assign and_ln103_fu_307_p2 = (write4_read_reg_567 & icmp_ln103_fu_301_p2);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state25 = ap_CS_fsm[32'd2];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (write4_empty_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1));
end

assign ap_block_state10_pp0_stage0_iter8 = ~(1'b1 == 1'b1);

assign ap_block_state11_pp0_stage0_iter9 = ~(1'b1 == 1'b1);

assign ap_block_state12_pp0_stage0_iter10 = ~(1'b1 == 1'b1);

assign ap_block_state13_pp0_stage0_iter11 = ~(1'b1 == 1'b1);

assign ap_block_state14_pp0_stage0_iter12 = ~(1'b1 == 1'b1);

assign ap_block_state15_pp0_stage0_iter13 = ~(1'b1 == 1'b1);

assign ap_block_state16_pp0_stage0_iter14 = ~(1'b1 == 1'b1);

assign ap_block_state17_pp0_stage0_iter15 = ~(1'b1 == 1'b1);

assign ap_block_state18_pp0_stage0_iter16 = ~(1'b1 == 1'b1);

assign ap_block_state19_pp0_stage0_iter17 = ~(1'b1 == 1'b1);

assign ap_block_state20_pp0_stage0_iter18 = ~(1'b1 == 1'b1);

assign ap_block_state21_pp0_stage0_iter19 = ~(1'b1 == 1'b1);

assign ap_block_state22_pp0_stage0_iter20 = ~(1'b1 == 1'b1);

assign ap_block_state23_pp0_stage0_iter21 = ~(1'b1 == 1'b1);

assign ap_block_state24_pp0_stage0_iter22 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter4 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage0_iter5 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage0_iter6 = ~(1'b1 == 1'b1);

assign ap_block_state9_pp0_stage0_iter7 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign bitcast_ln109_4_fu_518_p1 = quad_3_25_fu_467_p3;

assign bitcast_ln109_5_fu_522_p1 = quad_3_23_fu_451_p3;

assign bitcast_ln109_6_fu_526_p1 = quad_3_20_fu_427_p3;

assign bitcast_ln109_fu_514_p1 = quad_3_26_fu_475_p3;

assign data_V_fu_378_p1 = biased_reg_675;

assign grp_fu_223_p1 = tmp_48_i_i_reg_650_pp0_iter15_reg;

assign grp_fu_227_p1 = trunc_ln95_fu_329_p1;

assign grp_fu_231_p1 = tmp_47_i_i_reg_645_pp0_iter11_reg;

assign icmp_ln103_fu_301_p2 = ((trunc_ln99_fu_297_p1 == 2'd3) ? 1'b1 : 1'b0);

assign icmp_ln86_fu_285_p2 = ((ochan_reg_208 == 5'd16) ? 1'b1 : 1'b0);

assign icmp_ln99_3_fu_409_p2 = ((trunc_ln99_reg_603_pp0_iter20_reg == 2'd1) ? 1'b1 : 1'b0);

assign icmp_ln99_4_fu_422_p2 = ((trunc_ln99_reg_603_pp0_iter20_reg == 2'd0) ? 1'b1 : 1'b0);

assign icmp_ln99_fu_396_p2 = ((trunc_ln99_reg_603_pp0_iter20_reg == 2'd2) ? 1'b1 : 1'b0);

assign l2_adjustments_address0 = zext_ln86_reg_587_pp0_iter3_reg;

assign l2_partial_sums_address0 = zext_ln86_fu_291_p1;

assign out_data_address1 = sext_ln109_fu_509_p1;

assign out_data_d1 = {{{{bitcast_ln109_6_fu_526_p1}, {bitcast_ln109_5_fu_522_p1}}, {bitcast_ln109_4_fu_518_p1}}, {bitcast_ln109_fu_514_p1}};

assign p_Result_s_fu_381_p3 = data_V_fu_378_p1[32'd15];

assign quad_0_fu_389_p3 = ((p_Result_s_fu_381_p3[0:0] == 1'b1) ? 16'd0 : biased_reg_675);

assign quad_3_19_fu_414_p3 = ((icmp_ln99_3_fu_409_p2[0:0] == 1'b1) ? quad_3_17_fu_126 : quad_3_fu_401_p3);

assign quad_3_20_fu_427_p3 = ((icmp_ln99_4_fu_422_p2[0:0] == 1'b1) ? quad_3_17_fu_126 : quad_3_19_fu_414_p3);

assign quad_3_21_fu_435_p3 = ((icmp_ln99_fu_396_p2[0:0] == 1'b1) ? quad_0_fu_389_p3 : quad_3_16_fu_122);

assign quad_3_22_fu_443_p3 = ((icmp_ln99_3_fu_409_p2[0:0] == 1'b1) ? quad_3_16_fu_122 : quad_3_21_fu_435_p3);

assign quad_3_23_fu_451_p3 = ((icmp_ln99_4_fu_422_p2[0:0] == 1'b1) ? quad_3_16_fu_122 : quad_3_22_fu_443_p3);

assign quad_3_24_fu_459_p3 = ((icmp_ln99_3_fu_409_p2[0:0] == 1'b1) ? quad_0_fu_389_p3 : quad_3_15_fu_118);

assign quad_3_25_fu_467_p3 = ((icmp_ln99_4_fu_422_p2[0:0] == 1'b1) ? quad_3_15_fu_118 : quad_3_24_fu_459_p3);

assign quad_3_26_fu_475_p3 = ((icmp_ln99_4_fu_422_p2[0:0] == 1'b1) ? quad_0_fu_389_p3 : quad_3_14_fu_114);

assign quad_3_fu_401_p3 = ((icmp_ln99_fu_396_p2[0:0] == 1'b1) ? quad_3_17_fu_126 : quad_0_fu_389_p3);

assign running_sums_1_address1 = zext_ln86_fu_291_p1;

assign running_sums_1_d0 = ((write4_read_reg_567[0:0] == 1'b1) ? 16'd0 : sum_reg_634);

assign sext_ln109_fu_509_p1 = (tmp_34_fu_503_p3);

assign sub_ln109_cast_fu_265_p1 = (sub_ln109_fu_259_p2);

assign sub_ln109_fu_259_p2 = (zext_ln109_fu_243_p1 - zext_ln109_3_fu_255_p1);

assign tmp_34_fu_503_p3 = {{add_ln109_reg_573}, {lshr_ln_reg_614_pp0_iter20_reg}};

assign tmp_fu_235_p3 = {{indices_01_dout}, {6'd0}};

assign tmp_s_fu_247_p3 = {{indices_01_dout}, {3'd0}};

assign trunc_ln95_fu_329_p1 = l2_adjustments_q0[15:0];

assign trunc_ln99_fu_297_p1 = ochan_reg_208[1:0];

assign zext_ln109_3_fu_255_p1 = tmp_s_fu_247_p3;

assign zext_ln109_4_fu_269_p1 = indices_12_dout;

assign zext_ln109_fu_243_p1 = tmp_fu_235_p3;

assign zext_ln86_fu_291_p1 = ochan_reg_208;

always @ (posedge ap_clk) begin
    zext_ln86_reg_587[63:5] <= 59'b00000000000000000000000000000000000000000000000000000000000;
    zext_ln86_reg_587_pp0_iter1_reg[63:5] <= 59'b00000000000000000000000000000000000000000000000000000000000;
    zext_ln86_reg_587_pp0_iter2_reg[63:5] <= 59'b00000000000000000000000000000000000000000000000000000000000;
    zext_ln86_reg_587_pp0_iter3_reg[63:5] <= 59'b00000000000000000000000000000000000000000000000000000000000;
end

endmodule //td_fused_top_tdf4_l2_writeOutputs_133
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf4_readFilters36 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        filter_data_address0,
        filter_data_ce0,
        filter_data_q0,
        indices_23_dout,
        indices_23_empty_n,
        indices_23_read,
        weight_vecs_0_address0,
        weight_vecs_0_ce0,
        weight_vecs_0_we0,
        weight_vecs_0_d0
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state7 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [14:0] filter_data_address0;
output   filter_data_ce0;
input  [15:0] filter_data_q0;
input  [6:0] indices_23_dout;
input   indices_23_empty_n;
output   indices_23_read;
output  [7:0] weight_vecs_0_address0;
output   weight_vecs_0_ce0;
output   weight_vecs_0_we0;
output  [15:0] weight_vecs_0_d0;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg filter_data_ce0;
reg indices_23_read;
reg weight_vecs_0_ce0;
reg weight_vecs_0_we0;

reg    ap_done_reg;
  reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    indices_23_blk_n;
reg   [7:0] indvar_flatten13_reg_123;
reg   [1:0] ii_reg_134;
reg   [6:0] indvar_flatten_reg_145;
reg   [1:0] jj_reg_156;
reg   [4:0] kk_reg_167;
wire   [10:0] sext_ln47_fu_200_p1;
reg   [10:0] sext_ln47_reg_408;
wire   [7:0] add_ln47_4_fu_204_p2;
wire    ap_CS_fsm_pp0_stage0;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
wire    ap_block_state4_pp0_stage0_iter2;
wire    ap_block_state5_pp0_stage0_iter3;
wire    ap_block_state6_pp0_stage0_iter4;
wire    ap_block_pp0_stage0_11001;
wire   [0:0] icmp_ln47_fu_210_p2;
reg   [0:0] icmp_ln47_reg_418;
reg   [0:0] icmp_ln47_reg_418_pp0_iter1_reg;
reg   [0:0] icmp_ln47_reg_418_pp0_iter2_reg;
reg   [0:0] icmp_ln47_reg_418_pp0_iter3_reg;
wire   [0:0] icmp_ln48_fu_222_p2;
reg   [0:0] icmp_ln48_reg_422;
wire   [1:0] select_ln47_4_fu_228_p3;
reg   [1:0] select_ln47_4_reg_429;
wire   [6:0] select_ln48_8_fu_242_p3;
wire   [1:0] select_ln48_7_fu_329_p3;
reg   [1:0] select_ln48_7_reg_442;
reg    ap_enable_reg_pp0_iter1;
wire   [7:0] add_ln55_16_fu_392_p2;
reg   [7:0] add_ln55_16_reg_452;
reg   [7:0] add_ln55_16_reg_452_pp0_iter2_reg;
reg   [7:0] add_ln55_16_reg_452_pp0_iter3_reg;
wire   [4:0] add_ln49_fu_398_p2;
reg    ap_block_state1;
wire    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_flush_enable;
reg    ap_enable_reg_pp0_iter2;
reg    ap_condition_pp0_exit_iter1_state3;
reg    ap_enable_reg_pp0_iter3;
reg    ap_enable_reg_pp0_iter4;
reg   [1:0] ap_phi_mux_ii_phi_fu_138_p4;
wire    ap_block_pp0_stage0;
reg   [1:0] ap_phi_mux_jj_phi_fu_160_p4;
wire   [63:0] zext_ln55_37_fu_387_p1;
wire   [63:0] zext_ln55_38_fu_404_p1;
wire   [8:0] tmp_fu_182_p3;
wire   [9:0] zext_ln55_30_fu_190_p1;
wire   [9:0] zext_ln55_fu_178_p1;
wire   [9:0] sub_ln55_fu_194_p2;
wire   [1:0] add_ln47_fu_216_p2;
wire   [6:0] add_ln48_4_fu_236_p2;
wire   [10:0] zext_ln55_32_fu_260_p1;
wire   [10:0] add_ln55_fu_263_p2;
wire   [10:0] shl_ln55_fu_268_p2;
wire   [3:0] tmp_s_fu_280_p3;
wire   [3:0] zext_ln55_31_fu_257_p1;
wire   [0:0] icmp_ln49_fu_298_p2;
wire   [0:0] xor_ln47_fu_293_p2;
wire   [1:0] select_ln47_fu_250_p3;
wire   [0:0] and_ln47_fu_304_p2;
wire   [0:0] or_ln48_fu_316_p2;
wire   [1:0] add_ln48_fu_310_p2;
wire   [10:0] sub_ln55_7_fu_274_p2;
wire   [10:0] zext_ln55_34_fu_341_p1;
wire   [10:0] add_ln55_13_fu_345_p2;
wire   [3:0] sub_ln55_8_fu_287_p2;
wire   [3:0] zext_ln55_33_fu_337_p1;
wire   [3:0] add_ln55_14_fu_359_p2;
wire   [4:0] select_ln48_fu_321_p3;
wire   [14:0] tmp_91_cast_fu_351_p3;
wire   [14:0] zext_ln55_36_fu_377_p1;
wire   [14:0] add_ln55_15_fu_381_p2;
wire   [7:0] tmp_93_cast_fu_365_p3;
wire   [7:0] zext_ln55_35_fu_373_p1;
wire    ap_CS_fsm_state7;
reg   [2:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
#0 ap_enable_reg_pp0_iter4 = 1'b0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state7)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if ((1'b1 == ap_condition_pp0_flush_enable)) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            if ((1'b1 == ap_condition_pp0_exit_iter1_state3)) begin
                ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter0;
            end else if ((1'b1 == 1'b1)) begin
                ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
            end
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter4 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
        end else if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter4 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln47_reg_418 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ii_reg_134 <= select_ln47_4_reg_429;
    end else if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ii_reg_134 <= 2'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_fu_210_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        indvar_flatten13_reg_123 <= add_ln47_4_fu_204_p2;
    end else if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indvar_flatten13_reg_123 <= 8'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_fu_210_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        indvar_flatten_reg_145 <= select_ln48_8_fu_242_p3;
    end else if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indvar_flatten_reg_145 <= 7'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_reg_418_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        jj_reg_156 <= select_ln48_7_reg_442;
    end else if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        jj_reg_156 <= 2'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln47_reg_418 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        kk_reg_167 <= add_ln49_fu_398_p2;
    end else if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        kk_reg_167 <= 5'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_reg_418 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        add_ln55_16_reg_452 <= add_ln55_16_fu_392_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        add_ln55_16_reg_452_pp0_iter2_reg <= add_ln55_16_reg_452;
        add_ln55_16_reg_452_pp0_iter3_reg <= add_ln55_16_reg_452_pp0_iter2_reg;
        icmp_ln47_reg_418_pp0_iter2_reg <= icmp_ln47_reg_418_pp0_iter1_reg;
        icmp_ln47_reg_418_pp0_iter3_reg <= icmp_ln47_reg_418_pp0_iter2_reg;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln47_reg_418 <= icmp_ln47_fu_210_p2;
        icmp_ln47_reg_418_pp0_iter1_reg <= icmp_ln47_reg_418;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_fu_210_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln48_reg_422 <= icmp_ln48_fu_222_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_fu_210_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        select_ln47_4_reg_429 <= select_ln47_4_fu_228_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln47_reg_418 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        select_ln48_7_reg_442 <= select_ln48_7_fu_329_p3;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state1)) begin
        sext_ln47_reg_408 <= sext_ln47_fu_200_p1;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_condition_pp0_exit_iter1_state3 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter1_state3 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln47_fu_210_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_condition_pp0_flush_enable = 1'b1;
    end else begin
        ap_condition_pp0_flush_enable = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state7)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln47_reg_418 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_phi_mux_ii_phi_fu_138_p4 = select_ln47_4_reg_429;
    end else begin
        ap_phi_mux_ii_phi_fu_138_p4 = ii_reg_134;
    end
end

always @ (*) begin
    if (((icmp_ln47_reg_418_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        ap_phi_mux_jj_phi_fu_160_p4 = select_ln48_7_reg_442;
    end else begin
        ap_phi_mux_jj_phi_fu_160_p4 = jj_reg_156;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state7)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter3 == 1'b1)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter4 == 1'b1)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1)))) begin
        filter_data_ce0 = 1'b1;
    end else begin
        filter_data_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_23_blk_n = indices_23_empty_n;
    end else begin
        indices_23_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_23_read = 1'b1;
    end else begin
        indices_23_read = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter4 == 1'b1))) begin
        weight_vecs_0_ce0 = 1'b1;
    end else begin
        weight_vecs_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln47_reg_418_pp0_iter3_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter4 == 1'b1))) begin
        weight_vecs_0_we0 = 1'b1;
    end else begin
        weight_vecs_0_we0 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((~((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b0)) & ~((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter4 == 1'b1) & (ap_enable_reg_pp0_iter3 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if ((((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b0)) | ((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter4 == 1'b1) & (ap_enable_reg_pp0_iter3 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_state7;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state7 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln47_4_fu_204_p2 = (indvar_flatten13_reg_123 + 8'd1);

assign add_ln47_fu_216_p2 = (ap_phi_mux_ii_phi_fu_138_p4 + 2'd1);

assign add_ln48_4_fu_236_p2 = (indvar_flatten_reg_145 + 7'd1);

assign add_ln48_fu_310_p2 = (select_ln47_fu_250_p3 + 2'd1);

assign add_ln49_fu_398_p2 = (select_ln48_fu_321_p3 + 5'd1);

assign add_ln55_13_fu_345_p2 = (sub_ln55_7_fu_274_p2 + zext_ln55_34_fu_341_p1);

assign add_ln55_14_fu_359_p2 = (sub_ln55_8_fu_287_p2 + zext_ln55_33_fu_337_p1);

assign add_ln55_15_fu_381_p2 = (tmp_91_cast_fu_351_p3 + zext_ln55_36_fu_377_p1);

assign add_ln55_16_fu_392_p2 = (tmp_93_cast_fu_365_p3 + zext_ln55_35_fu_373_p1);

assign add_ln55_fu_263_p2 = ((sext_ln47_reg_408) + (zext_ln55_32_fu_260_p1));

assign and_ln47_fu_304_p2 = (xor_ln47_fu_293_p2 & icmp_ln49_fu_298_p2);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state7 = ap_CS_fsm[32'd2];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1));
end

assign ap_block_state2_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter4 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign filter_data_address0 = zext_ln55_37_fu_387_p1;

assign icmp_ln47_fu_210_p2 = ((indvar_flatten13_reg_123 == 8'd144) ? 1'b1 : 1'b0);

assign icmp_ln48_fu_222_p2 = ((indvar_flatten_reg_145 == 7'd48) ? 1'b1 : 1'b0);

assign icmp_ln49_fu_298_p2 = ((kk_reg_167 == 5'd16) ? 1'b1 : 1'b0);

assign or_ln48_fu_316_p2 = (icmp_ln48_reg_422 | and_ln47_fu_304_p2);

assign select_ln47_4_fu_228_p3 = ((icmp_ln48_fu_222_p2[0:0] == 1'b1) ? add_ln47_fu_216_p2 : ap_phi_mux_ii_phi_fu_138_p4);

assign select_ln47_fu_250_p3 = ((icmp_ln48_reg_422[0:0] == 1'b1) ? 2'd0 : ap_phi_mux_jj_phi_fu_160_p4);

assign select_ln48_7_fu_329_p3 = ((and_ln47_fu_304_p2[0:0] == 1'b1) ? add_ln48_fu_310_p2 : select_ln47_fu_250_p3);

assign select_ln48_8_fu_242_p3 = ((icmp_ln48_fu_222_p2[0:0] == 1'b1) ? 7'd1 : add_ln48_4_fu_236_p2);

assign select_ln48_fu_321_p3 = ((or_ln48_fu_316_p2[0:0] == 1'b1) ? 5'd0 : kk_reg_167);

assign sext_ln47_fu_200_p1 = (sub_ln55_fu_194_p2);

assign shl_ln55_fu_268_p2 = add_ln55_fu_263_p2 << 11'd2;

assign sub_ln55_7_fu_274_p2 = (shl_ln55_fu_268_p2 - add_ln55_fu_263_p2);

assign sub_ln55_8_fu_287_p2 = (tmp_s_fu_280_p3 - zext_ln55_31_fu_257_p1);

assign sub_ln55_fu_194_p2 = (zext_ln55_30_fu_190_p1 - zext_ln55_fu_178_p1);

assign tmp_91_cast_fu_351_p3 = {{add_ln55_13_fu_345_p2}, {4'd0}};

assign tmp_93_cast_fu_365_p3 = {{add_ln55_14_fu_359_p2}, {4'd0}};

assign tmp_fu_182_p3 = {{indices_23_dout}, {2'd0}};

assign tmp_s_fu_280_p3 = {{select_ln47_4_reg_429}, {2'd0}};

assign weight_vecs_0_address0 = zext_ln55_38_fu_404_p1;

assign weight_vecs_0_d0 = filter_data_q0;

assign xor_ln47_fu_293_p2 = (icmp_ln48_reg_422 ^ 1'd1);

assign zext_ln55_30_fu_190_p1 = tmp_fu_182_p3;

assign zext_ln55_31_fu_257_p1 = select_ln47_4_reg_429;

assign zext_ln55_32_fu_260_p1 = select_ln47_4_reg_429;

assign zext_ln55_33_fu_337_p1 = select_ln48_7_fu_329_p3;

assign zext_ln55_34_fu_341_p1 = select_ln48_7_fu_329_p3;

assign zext_ln55_35_fu_373_p1 = select_ln48_fu_321_p3;

assign zext_ln55_36_fu_377_p1 = select_ln48_fu_321_p3;

assign zext_ln55_37_fu_387_p1 = add_ln55_15_fu_381_p2;

assign zext_ln55_38_fu_404_p1 = add_ln55_16_reg_452_pp0_iter3_reg;

assign zext_ln55_fu_178_p1 = indices_23_dout;

endmodule //td_fused_top_tdf4_readFilters36
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf4_readInputs37 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        in_data_address0,
        in_data_ce0,
        in_data_q0,
        indices_01_dout,
        indices_01_empty_n,
        indices_01_read,
        indices_12_dout,
        indices_12_empty_n,
        indices_12_read,
        ifmap_vec_address0,
        ifmap_vec_ce0,
        ifmap_vec_we0,
        ifmap_vec_d0,
        ifmap_vec_address1,
        ifmap_vec_ce1,
        ifmap_vec_we1,
        ifmap_vec_d1,
        indices_01_out_din,
        indices_01_out_full_n,
        indices_01_out_write,
        indices_12_out_din,
        indices_12_out_full_n,
        indices_12_out_write
);

parameter    ap_ST_fsm_state1 = 5'd1;
parameter    ap_ST_fsm_state2 = 5'd2;
parameter    ap_ST_fsm_pp0_stage0 = 5'd4;
parameter    ap_ST_fsm_pp0_stage1 = 5'd8;
parameter    ap_ST_fsm_state9 = 5'd16;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [13:0] in_data_address0;
output   in_data_ce0;
input  [63:0] in_data_q0;
input  [15:0] indices_01_dout;
input   indices_01_empty_n;
output   indices_01_read;
input  [15:0] indices_12_dout;
input   indices_12_empty_n;
output   indices_12_read;
output  [7:0] ifmap_vec_address0;
output   ifmap_vec_ce0;
output   ifmap_vec_we0;
output  [15:0] ifmap_vec_d0;
output  [7:0] ifmap_vec_address1;
output   ifmap_vec_ce1;
output   ifmap_vec_we1;
output  [15:0] ifmap_vec_d1;
output  [5:0] indices_01_out_din;
input   indices_01_out_full_n;
output   indices_01_out_write;
output  [11:0] indices_12_out_din;
input   indices_12_out_full_n;
output   indices_12_out_write;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg in_data_ce0;
reg indices_01_read;
reg indices_12_read;
reg[7:0] ifmap_vec_address0;
reg ifmap_vec_ce0;
reg ifmap_vec_we0;
reg[15:0] ifmap_vec_d0;
reg[7:0] ifmap_vec_address1;
reg ifmap_vec_ce1;
reg ifmap_vec_we1;
reg[15:0] ifmap_vec_d1;
reg indices_01_out_write;
reg indices_12_out_write;

reg    ap_done_reg;
  reg   [4:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    indices_01_blk_n;
reg    indices_12_blk_n;
reg    indices_01_out_blk_n;
reg    indices_12_out_blk_n;
reg   [5:0] indvar_flatten47_reg_224;
reg   [1:0] ii_reg_236;
reg   [4:0] indvar_flatten_reg_248;
reg   [1:0] jj_reg_259;
reg   [4:0] kk_0_i_i_reg_271;
reg   [15:0] indices_01_read_reg_959;
wire   [5:0] trunc_ln250_fu_282_p1;
reg   [5:0] trunc_ln250_reg_964;
reg   [15:0] indices_12_read_reg_969;
wire   [11:0] empty_fu_287_p1;
reg   [11:0] empty_reg_974;
wire   [17:0] p_cast_i_i_fu_304_p1;
reg   [17:0] p_cast_i_i_reg_981;
wire    ap_CS_fsm_state2;
wire   [17:0] sext_ln22_fu_314_p1;
reg   [17:0] sext_ln22_reg_987;
wire   [5:0] p_cast_fu_318_p2;
reg   [5:0] p_cast_reg_993;
wire   [0:0] or_ln23_16_fu_337_p2;
reg   [0:0] or_ln23_16_reg_999;
wire   [11:0] p_mid137_fu_343_p2;
reg   [11:0] p_mid137_reg_1004;
wire   [5:0] p_cast5_i_i_fu_361_p2;
reg   [5:0] p_cast5_i_i_reg_1009;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_block_state3_pp0_stage0_iter0;
wire    ap_block_state5_pp0_stage0_iter1;
wire    ap_block_state7_pp0_stage0_iter2;
wire    ap_block_pp0_stage0_11001;
wire   [0:0] is_padding_fu_401_p2;
reg   [0:0] is_padding_reg_1015;
wire   [0:0] icmp_ln19_fu_407_p2;
reg   [0:0] icmp_ln19_reg_1022;
reg   [0:0] icmp_ln19_reg_1022_pp0_iter1_reg;
reg   [0:0] icmp_ln19_reg_1022_pp0_iter2_reg;
wire   [1:0] add_ln19_fu_413_p2;
reg   [1:0] add_ln19_reg_1026;
wire   [0:0] icmp_ln20_fu_419_p2;
reg   [0:0] icmp_ln20_reg_1031;
wire   [1:0] select_ln19_fu_425_p3;
reg   [1:0] select_ln19_reg_1043;
wire   [5:0] p_cast5_i_i_mid1_fu_446_p2;
reg   [5:0] p_cast5_i_i_mid1_reg_1048;
wire   [0:0] or_ln23_18_fu_465_p2;
reg   [0:0] or_ln23_18_reg_1054;
wire   [1:0] add_ln20_fu_470_p2;
reg   [1:0] add_ln20_reg_1061;
wire   [0:0] or_ln23_20_fu_505_p2;
reg   [0:0] or_ln23_20_reg_1067;
wire   [4:0] add_ln20_4_fu_511_p2;
reg   [4:0] add_ln20_4_reg_1074;
wire   [5:0] add_ln19_4_fu_517_p2;
reg   [5:0] add_ln19_4_reg_1079;
wire    ap_CS_fsm_pp0_stage1;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_state4_pp0_stage1_iter0;
wire    ap_block_state6_pp0_stage1_iter1;
wire    ap_block_state8_pp0_stage1_iter2;
wire    ap_block_pp0_stage1_11001;
wire   [1:0] select_ln19_19_fu_555_p3;
reg   [1:0] select_ln19_19_reg_1084;
wire   [4:0] select_ln20_fu_619_p3;
reg   [4:0] select_ln20_reg_1091;
wire   [1:0] select_ln20_16_fu_627_p3;
reg   [1:0] select_ln20_16_reg_1097;
wire   [0:0] select_ln20_17_fu_636_p3;
reg   [0:0] select_ln20_17_reg_1103;
reg   [0:0] select_ln20_17_reg_1103_pp0_iter1_reg;
wire   [3:0] empty_97_fu_732_p1;
reg   [3:0] empty_97_reg_1111;
reg   [3:0] empty_97_reg_1111_pp0_iter1_reg;
wire   [4:0] select_ln20_20_fu_759_p3;
reg   [4:0] select_ln20_20_reg_1123;
wire   [4:0] add_ln25_fu_765_p2;
reg   [4:0] add_ln25_reg_1128;
reg    ap_enable_reg_pp0_iter1;
wire   [5:0] add_ln33_fu_797_p2;
reg   [5:0] add_ln33_reg_1133;
wire   [7:0] add_ln33_4_fu_818_p2;
reg   [7:0] add_ln33_4_reg_1140;
wire   [15:0] select_ln33_17_fu_897_p3;
reg   [15:0] select_ln33_17_reg_1145;
wire   [15:0] select_ln33_18_fu_918_p3;
reg   [15:0] select_ln33_18_reg_1150;
wire    ap_block_pp0_stage1_subdone;
reg    ap_condition_pp0_exit_iter0_state4;
reg    ap_enable_reg_pp0_iter2;
reg   [5:0] ap_phi_mux_indvar_flatten47_phi_fu_228_p4;
wire    ap_block_pp0_stage0;
reg   [1:0] ap_phi_mux_ii_phi_fu_240_p4;
reg   [4:0] ap_phi_mux_indvar_flatten_phi_fu_252_p4;
reg   [1:0] ap_phi_mux_jj_phi_fu_263_p4;
reg   [4:0] ap_phi_mux_kk_0_i_i_phi_fu_275_p4;
wire    ap_block_pp0_stage1;
wire   [63:0] sext_ln32_fu_754_p1;
wire   [63:0] zext_ln33_17_fu_824_p1;
wire   [63:0] sext_ln33_fu_856_p1;
wire   [63:0] sext_ln33_7_fu_937_p1;
wire   [63:0] sext_ln33_8_fu_954_p1;
reg    ap_block_state1;
wire   [15:0] select_ln33_fu_836_p3;
wire   [15:0] select_ln33_16_fu_875_p3;
wire   [16:0] zext_ln19_fu_295_p1;
wire   [16:0] empty_92_fu_298_p2;
wire   [16:0] j_cast_i_i_fu_292_p1;
wire   [16:0] add_ln22_fu_308_p2;
wire   [0:0] tmp_26_fu_323_p3;
wire   [0:0] icmp_ln24_fu_331_p2;
wire   [17:0] ii_cast_i_i_fu_348_p1;
wire   [5:0] ii_cast_fu_352_p1;
wire   [17:0] empty_93_fu_356_p2;
wire   [17:0] zext_ln20_fu_372_p1;
wire   [17:0] add_ln22_4_fu_376_p2;
wire   [0:0] tmp_27_fu_381_p3;
wire   [0:0] icmp_ln24_4_fu_389_p2;
wire   [0:0] or_ln23_fu_395_p2;
wire   [0:0] empty_94_fu_366_p2;
wire   [17:0] ii_cast_i_i_mid1_fu_433_p1;
wire   [5:0] ii_cast_mid1_fu_437_p1;
wire   [17:0] p_mid111_fu_441_p2;
wire   [0:0] p_mid113_fu_451_p2;
wire   [17:0] zext_ln20_4_fu_476_p1;
wire   [17:0] add_ln22_5_fu_480_p2;
wire   [0:0] tmp_28_fu_485_p3;
wire   [0:0] icmp_ln24_5_fu_493_p2;
wire   [0:0] or_ln23_19_fu_499_p2;
wire   [0:0] select_ln19_21_fu_457_p3;
wire   [2:0] zext_ln22_fu_523_p1;
wire   [2:0] tmp1_fu_533_p2;
wire   [11:0] tmp1_cast_fu_539_p1;
wire   [11:0] empty_95_fu_543_p2;
wire   [5:0] row_coord_int_mid131_fu_571_p3;
wire   [5:0] row_coord_int_fu_527_p3;
wire   [11:0] col_coord_int_mid139_fu_577_p3;
wire   [11:0] col_coord_int_fu_548_p3;
wire   [0:0] icmp_ln25_fu_602_p2;
wire   [0:0] xor_ln19_fu_597_p2;
wire   [0:0] and_ln19_fu_608_p2;
wire   [0:0] or_ln20_fu_614_p2;
wire   [0:0] select_ln19_22_fu_566_p3;
wire   [5:0] select_ln19_20_fu_561_p3;
wire   [2:0] zext_ln22_4_fu_633_p1;
wire   [2:0] tmp1_mid1_fu_650_p2;
wire   [11:0] tmp1_cast_mid1_fu_656_p1;
wire   [11:0] p_mid1_fu_660_p2;
wire   [5:0] row_coord_int_mid1_fu_643_p3;
wire   [5:0] select_ln19_23_fu_583_p3;
wire   [5:0] select_ln20_18_fu_672_p3;
wire   [11:0] tmp_s_fu_680_p3;
wire   [8:0] tmp_6_fu_692_p3;
wire   [12:0] zext_ln32_fu_688_p1;
wire   [12:0] zext_ln32_18_fu_700_p1;
wire   [12:0] sub_ln32_fu_704_p2;
wire   [11:0] col_coord_int_mid1_fu_665_p3;
wire   [11:0] select_ln19_24_fu_590_p3;
wire   [11:0] select_ln20_19_fu_714_p3;
wire   [13:0] sext_ln20_fu_710_p1;
wire   [13:0] zext_ln32_19_fu_722_p1;
wire   [13:0] add_ln32_fu_726_p2;
wire   [1:0] lshr_ln_fu_736_p4;
wire   [15:0] tmp_29_fu_746_p3;
wire   [3:0] tmp_fu_773_p3;
wire   [4:0] zext_ln33_14_fu_780_p1;
wire   [4:0] zext_ln33_fu_770_p1;
wire   [4:0] sub_ln33_fu_784_p2;
wire   [5:0] sub_ln33_cast_fu_790_p1;
wire   [5:0] zext_ln33_15_fu_794_p1;
wire   [3:0] trunc_ln33_fu_803_p1;
wire   [7:0] tmp_80_cast_fu_807_p3;
wire   [7:0] zext_ln33_16_fu_815_p1;
wire   [15:0] trunc_ln32_fu_828_p1;
wire   [15:0] bitcast_ln32_fu_832_p1;
wire   [3:0] or_ln25_fu_844_p2;
wire   [9:0] tmp_30_fu_849_p3;
wire   [15:0] tmp_44_i_i_fu_861_p4;
wire   [15:0] bitcast_ln32_16_fu_871_p1;
wire   [15:0] tmp_45_i_i_fu_883_p4;
wire   [15:0] bitcast_ln32_17_fu_893_p1;
wire   [15:0] tmp_46_i_i_fu_904_p4;
wire   [15:0] bitcast_ln32_18_fu_914_p1;
wire   [3:0] or_ln25_11_fu_925_p2;
wire   [9:0] tmp_31_fu_930_p3;
wire   [3:0] or_ln25_12_fu_942_p2;
wire   [9:0] tmp_32_fu_947_p3;
wire    ap_CS_fsm_state9;
reg   [4:0] ap_NS_fsm;
wire    ap_block_pp0_stage0_subdone;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 5'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b1 == ap_condition_pp0_exit_iter0_state4) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_subdone))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_subdone))) begin
            if ((1'b1 == ap_condition_pp0_exit_iter0_state4)) begin
                ap_enable_reg_pp0_iter1 <= (1'b1 ^ ap_condition_pp0_exit_iter0_state4);
            end else if ((1'b1 == 1'b1)) begin
                ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
            end
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_subdone))) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            ap_enable_reg_pp0_iter2 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln19_reg_1022 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        ii_reg_236 <= select_ln19_19_reg_1084;
    end else if ((1'b1 == ap_CS_fsm_state2)) begin
        ii_reg_236 <= 2'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln19_reg_1022 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        indvar_flatten47_reg_224 <= add_ln19_4_reg_1079;
    end else if ((1'b1 == ap_CS_fsm_state2)) begin
        indvar_flatten47_reg_224 <= 6'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln19_reg_1022 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        indvar_flatten_reg_248 <= select_ln20_20_reg_1123;
    end else if ((1'b1 == ap_CS_fsm_state2)) begin
        indvar_flatten_reg_248 <= 5'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln19_reg_1022 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        jj_reg_259 <= select_ln20_16_reg_1097;
    end else if ((1'b1 == ap_CS_fsm_state2)) begin
        jj_reg_259 <= 2'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln19_reg_1022_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001))) begin
        kk_0_i_i_reg_271 <= add_ln25_reg_1128;
    end else if ((1'b1 == ap_CS_fsm_state2)) begin
        kk_0_i_i_reg_271 <= 5'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
        add_ln19_4_reg_1079 <= add_ln19_4_fu_517_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (icmp_ln19_fu_407_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        add_ln19_reg_1026 <= add_ln19_fu_413_p2;
        add_ln20_4_reg_1074 <= add_ln20_4_fu_511_p2;
        add_ln20_reg_1061 <= add_ln20_fu_470_p2;
        icmp_ln20_reg_1031 <= icmp_ln20_fu_419_p2;
        or_ln23_18_reg_1054 <= or_ln23_18_fu_465_p2;
        or_ln23_20_reg_1067 <= or_ln23_20_fu_505_p2;
        p_cast5_i_i_mid1_reg_1048 <= p_cast5_i_i_mid1_fu_446_p2;
        select_ln19_reg_1043 <= select_ln19_fu_425_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln19_reg_1022 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        add_ln25_reg_1128 <= add_ln25_fu_765_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln19_reg_1022_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001))) begin
        add_ln33_4_reg_1140 <= add_ln33_4_fu_818_p2;
        add_ln33_reg_1133 <= add_ln33_fu_797_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln19_reg_1022 == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001))) begin
        empty_97_reg_1111 <= empty_97_fu_732_p1;
        select_ln20_17_reg_1103 <= select_ln20_17_fu_636_p3;
        select_ln20_reg_1091 <= select_ln20_fu_619_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
        empty_97_reg_1111_pp0_iter1_reg <= empty_97_reg_1111;
        select_ln20_17_reg_1103_pp0_iter1_reg <= select_ln20_17_reg_1103;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state1)) begin
        empty_reg_974 <= empty_fu_287_p1;
        indices_01_read_reg_959 <= indices_01_dout;
        indices_12_read_reg_969 <= indices_12_dout;
        trunc_ln250_reg_964 <= trunc_ln250_fu_282_p1;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        icmp_ln19_reg_1022 <= icmp_ln19_fu_407_p2;
        icmp_ln19_reg_1022_pp0_iter1_reg <= icmp_ln19_reg_1022;
        icmp_ln19_reg_1022_pp0_iter2_reg <= icmp_ln19_reg_1022_pp0_iter1_reg;
        is_padding_reg_1015 <= is_padding_fu_401_p2;
        p_cast5_i_i_reg_1009 <= p_cast5_i_i_fu_361_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        or_ln23_16_reg_999 <= or_ln23_16_fu_337_p2;
        p_cast_i_i_reg_981 <= p_cast_i_i_fu_304_p1;
        p_cast_reg_993 <= p_cast_fu_318_p2;
        p_mid137_reg_1004 <= p_mid137_fu_343_p2;
        sext_ln22_reg_987 <= sext_ln22_fu_314_p1;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln19_reg_1022 == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001))) begin
        select_ln19_19_reg_1084 <= select_ln19_19_fu_555_p3;
        select_ln20_16_reg_1097 <= select_ln20_16_fu_627_p3;
        select_ln20_20_reg_1123 <= select_ln20_20_fu_759_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (icmp_ln19_reg_1022_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        select_ln33_17_reg_1145 <= select_ln33_17_fu_897_p3;
        select_ln33_18_reg_1150 <= select_ln33_18_fu_918_p3;
    end
end

always @ (*) begin
    if ((icmp_ln19_reg_1022 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state4 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state4 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state9)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln19_reg_1022 == 1'd0) & (1'b0 == ap_block_pp0_stage0))) begin
        ap_phi_mux_ii_phi_fu_240_p4 = select_ln19_19_reg_1084;
    end else begin
        ap_phi_mux_ii_phi_fu_240_p4 = ii_reg_236;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln19_reg_1022 == 1'd0) & (1'b0 == ap_block_pp0_stage0))) begin
        ap_phi_mux_indvar_flatten47_phi_fu_228_p4 = add_ln19_4_reg_1079;
    end else begin
        ap_phi_mux_indvar_flatten47_phi_fu_228_p4 = indvar_flatten47_reg_224;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln19_reg_1022 == 1'd0) & (1'b0 == ap_block_pp0_stage0))) begin
        ap_phi_mux_indvar_flatten_phi_fu_252_p4 = select_ln20_20_reg_1123;
    end else begin
        ap_phi_mux_indvar_flatten_phi_fu_252_p4 = indvar_flatten_reg_248;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln19_reg_1022 == 1'd0) & (1'b0 == ap_block_pp0_stage0))) begin
        ap_phi_mux_jj_phi_fu_263_p4 = select_ln20_16_reg_1097;
    end else begin
        ap_phi_mux_jj_phi_fu_263_p4 = jj_reg_259;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln19_reg_1022_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage1))) begin
        ap_phi_mux_kk_0_i_i_phi_fu_275_p4 = add_ln25_reg_1128;
    end else begin
        ap_phi_mux_kk_0_i_i_phi_fu_275_p4 = kk_0_i_i_reg_271;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state9)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((ap_enable_reg_pp0_iter2 == 1'b1)) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ifmap_vec_address0 = sext_ln33_8_fu_954_p1;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0))) begin
            ifmap_vec_address0 = sext_ln33_fu_856_p1;
        end else begin
            ifmap_vec_address0 = 'bx;
        end
    end else begin
        ifmap_vec_address0 = 'bx;
    end
end

always @ (*) begin
    if ((ap_enable_reg_pp0_iter2 == 1'b1)) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ifmap_vec_address1 = sext_ln33_7_fu_937_p1;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0))) begin
            ifmap_vec_address1 = zext_ln33_17_fu_824_p1;
        end else begin
            ifmap_vec_address1 = 'bx;
        end
    end else begin
        ifmap_vec_address1 = 'bx;
    end
end

always @ (*) begin
    if ((((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_11001)) | ((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
        ifmap_vec_ce0 = 1'b1;
    end else begin
        ifmap_vec_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_11001)) | ((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
        ifmap_vec_ce1 = 1'b1;
    end else begin
        ifmap_vec_ce1 = 1'b0;
    end
end

always @ (*) begin
    if ((ap_enable_reg_pp0_iter2 == 1'b1)) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ifmap_vec_d0 = select_ln33_18_reg_1150;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0))) begin
            ifmap_vec_d0 = select_ln33_16_fu_875_p3;
        end else begin
            ifmap_vec_d0 = 'bx;
        end
    end else begin
        ifmap_vec_d0 = 'bx;
    end
end

always @ (*) begin
    if ((ap_enable_reg_pp0_iter2 == 1'b1)) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ifmap_vec_d1 = select_ln33_17_reg_1145;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0))) begin
            ifmap_vec_d1 = select_ln33_fu_836_p3;
        end else begin
            ifmap_vec_d1 = 'bx;
        end
    end else begin
        ifmap_vec_d1 = 'bx;
    end
end

always @ (*) begin
    if ((((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln19_reg_1022_pp0_iter2_reg == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001)) | ((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (icmp_ln19_reg_1022_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
        ifmap_vec_we0 = 1'b1;
    end else begin
        ifmap_vec_we0 = 1'b0;
    end
end

always @ (*) begin
    if ((((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln19_reg_1022_pp0_iter2_reg == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001)) | ((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (icmp_ln19_reg_1022_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
        ifmap_vec_we1 = 1'b1;
    end else begin
        ifmap_vec_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001)) | ((1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b0 == ap_block_pp0_stage1_11001)) | ((1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage1_11001)) | ((1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
        in_data_ce0 = 1'b1;
    end else begin
        in_data_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_01_blk_n = indices_01_empty_n;
    end else begin
        indices_01_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_01_out_blk_n = indices_01_out_full_n;
    end else begin
        indices_01_out_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((indices_12_out_full_n == 1'b0) | (indices_01_out_full_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_01_out_write = 1'b1;
    end else begin
        indices_01_out_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((indices_12_out_full_n == 1'b0) | (indices_01_out_full_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_01_read = 1'b1;
    end else begin
        indices_01_read = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_12_blk_n = indices_12_empty_n;
    end else begin
        indices_12_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_12_out_blk_n = indices_12_out_full_n;
    end else begin
        indices_12_out_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((indices_12_out_full_n == 1'b0) | (indices_01_out_full_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_12_out_write = 1'b1;
    end else begin
        indices_12_out_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((indices_12_out_full_n == 1'b0) | (indices_01_out_full_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_12_read = 1'b1;
    end else begin
        indices_12_read = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((indices_12_out_full_n == 1'b0) | (indices_01_out_full_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_state2 : begin
            ap_NS_fsm = ap_ST_fsm_pp0_stage0;
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_pp0_stage1 : begin
            if ((~((ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln19_reg_1022 == 1'd1) & (1'b0 == ap_block_pp0_stage1_subdone)) & ~((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b0) & (1'b0 == ap_block_pp0_stage1_subdone)) & (1'b0 == ap_block_pp0_stage1_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if ((((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b0) & (1'b0 == ap_block_pp0_stage1_subdone)) | ((ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln19_reg_1022 == 1'd1) & (1'b0 == ap_block_pp0_stage1_subdone)))) begin
                ap_NS_fsm = ap_ST_fsm_state9;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end
        end
        ap_ST_fsm_state9 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln19_4_fu_517_p2 = (indvar_flatten47_reg_224 + 6'd1);

assign add_ln19_fu_413_p2 = (ap_phi_mux_ii_phi_fu_240_p4 + 2'd1);

assign add_ln20_4_fu_511_p2 = (ap_phi_mux_indvar_flatten_phi_fu_252_p4 + 5'd1);

assign add_ln20_fu_470_p2 = (select_ln19_fu_425_p3 + 2'd1);

assign add_ln22_4_fu_376_p2 = ((sext_ln22_reg_987) + (zext_ln20_fu_372_p1));

assign add_ln22_5_fu_480_p2 = ((sext_ln22_reg_987) + (zext_ln20_4_fu_476_p1));

assign add_ln22_fu_308_p2 = ((j_cast_i_i_fu_292_p1) + (17'd131071));

assign add_ln25_fu_765_p2 = (select_ln20_reg_1091 + 5'd4);

assign add_ln32_fu_726_p2 = ((sext_ln20_fu_710_p1) + (zext_ln32_19_fu_722_p1));

assign add_ln33_4_fu_818_p2 = (tmp_80_cast_fu_807_p3 + zext_ln33_16_fu_815_p1);

assign add_ln33_fu_797_p2 = ((sub_ln33_cast_fu_790_p1) + (zext_ln33_15_fu_794_p1));

assign and_ln19_fu_608_p2 = (xor_ln19_fu_597_p2 & icmp_ln25_fu_602_p2);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_pp0_stage1 = ap_CS_fsm[32'd3];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state9 = ap_CS_fsm[32'd4];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((indices_12_out_full_n == 1'b0) | (indices_01_out_full_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0));
end

assign ap_block_state3_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage1_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage1_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage1_iter2 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign bitcast_ln32_16_fu_871_p1 = tmp_44_i_i_fu_861_p4;

assign bitcast_ln32_17_fu_893_p1 = tmp_45_i_i_fu_883_p4;

assign bitcast_ln32_18_fu_914_p1 = tmp_46_i_i_fu_904_p4;

assign bitcast_ln32_fu_832_p1 = trunc_ln32_fu_828_p1;

assign col_coord_int_fu_548_p3 = ((is_padding_reg_1015[0:0] == 1'b1) ? 12'd0 : empty_95_fu_543_p2);

assign col_coord_int_mid139_fu_577_p3 = ((or_ln23_18_reg_1054[0:0] == 1'b1) ? 12'd0 : p_mid137_reg_1004);

assign col_coord_int_mid1_fu_665_p3 = ((or_ln23_20_reg_1067[0:0] == 1'b1) ? 12'd0 : p_mid1_fu_660_p2);

assign empty_92_fu_298_p2 = ((zext_ln19_fu_295_p1) + (17'd131071));

assign empty_93_fu_356_p2 = ((p_cast_i_i_reg_981) + (ii_cast_i_i_fu_348_p1));

assign empty_94_fu_366_p2 = ((empty_93_fu_356_p2 > 18'd55) ? 1'b1 : 1'b0);

assign empty_95_fu_543_p2 = ((tmp1_cast_fu_539_p1) + (empty_reg_974));

assign empty_97_fu_732_p1 = select_ln20_fu_619_p3[3:0];

assign empty_fu_287_p1 = indices_12_dout[11:0];

assign icmp_ln19_fu_407_p2 = ((ap_phi_mux_indvar_flatten47_phi_fu_228_p4 == 6'd36) ? 1'b1 : 1'b0);

assign icmp_ln20_fu_419_p2 = ((ap_phi_mux_indvar_flatten_phi_fu_252_p4 == 5'd12) ? 1'b1 : 1'b0);

assign icmp_ln24_4_fu_389_p2 = (((add_ln22_4_fu_376_p2) > (18'd55)) ? 1'b1 : 1'b0);

assign icmp_ln24_5_fu_493_p2 = (((add_ln22_5_fu_480_p2) > (18'd55)) ? 1'b1 : 1'b0);

assign icmp_ln24_fu_331_p2 = (((add_ln22_fu_308_p2) > (17'd55)) ? 1'b1 : 1'b0);

assign icmp_ln25_fu_602_p2 = ((ap_phi_mux_kk_0_i_i_phi_fu_275_p4 == 5'd16) ? 1'b1 : 1'b0);

assign ii_cast_fu_352_p1 = ap_phi_mux_ii_phi_fu_240_p4;

assign ii_cast_i_i_fu_348_p1 = ap_phi_mux_ii_phi_fu_240_p4;

assign ii_cast_i_i_mid1_fu_433_p1 = add_ln19_fu_413_p2;

assign ii_cast_mid1_fu_437_p1 = add_ln19_fu_413_p2;

assign in_data_address0 = sext_ln32_fu_754_p1;

assign indices_01_out_din = indices_01_dout[5:0];

assign indices_12_out_din = indices_12_dout[11:0];

assign is_padding_fu_401_p2 = (or_ln23_fu_395_p2 | empty_94_fu_366_p2);

assign j_cast_i_i_fu_292_p1 = indices_12_read_reg_969;

assign lshr_ln_fu_736_p4 = {{select_ln20_fu_619_p3[3:2]}};

assign or_ln20_fu_614_p2 = (icmp_ln20_reg_1031 | and_ln19_fu_608_p2);

assign or_ln23_16_fu_337_p2 = (tmp_26_fu_323_p3 | icmp_ln24_fu_331_p2);

assign or_ln23_18_fu_465_p2 = (p_mid113_fu_451_p2 | or_ln23_16_reg_999);

assign or_ln23_19_fu_499_p2 = (tmp_28_fu_485_p3 | icmp_ln24_5_fu_493_p2);

assign or_ln23_20_fu_505_p2 = (select_ln19_21_fu_457_p3 | or_ln23_19_fu_499_p2);

assign or_ln23_fu_395_p2 = (tmp_27_fu_381_p3 | icmp_ln24_4_fu_389_p2);

assign or_ln25_11_fu_925_p2 = (empty_97_reg_1111_pp0_iter1_reg | 4'd2);

assign or_ln25_12_fu_942_p2 = (empty_97_reg_1111_pp0_iter1_reg | 4'd3);

assign or_ln25_fu_844_p2 = (empty_97_reg_1111_pp0_iter1_reg | 4'd1);

assign p_cast5_i_i_fu_361_p2 = (p_cast_reg_993 + ii_cast_fu_352_p1);

assign p_cast5_i_i_mid1_fu_446_p2 = (p_cast_reg_993 + ii_cast_mid1_fu_437_p1);

assign p_cast_fu_318_p2 = ((trunc_ln250_reg_964) + (6'd63));

assign p_cast_i_i_fu_304_p1 = (empty_92_fu_298_p2);

assign p_mid111_fu_441_p2 = ((p_cast_i_i_reg_981) + (ii_cast_i_i_mid1_fu_433_p1));

assign p_mid113_fu_451_p2 = ((p_mid111_fu_441_p2 > 18'd55) ? 1'b1 : 1'b0);

assign p_mid137_fu_343_p2 = ((empty_reg_974) + (12'd4095));

assign p_mid1_fu_660_p2 = ((tmp1_cast_mid1_fu_656_p1) + (empty_reg_974));

assign row_coord_int_fu_527_p3 = ((is_padding_reg_1015[0:0] == 1'b1) ? 6'd0 : p_cast5_i_i_reg_1009);

assign row_coord_int_mid131_fu_571_p3 = ((or_ln23_18_reg_1054[0:0] == 1'b1) ? 6'd0 : p_cast5_i_i_mid1_reg_1048);

assign row_coord_int_mid1_fu_643_p3 = ((or_ln23_20_reg_1067[0:0] == 1'b1) ? 6'd0 : select_ln19_20_fu_561_p3);

assign select_ln19_19_fu_555_p3 = ((icmp_ln20_reg_1031[0:0] == 1'b1) ? add_ln19_reg_1026 : ii_reg_236);

assign select_ln19_20_fu_561_p3 = ((icmp_ln20_reg_1031[0:0] == 1'b1) ? p_cast5_i_i_mid1_reg_1048 : p_cast5_i_i_reg_1009);

assign select_ln19_21_fu_457_p3 = ((icmp_ln20_fu_419_p2[0:0] == 1'b1) ? p_mid113_fu_451_p2 : empty_94_fu_366_p2);

assign select_ln19_22_fu_566_p3 = ((icmp_ln20_reg_1031[0:0] == 1'b1) ? or_ln23_18_reg_1054 : is_padding_reg_1015);

assign select_ln19_23_fu_583_p3 = ((icmp_ln20_reg_1031[0:0] == 1'b1) ? row_coord_int_mid131_fu_571_p3 : row_coord_int_fu_527_p3);

assign select_ln19_24_fu_590_p3 = ((icmp_ln20_reg_1031[0:0] == 1'b1) ? col_coord_int_mid139_fu_577_p3 : col_coord_int_fu_548_p3);

assign select_ln19_fu_425_p3 = ((icmp_ln20_fu_419_p2[0:0] == 1'b1) ? 2'd0 : ap_phi_mux_jj_phi_fu_263_p4);

assign select_ln20_16_fu_627_p3 = ((and_ln19_fu_608_p2[0:0] == 1'b1) ? add_ln20_reg_1061 : select_ln19_reg_1043);

assign select_ln20_17_fu_636_p3 = ((and_ln19_fu_608_p2[0:0] == 1'b1) ? or_ln23_20_reg_1067 : select_ln19_22_fu_566_p3);

assign select_ln20_18_fu_672_p3 = ((and_ln19_fu_608_p2[0:0] == 1'b1) ? row_coord_int_mid1_fu_643_p3 : select_ln19_23_fu_583_p3);

assign select_ln20_19_fu_714_p3 = ((and_ln19_fu_608_p2[0:0] == 1'b1) ? col_coord_int_mid1_fu_665_p3 : select_ln19_24_fu_590_p3);

assign select_ln20_20_fu_759_p3 = ((icmp_ln20_reg_1031[0:0] == 1'b1) ? 5'd1 : add_ln20_4_reg_1074);

assign select_ln20_fu_619_p3 = ((or_ln20_fu_614_p2[0:0] == 1'b1) ? 5'd0 : ap_phi_mux_kk_0_i_i_phi_fu_275_p4);

assign select_ln33_16_fu_875_p3 = ((select_ln20_17_reg_1103_pp0_iter1_reg[0:0] == 1'b1) ? 16'd0 : bitcast_ln32_16_fu_871_p1);

assign select_ln33_17_fu_897_p3 = ((select_ln20_17_reg_1103_pp0_iter1_reg[0:0] == 1'b1) ? 16'd0 : bitcast_ln32_17_fu_893_p1);

assign select_ln33_18_fu_918_p3 = ((select_ln20_17_reg_1103_pp0_iter1_reg[0:0] == 1'b1) ? 16'd0 : bitcast_ln32_18_fu_914_p1);

assign select_ln33_fu_836_p3 = ((select_ln20_17_reg_1103_pp0_iter1_reg[0:0] == 1'b1) ? 16'd0 : bitcast_ln32_fu_832_p1);

assign sext_ln20_fu_710_p1 = (sub_ln32_fu_704_p2);

assign sext_ln22_fu_314_p1 = add_ln22_fu_308_p2;

assign sext_ln32_fu_754_p1 = (tmp_29_fu_746_p3);

assign sext_ln33_7_fu_937_p1 = (tmp_31_fu_930_p3);

assign sext_ln33_8_fu_954_p1 = (tmp_32_fu_947_p3);

assign sext_ln33_fu_856_p1 = (tmp_30_fu_849_p3);

assign sub_ln32_fu_704_p2 = (zext_ln32_fu_688_p1 - zext_ln32_18_fu_700_p1);

assign sub_ln33_cast_fu_790_p1 = (sub_ln33_fu_784_p2);

assign sub_ln33_fu_784_p2 = (zext_ln33_14_fu_780_p1 - zext_ln33_fu_770_p1);

assign tmp1_cast_fu_539_p1 = (tmp1_fu_533_p2);

assign tmp1_cast_mid1_fu_656_p1 = (tmp1_mid1_fu_650_p2);

assign tmp1_fu_533_p2 = ((zext_ln22_fu_523_p1) + (3'd7));

assign tmp1_mid1_fu_650_p2 = ((zext_ln22_4_fu_633_p1) + (3'd7));

assign tmp_26_fu_323_p3 = add_ln22_fu_308_p2[32'd16];

assign tmp_27_fu_381_p3 = add_ln22_4_fu_376_p2[32'd17];

assign tmp_28_fu_485_p3 = add_ln22_5_fu_480_p2[32'd17];

assign tmp_29_fu_746_p3 = {{add_ln32_fu_726_p2}, {lshr_ln_fu_736_p4}};

assign tmp_30_fu_849_p3 = {{add_ln33_reg_1133}, {or_ln25_fu_844_p2}};

assign tmp_31_fu_930_p3 = {{add_ln33_reg_1133}, {or_ln25_11_fu_925_p2}};

assign tmp_32_fu_947_p3 = {{add_ln33_reg_1133}, {or_ln25_12_fu_942_p2}};

assign tmp_44_i_i_fu_861_p4 = {{in_data_q0[31:16]}};

assign tmp_45_i_i_fu_883_p4 = {{in_data_q0[47:32]}};

assign tmp_46_i_i_fu_904_p4 = {{in_data_q0[63:48]}};

assign tmp_6_fu_692_p3 = {{select_ln20_18_fu_672_p3}, {3'd0}};

assign tmp_80_cast_fu_807_p3 = {{trunc_ln33_fu_803_p1}, {4'd0}};

assign tmp_fu_773_p3 = {{select_ln19_19_reg_1084}, {2'd0}};

assign tmp_s_fu_680_p3 = {{select_ln20_18_fu_672_p3}, {6'd0}};

assign trunc_ln250_fu_282_p1 = indices_01_dout[5:0];

assign trunc_ln32_fu_828_p1 = in_data_q0[15:0];

assign trunc_ln33_fu_803_p1 = add_ln33_fu_797_p2[3:0];

assign xor_ln19_fu_597_p2 = (icmp_ln20_reg_1031 ^ 1'd1);

assign zext_ln19_fu_295_p1 = indices_01_read_reg_959;

assign zext_ln20_4_fu_476_p1 = add_ln20_fu_470_p2;

assign zext_ln20_fu_372_p1 = ap_phi_mux_jj_phi_fu_263_p4;

assign zext_ln22_4_fu_633_p1 = add_ln20_reg_1061;

assign zext_ln22_fu_523_p1 = jj_reg_259;

assign zext_ln32_18_fu_700_p1 = tmp_6_fu_692_p3;

assign zext_ln32_19_fu_722_p1 = select_ln20_19_fu_714_p3;

assign zext_ln32_fu_688_p1 = tmp_s_fu_680_p3;

assign zext_ln33_14_fu_780_p1 = tmp_fu_773_p3;

assign zext_ln33_15_fu_794_p1 = select_ln20_16_reg_1097;

assign zext_ln33_16_fu_815_p1 = select_ln20_reg_1091;

assign zext_ln33_17_fu_824_p1 = add_ln33_4_reg_1140;

assign zext_ln33_fu_770_p1 = select_ln19_19_reg_1084;

endmodule //td_fused_top_tdf4_readInputs37
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf5_110 (
        in_data_address0,
        in_data_ce0,
        in_data_d0,
        in_data_q0,
        in_data_we0,
        in_data_address1,
        in_data_ce1,
        in_data_d1,
        in_data_q1,
        in_data_we1,
        out_data_address0,
        out_data_ce0,
        out_data_d0,
        out_data_q0,
        out_data_we0,
        out_data_address1,
        out_data_ce1,
        out_data_d1,
        out_data_q1,
        out_data_we1,
        filter_data_address0,
        filter_data_ce0,
        filter_data_d0,
        filter_data_q0,
        filter_data_we0,
        filter_data_address1,
        filter_data_ce1,
        filter_data_d1,
        filter_data_q1,
        filter_data_we1,
        adjustments_address0,
        adjustments_ce0,
        adjustments_d0,
        adjustments_q0,
        adjustments_we0,
        adjustments_address1,
        adjustments_ce1,
        adjustments_d1,
        adjustments_q1,
        adjustments_we1,
        ap_clk,
        ap_rst,
        in_data_empty_n,
        in_data_read,
        out_data_full_n,
        out_data_write,
        ap_start,
        ap_done,
        ap_ready,
        ap_idle,
        ap_continue
);


output  [13:0] in_data_address0;
output   in_data_ce0;
output  [63:0] in_data_d0;
input  [63:0] in_data_q0;
output   in_data_we0;
output  [13:0] in_data_address1;
output   in_data_ce1;
output  [63:0] in_data_d1;
input  [63:0] in_data_q1;
output   in_data_we1;
output  [14:0] out_data_address0;
output   out_data_ce0;
output  [63:0] out_data_d0;
input  [63:0] out_data_q0;
output   out_data_we0;
output  [14:0] out_data_address1;
output   out_data_ce1;
output  [63:0] out_data_d1;
input  [63:0] out_data_q1;
output   out_data_we1;
output  [14:0] filter_data_address0;
output   filter_data_ce0;
output  [15:0] filter_data_d0;
input  [15:0] filter_data_q0;
output   filter_data_we0;
output  [14:0] filter_data_address1;
output   filter_data_ce1;
output  [15:0] filter_data_d1;
input  [15:0] filter_data_q1;
output   filter_data_we1;
output  [6:0] adjustments_address0;
output   adjustments_ce0;
output  [47:0] adjustments_d0;
input  [47:0] adjustments_q0;
output   adjustments_we0;
output  [6:0] adjustments_address1;
output   adjustments_ce1;
output  [47:0] adjustments_d1;
input  [47:0] adjustments_q1;
output   adjustments_we1;
input   ap_clk;
input   ap_rst;
input   in_data_empty_n;
output   in_data_read;
input   out_data_full_n;
output   out_data_write;
input   ap_start;
output   ap_done;
output   ap_ready;
output   ap_idle;
input   ap_continue;

reg ap_done;
reg ap_ready;
reg ap_idle;

wire   [13:0] dataflow_in_loop_TOP_LOOP37738_U0_in_data_address0;
wire    dataflow_in_loop_TOP_LOOP37738_U0_in_data_ce0;
wire   [63:0] dataflow_in_loop_TOP_LOOP37738_U0_in_data_d0;
wire    dataflow_in_loop_TOP_LOOP37738_U0_in_data_we0;
wire   [13:0] dataflow_in_loop_TOP_LOOP37738_U0_in_data_address1;
wire    dataflow_in_loop_TOP_LOOP37738_U0_in_data_ce1;
wire   [63:0] dataflow_in_loop_TOP_LOOP37738_U0_in_data_d1;
wire    dataflow_in_loop_TOP_LOOP37738_U0_in_data_we1;
wire   [14:0] dataflow_in_loop_TOP_LOOP37738_U0_filter_data_address0;
wire    dataflow_in_loop_TOP_LOOP37738_U0_filter_data_ce0;
wire   [15:0] dataflow_in_loop_TOP_LOOP37738_U0_filter_data_d0;
wire    dataflow_in_loop_TOP_LOOP37738_U0_filter_data_we0;
wire   [14:0] dataflow_in_loop_TOP_LOOP37738_U0_filter_data_address1;
wire    dataflow_in_loop_TOP_LOOP37738_U0_filter_data_ce1;
wire   [15:0] dataflow_in_loop_TOP_LOOP37738_U0_filter_data_d1;
wire    dataflow_in_loop_TOP_LOOP37738_U0_filter_data_we1;
wire   [6:0] dataflow_in_loop_TOP_LOOP37738_U0_adjustments_address0;
wire    dataflow_in_loop_TOP_LOOP37738_U0_adjustments_ce0;
wire   [47:0] dataflow_in_loop_TOP_LOOP37738_U0_adjustments_d0;
wire    dataflow_in_loop_TOP_LOOP37738_U0_adjustments_we0;
wire   [6:0] dataflow_in_loop_TOP_LOOP37738_U0_adjustments_address1;
wire    dataflow_in_loop_TOP_LOOP37738_U0_adjustments_ce1;
wire   [47:0] dataflow_in_loop_TOP_LOOP37738_U0_adjustments_d1;
wire    dataflow_in_loop_TOP_LOOP37738_U0_adjustments_we1;
wire   [14:0] dataflow_in_loop_TOP_LOOP37738_U0_out_data_address0;
wire    dataflow_in_loop_TOP_LOOP37738_U0_out_data_ce0;
wire   [63:0] dataflow_in_loop_TOP_LOOP37738_U0_out_data_d0;
wire    dataflow_in_loop_TOP_LOOP37738_U0_out_data_we0;
wire   [14:0] dataflow_in_loop_TOP_LOOP37738_U0_out_data_address1;
wire    dataflow_in_loop_TOP_LOOP37738_U0_out_data_ce1;
wire   [63:0] dataflow_in_loop_TOP_LOOP37738_U0_out_data_d1;
wire    dataflow_in_loop_TOP_LOOP37738_U0_out_data_we1;
wire    dataflow_in_loop_TOP_LOOP37738_U0_ap_start;
wire    dataflow_in_loop_TOP_LOOP37738_U0_in_data_read;
wire    dataflow_in_loop_TOP_LOOP37738_U0_out_data_write;
wire    dataflow_in_loop_TOP_LOOP37738_U0_ap_done;
wire    dataflow_in_loop_TOP_LOOP37738_U0_ap_ready;
wire    dataflow_in_loop_TOP_LOOP37738_U0_ap_idle;
reg    dataflow_in_loop_TOP_LOOP37738_U0_ap_continue;
wire    dataflow_in_loop_TOP_LOOP37738_U0_in_data_full_n;
wire    dataflow_in_loop_TOP_LOOP37738_U0_in_data_write;
wire    ap_sync_continue;
wire    ap_sync_done;
wire    ap_sync_ready;
reg   [18:0] loop_dataflow_input_count;
reg   [18:0] loop_dataflow_output_count;
wire   [18:0] bound_minus_1;
wire    dataflow_in_loop_TOP_LOOP37738_U0_start_full_n;
wire    dataflow_in_loop_TOP_LOOP37738_U0_start_write;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 loop_dataflow_input_count = 19'd0;
#0 loop_dataflow_output_count = 19'd0;
end

td_fused_top_dataflow_in_loop_TOP_LOOP37738 dataflow_in_loop_TOP_LOOP37738_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .in_data_address0(dataflow_in_loop_TOP_LOOP37738_U0_in_data_address0),
    .in_data_ce0(dataflow_in_loop_TOP_LOOP37738_U0_in_data_ce0),
    .in_data_d0(dataflow_in_loop_TOP_LOOP37738_U0_in_data_d0),
    .in_data_q0(in_data_q0),
    .in_data_we0(dataflow_in_loop_TOP_LOOP37738_U0_in_data_we0),
    .in_data_address1(dataflow_in_loop_TOP_LOOP37738_U0_in_data_address1),
    .in_data_ce1(dataflow_in_loop_TOP_LOOP37738_U0_in_data_ce1),
    .in_data_d1(dataflow_in_loop_TOP_LOOP37738_U0_in_data_d1),
    .in_data_q1(64'd0),
    .in_data_we1(dataflow_in_loop_TOP_LOOP37738_U0_in_data_we1),
    .filter_data_address0(dataflow_in_loop_TOP_LOOP37738_U0_filter_data_address0),
    .filter_data_ce0(dataflow_in_loop_TOP_LOOP37738_U0_filter_data_ce0),
    .filter_data_d0(dataflow_in_loop_TOP_LOOP37738_U0_filter_data_d0),
    .filter_data_q0(filter_data_q0),
    .filter_data_we0(dataflow_in_loop_TOP_LOOP37738_U0_filter_data_we0),
    .filter_data_address1(dataflow_in_loop_TOP_LOOP37738_U0_filter_data_address1),
    .filter_data_ce1(dataflow_in_loop_TOP_LOOP37738_U0_filter_data_ce1),
    .filter_data_d1(dataflow_in_loop_TOP_LOOP37738_U0_filter_data_d1),
    .filter_data_q1(16'd0),
    .filter_data_we1(dataflow_in_loop_TOP_LOOP37738_U0_filter_data_we1),
    .adjustments_address0(dataflow_in_loop_TOP_LOOP37738_U0_adjustments_address0),
    .adjustments_ce0(dataflow_in_loop_TOP_LOOP37738_U0_adjustments_ce0),
    .adjustments_d0(dataflow_in_loop_TOP_LOOP37738_U0_adjustments_d0),
    .adjustments_q0(adjustments_q0),
    .adjustments_we0(dataflow_in_loop_TOP_LOOP37738_U0_adjustments_we0),
    .adjustments_address1(dataflow_in_loop_TOP_LOOP37738_U0_adjustments_address1),
    .adjustments_ce1(dataflow_in_loop_TOP_LOOP37738_U0_adjustments_ce1),
    .adjustments_d1(dataflow_in_loop_TOP_LOOP37738_U0_adjustments_d1),
    .adjustments_q1(48'd0),
    .adjustments_we1(dataflow_in_loop_TOP_LOOP37738_U0_adjustments_we1),
    .out_data_address0(dataflow_in_loop_TOP_LOOP37738_U0_out_data_address0),
    .out_data_ce0(dataflow_in_loop_TOP_LOOP37738_U0_out_data_ce0),
    .out_data_d0(dataflow_in_loop_TOP_LOOP37738_U0_out_data_d0),
    .out_data_q0(64'd0),
    .out_data_we0(dataflow_in_loop_TOP_LOOP37738_U0_out_data_we0),
    .out_data_address1(dataflow_in_loop_TOP_LOOP37738_U0_out_data_address1),
    .out_data_ce1(dataflow_in_loop_TOP_LOOP37738_U0_out_data_ce1),
    .out_data_d1(dataflow_in_loop_TOP_LOOP37738_U0_out_data_d1),
    .out_data_q1(64'd0),
    .out_data_we1(dataflow_in_loop_TOP_LOOP37738_U0_out_data_we1),
    .ap_start(dataflow_in_loop_TOP_LOOP37738_U0_ap_start),
    .in_data_empty_n(1'b0),
    .in_data_read(dataflow_in_loop_TOP_LOOP37738_U0_in_data_read),
    .out_data_full_n(out_data_full_n),
    .out_data_write(dataflow_in_loop_TOP_LOOP37738_U0_out_data_write),
    .ap_done(dataflow_in_loop_TOP_LOOP37738_U0_ap_done),
    .ap_ready(dataflow_in_loop_TOP_LOOP37738_U0_ap_ready),
    .ap_idle(dataflow_in_loop_TOP_LOOP37738_U0_ap_idle),
    .ap_continue(dataflow_in_loop_TOP_LOOP37738_U0_ap_continue)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        loop_dataflow_input_count <= 19'd0;
    end else begin
        if ((~(loop_dataflow_input_count == bound_minus_1) & (dataflow_in_loop_TOP_LOOP37738_U0_ap_ready == 1'b1) & (ap_start == 1'b1))) begin
            loop_dataflow_input_count <= (loop_dataflow_input_count + 19'd1);
        end else if (((dataflow_in_loop_TOP_LOOP37738_U0_ap_ready == 1'b1) & (loop_dataflow_input_count == bound_minus_1) & (ap_start == 1'b1))) begin
            loop_dataflow_input_count <= 19'd0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        loop_dataflow_output_count <= 19'd0;
    end else begin
        if ((~(loop_dataflow_output_count == bound_minus_1) & (dataflow_in_loop_TOP_LOOP37738_U0_ap_continue == 1'b1) & (dataflow_in_loop_TOP_LOOP37738_U0_ap_done == 1'b1))) begin
            loop_dataflow_output_count <= (loop_dataflow_output_count + 19'd1);
        end else if (((dataflow_in_loop_TOP_LOOP37738_U0_ap_continue == 1'b1) & (dataflow_in_loop_TOP_LOOP37738_U0_ap_done == 1'b1) & (loop_dataflow_output_count == bound_minus_1))) begin
            loop_dataflow_output_count <= 19'd0;
        end
    end
end

always @ (*) begin
    if (((dataflow_in_loop_TOP_LOOP37738_U0_ap_done == 1'b1) & (loop_dataflow_output_count == bound_minus_1))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = 1'b0;
    end
end

always @ (*) begin
    if (((dataflow_in_loop_TOP_LOOP37738_U0_ap_idle == 1'b1) & (loop_dataflow_output_count == 19'd0) & (ap_start == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((dataflow_in_loop_TOP_LOOP37738_U0_ap_ready == 1'b1) & (loop_dataflow_input_count == bound_minus_1) & (ap_start == 1'b1))) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((~(loop_dataflow_output_count == bound_minus_1) | (ap_continue == 1'b1))) begin
        dataflow_in_loop_TOP_LOOP37738_U0_ap_continue = 1'b1;
    end else begin
        dataflow_in_loop_TOP_LOOP37738_U0_ap_continue = 1'b0;
    end
end

assign adjustments_address0 = dataflow_in_loop_TOP_LOOP37738_U0_adjustments_address0;

assign adjustments_address1 = 7'd0;

assign adjustments_ce0 = dataflow_in_loop_TOP_LOOP37738_U0_adjustments_ce0;

assign adjustments_ce1 = 1'b0;

assign adjustments_d0 = 48'd0;

assign adjustments_d1 = 48'd0;

assign adjustments_we0 = 1'b0;

assign adjustments_we1 = 1'b0;

assign ap_sync_continue = ap_continue;

assign ap_sync_done = dataflow_in_loop_TOP_LOOP37738_U0_ap_done;

assign ap_sync_ready = dataflow_in_loop_TOP_LOOP37738_U0_ap_ready;

assign bound_minus_1 = (19'd401408 - 19'd1);

assign dataflow_in_loop_TOP_LOOP37738_U0_ap_start = ap_start;

assign dataflow_in_loop_TOP_LOOP37738_U0_in_data_full_n = in_data_empty_n;

assign dataflow_in_loop_TOP_LOOP37738_U0_in_data_write = 1'b0;

assign dataflow_in_loop_TOP_LOOP37738_U0_start_full_n = 1'b1;

assign dataflow_in_loop_TOP_LOOP37738_U0_start_write = 1'b0;

assign filter_data_address0 = dataflow_in_loop_TOP_LOOP37738_U0_filter_data_address0;

assign filter_data_address1 = 15'd0;

assign filter_data_ce0 = dataflow_in_loop_TOP_LOOP37738_U0_filter_data_ce0;

assign filter_data_ce1 = 1'b0;

assign filter_data_d0 = 16'd0;

assign filter_data_d1 = 16'd0;

assign filter_data_we0 = 1'b0;

assign filter_data_we1 = 1'b0;

assign in_data_address0 = dataflow_in_loop_TOP_LOOP37738_U0_in_data_address0;

assign in_data_address1 = 14'd0;

assign in_data_ce0 = dataflow_in_loop_TOP_LOOP37738_U0_in_data_ce0;

assign in_data_ce1 = 1'b0;

assign in_data_d0 = 64'd0;

assign in_data_d1 = 64'd0;

assign in_data_read = dataflow_in_loop_TOP_LOOP37738_U0_in_data_write;

assign in_data_we0 = 1'b0;

assign in_data_we1 = 1'b0;

assign out_data_address0 = 15'd0;

assign out_data_address1 = dataflow_in_loop_TOP_LOOP37738_U0_out_data_address1;

assign out_data_ce0 = 1'b0;

assign out_data_ce1 = dataflow_in_loop_TOP_LOOP37738_U0_out_data_ce1;

assign out_data_d0 = 64'd0;

assign out_data_d1 = dataflow_in_loop_TOP_LOOP37738_U0_out_data_d1;

assign out_data_we0 = 1'b0;

assign out_data_we1 = dataflow_in_loop_TOP_LOOP37738_U0_out_data_we1;

assign out_data_write = dataflow_in_loop_TOP_LOOP37738_U0_out_data_write;

endmodule //td_fused_top_tdf5_110
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf5_accum_1 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        accum_in_0_address0,
        accum_in_0_ce0,
        accum_in_0_q0,
        accum_in_0_address1,
        accum_in_0_ce1,
        accum_in_0_q1,
        accum_out_address0,
        accum_out_ce0,
        accum_out_we0,
        accum_out_d0,
        accum_out_address1,
        accum_out_ce1,
        accum_out_we1,
        accum_out_d1
);

parameter    ap_ST_fsm_state1 = 8'd1;
parameter    ap_ST_fsm_pp0_stage0 = 8'd2;
parameter    ap_ST_fsm_pp0_stage1 = 8'd4;
parameter    ap_ST_fsm_pp0_stage2 = 8'd8;
parameter    ap_ST_fsm_pp0_stage3 = 8'd16;
parameter    ap_ST_fsm_state12 = 8'd32;
parameter    ap_ST_fsm_state13 = 8'd64;
parameter    ap_ST_fsm_state14 = 8'd128;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [7:0] accum_in_0_address0;
output   accum_in_0_ce0;
input  [15:0] accum_in_0_q0;
output  [7:0] accum_in_0_address1;
output   accum_in_0_ce1;
input  [15:0] accum_in_0_q1;
output  [2:0] accum_out_address0;
output   accum_out_ce0;
output   accum_out_we0;
output  [15:0] accum_out_d0;
output  [2:0] accum_out_address1;
output   accum_out_ce1;
output   accum_out_we1;
output  [15:0] accum_out_d1;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg[7:0] accum_in_0_address0;
reg accum_in_0_ce0;
reg[7:0] accum_in_0_address1;
reg accum_in_0_ce1;
reg accum_out_ce0;
reg accum_out_we0;
reg accum_out_ce1;
reg accum_out_we1;

reg    ap_done_reg;
  reg   [7:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg   [7:0] x_reg_168;
reg   [15:0] psum_7_08_reg_180;
reg   [15:0] psum_6_07_reg_192;
reg   [15:0] psum_5_06_reg_204;
reg   [15:0] psum_4_05_reg_216;
reg   [15:0] psum_3_04_reg_228;
reg   [15:0] psum_2_03_reg_240;
reg   [15:0] psum_1_02_reg_252;
reg   [15:0] psum_0_01_reg_264;
wire   [0:0] icmp_ln49_fu_321_p2;
reg   [0:0] icmp_ln49_reg_492;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state6_pp0_stage0_iter1;
wire    ap_block_state10_pp0_stage0_iter2;
wire    ap_block_pp0_stage0_11001;
reg   [0:0] icmp_ln49_reg_492_pp0_iter1_reg;
reg   [0:0] icmp_ln49_reg_492_pp0_iter2_reg;
reg   [15:0] accum_in_0_load_reg_506;
wire    ap_CS_fsm_pp0_stage1;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_state3_pp0_stage1_iter0;
wire    ap_block_state7_pp0_stage1_iter1;
wire    ap_block_state11_pp0_stage1_iter2;
wire    ap_block_pp0_stage1_11001;
reg   [15:0] accum_in_0_load_29_reg_511;
reg   [15:0] accum_in_0_load_30_reg_526;
wire    ap_CS_fsm_pp0_stage2;
wire    ap_block_state4_pp0_stage2_iter0;
wire    ap_block_state8_pp0_stage2_iter1;
wire    ap_block_pp0_stage2_11001;
reg   [15:0] accum_in_0_load_31_reg_531;
wire   [7:0] add_ln49_fu_387_p2;
reg   [7:0] add_ln49_reg_546;
wire    ap_CS_fsm_pp0_stage3;
wire    ap_block_state5_pp0_stage3_iter0;
wire    ap_block_state9_pp0_stage3_iter1;
wire    ap_block_pp0_stage3_11001;
reg   [15:0] accum_in_0_load_32_reg_551;
reg   [15:0] accum_in_0_load_33_reg_556;
reg   [15:0] accum_in_0_load_34_reg_571;
reg    ap_enable_reg_pp0_iter1;
reg   [15:0] accum_in_0_load_35_reg_576;
wire   [15:0] grp_fu_305_p2;
wire   [15:0] grp_fu_310_p2;
reg    ap_enable_reg_pp0_iter2;
wire   [3:0] add_ln57_fu_432_p2;
wire    ap_CS_fsm_state13;
wire   [0:0] tmp_fu_415_p3;
reg    ap_block_state1;
wire    ap_block_pp0_stage2_subdone;
reg    ap_condition_pp0_exit_iter0_state4;
wire    ap_block_pp0_stage3_subdone;
wire    ap_block_pp0_stage1_subdone;
reg   [7:0] ap_phi_mux_x_phi_fu_172_p4;
wire    ap_block_pp0_stage0;
wire   [15:0] ap_phi_mux_psum_7_08_phi_fu_184_p4;
wire    ap_block_pp0_stage1;
wire   [15:0] ap_phi_mux_psum_6_07_phi_fu_196_p4;
wire   [15:0] ap_phi_mux_psum_5_06_phi_fu_208_p4;
wire   [15:0] ap_phi_mux_psum_4_05_phi_fu_220_p4;
wire   [15:0] ap_phi_mux_psum_3_04_phi_fu_232_p4;
wire    ap_block_pp0_stage3;
wire   [15:0] ap_phi_mux_psum_2_03_phi_fu_244_p4;
wire    ap_block_pp0_stage2;
reg   [3:0] q_reg_276;
wire    ap_CS_fsm_state12;
reg   [15:0] ap_phi_mux_phi_ln69_phi_fu_290_p8;
wire   [2:0] trunc_ln57_fu_428_p1;
wire   [63:0] zext_ln49_fu_327_p1;
wire   [63:0] zext_ln53_fu_338_p1;
wire   [63:0] zext_ln53_7_fu_349_p1;
wire   [63:0] zext_ln53_8_fu_360_p1;
wire   [63:0] zext_ln53_9_fu_371_p1;
wire   [63:0] zext_ln53_10_fu_382_p1;
wire   [63:0] zext_ln53_11_fu_399_p1;
wire   [63:0] zext_ln53_12_fu_410_p1;
wire   [63:0] zext_ln57_fu_423_p1;
wire   [63:0] zext_ln57_2_fu_444_p1;
reg   [15:0] grp_fu_305_p0;
reg   [15:0] grp_fu_305_p1;
reg   [15:0] grp_fu_310_p0;
reg   [15:0] grp_fu_310_p1;
wire   [7:0] or_ln53_fu_332_p2;
wire   [7:0] or_ln53_7_fu_343_p2;
wire   [7:0] or_ln53_8_fu_354_p2;
wire   [7:0] or_ln53_9_fu_365_p2;
wire   [7:0] or_ln53_10_fu_376_p2;
wire   [7:0] or_ln53_11_fu_393_p2;
wire   [7:0] or_ln53_12_fu_404_p2;
wire   [2:0] or_ln57_fu_438_p2;
wire   [0:0] icmp_ln69_fu_449_p2;
wire   [0:0] icmp_ln69_3_fu_463_p2;
wire   [15:0] select_ln69_fu_455_p3;
wire   [0:0] icmp_ln69_4_fu_477_p2;
wire   [15:0] select_ln69_3_fu_469_p3;
wire    ap_CS_fsm_state14;
reg   [7:0] ap_NS_fsm;
wire    ap_block_pp0_stage0_subdone;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
reg    ap_condition_514;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 8'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
end

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U297(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(grp_fu_305_p0),
    .din1(grp_fu_305_p1),
    .dout(grp_fu_305_p2)
);

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U298(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(grp_fu_310_p0),
    .din1(grp_fu_310_p1),
    .dout(grp_fu_310_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state14)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage2_subdone) & (1'b1 == ap_condition_pp0_exit_iter0_state4) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage3_subdone) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b0)) | ((1'b0 == ap_block_pp0_stage3_subdone) & (1'b1 == ap_CS_fsm_pp0_stage3)))) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end else if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter2 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state12)) begin
        q_reg_276 <= 4'd0;
    end else if (((tmp_fu_415_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state13))) begin
        q_reg_276 <= add_ln57_fu_432_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln49_reg_492 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        x_reg_168 <= add_ln49_reg_546;
    end else if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        x_reg_168 <= 8'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage1_11001) & (icmp_ln49_reg_492 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
        accum_in_0_load_29_reg_511 <= accum_in_0_q0;
        accum_in_0_load_reg_506 <= accum_in_0_q1;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2_11001) & (icmp_ln49_reg_492 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
        accum_in_0_load_30_reg_526 <= accum_in_0_q1;
        accum_in_0_load_31_reg_531 <= accum_in_0_q0;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage3_11001) & (icmp_ln49_reg_492 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
        accum_in_0_load_32_reg_551 <= accum_in_0_q1;
        accum_in_0_load_33_reg_556 <= accum_in_0_q0;
        add_ln49_reg_546 <= add_ln49_fu_387_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln49_reg_492 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        accum_in_0_load_34_reg_571 <= accum_in_0_q1;
        accum_in_0_load_35_reg_576 <= accum_in_0_q0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln49_reg_492 <= icmp_ln49_fu_321_p2;
        icmp_ln49_reg_492_pp0_iter1_reg <= icmp_ln49_reg_492;
        icmp_ln49_reg_492_pp0_iter2_reg <= icmp_ln49_reg_492_pp0_iter1_reg;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln49_reg_492_pp0_iter1_reg == 1'd1) & (1'b0 == ap_block_pp0_stage2_11001) & (1'b1 == ap_CS_fsm_pp0_stage2) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        psum_0_01_reg_264 <= grp_fu_305_p2;
        psum_1_02_reg_252 <= grp_fu_310_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln49_reg_492_pp0_iter1_reg == 1'd1) & (1'b0 == ap_block_pp0_stage3_11001) & (1'b1 == ap_CS_fsm_pp0_stage3) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        psum_2_03_reg_240 <= grp_fu_305_p2;
        psum_3_04_reg_228 <= grp_fu_310_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln49_reg_492_pp0_iter1_reg == 1'd1) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        psum_4_05_reg_216 <= grp_fu_305_p2;
        psum_5_06_reg_204 <= grp_fu_310_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln49_reg_492_pp0_iter2_reg == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        psum_6_07_reg_192 <= grp_fu_305_p2;
        psum_7_08_reg_180 <= grp_fu_310_p2;
    end
end

always @ (*) begin
    if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
        if (((1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            accum_in_0_address0 = zext_ln53_12_fu_410_p1;
        end else if (((1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            accum_in_0_address0 = zext_ln53_10_fu_382_p1;
        end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            accum_in_0_address0 = zext_ln53_8_fu_360_p1;
        end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            accum_in_0_address0 = zext_ln53_fu_338_p1;
        end else begin
            accum_in_0_address0 = 'bx;
        end
    end else begin
        accum_in_0_address0 = 'bx;
    end
end

always @ (*) begin
    if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
        if (((1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            accum_in_0_address1 = zext_ln53_11_fu_399_p1;
        end else if (((1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            accum_in_0_address1 = zext_ln53_9_fu_371_p1;
        end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            accum_in_0_address1 = zext_ln53_7_fu_349_p1;
        end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            accum_in_0_address1 = zext_ln49_fu_327_p1;
        end else begin
            accum_in_0_address1 = 'bx;
        end
    end else begin
        accum_in_0_address1 = 'bx;
    end
end

always @ (*) begin
    if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage3_11001) & (1'b1 == ap_CS_fsm_pp0_stage3)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2_11001) & (1'b1 == ap_CS_fsm_pp0_stage2)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1)))) begin
        accum_in_0_ce0 = 1'b1;
    end else begin
        accum_in_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage3_11001) & (1'b1 == ap_CS_fsm_pp0_stage3)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2_11001) & (1'b1 == ap_CS_fsm_pp0_stage2)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1)))) begin
        accum_in_0_ce1 = 1'b1;
    end else begin
        accum_in_0_ce1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state13)) begin
        accum_out_ce0 = 1'b1;
    end else begin
        accum_out_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state13)) begin
        accum_out_ce1 = 1'b1;
    end else begin
        accum_out_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((tmp_fu_415_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state13))) begin
        accum_out_we0 = 1'b1;
    end else begin
        accum_out_we0 = 1'b0;
    end
end

always @ (*) begin
    if (((tmp_fu_415_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state13))) begin
        accum_out_we1 = 1'b1;
    end else begin
        accum_out_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((icmp_ln49_reg_492 == 1'd0)) begin
        ap_condition_pp0_exit_iter0_state4 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state4 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state14)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((tmp_fu_415_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state13))) begin
        if ((trunc_ln57_fu_428_p1 == 3'd0)) begin
            ap_phi_mux_phi_ln69_phi_fu_290_p8 = psum_0_01_reg_264;
        end else if ((1'b1 == ap_condition_514)) begin
            ap_phi_mux_phi_ln69_phi_fu_290_p8 = psum_6_07_reg_192;
        end else if ((trunc_ln57_fu_428_p1 == 3'd4)) begin
            ap_phi_mux_phi_ln69_phi_fu_290_p8 = psum_4_05_reg_216;
        end else if ((trunc_ln57_fu_428_p1 == 3'd2)) begin
            ap_phi_mux_phi_ln69_phi_fu_290_p8 = psum_2_03_reg_240;
        end else begin
            ap_phi_mux_phi_ln69_phi_fu_290_p8 = 'bx;
        end
    end else begin
        ap_phi_mux_phi_ln69_phi_fu_290_p8 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0) & (icmp_ln49_reg_492 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_x_phi_fu_172_p4 = add_ln49_reg_546;
    end else begin
        ap_phi_mux_x_phi_fu_172_p4 = x_reg_168;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state14)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_305_p0 = ap_phi_mux_psum_6_07_phi_fu_196_p4;
    end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_305_p0 = ap_phi_mux_psum_4_05_phi_fu_220_p4;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
        grp_fu_305_p0 = ap_phi_mux_psum_2_03_phi_fu_244_p4;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
        grp_fu_305_p0 = grp_fu_305_p2;
    end else begin
        grp_fu_305_p0 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_305_p1 = accum_in_0_load_34_reg_571;
    end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_305_p1 = accum_in_0_load_32_reg_551;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
        grp_fu_305_p1 = accum_in_0_load_30_reg_526;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
        grp_fu_305_p1 = accum_in_0_load_reg_506;
    end else begin
        grp_fu_305_p1 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_310_p0 = ap_phi_mux_psum_7_08_phi_fu_184_p4;
    end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_310_p0 = ap_phi_mux_psum_5_06_phi_fu_208_p4;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
        grp_fu_310_p0 = ap_phi_mux_psum_3_04_phi_fu_232_p4;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
        grp_fu_310_p0 = grp_fu_310_p2;
    end else begin
        grp_fu_310_p0 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_310_p1 = accum_in_0_load_35_reg_576;
    end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_310_p1 = accum_in_0_load_33_reg_556;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
        grp_fu_310_p1 = accum_in_0_load_31_reg_531;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
        grp_fu_310_p1 = accum_in_0_load_29_reg_511;
    end else begin
        grp_fu_310_p1 = 'bx;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_pp0_stage1 : begin
            if ((~((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter2 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0)) & (1'b0 == ap_block_pp0_stage1_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage2;
            end else if (((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter2 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
                ap_NS_fsm = ap_ST_fsm_state12;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end
        end
        ap_ST_fsm_pp0_stage2 : begin
            if ((~((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2_subdone) & (icmp_ln49_reg_492 == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b0)) & (1'b0 == ap_block_pp0_stage2_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage3;
            end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2_subdone) & (icmp_ln49_reg_492 == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
                ap_NS_fsm = ap_ST_fsm_state12;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage2;
            end
        end
        ap_ST_fsm_pp0_stage3 : begin
            if ((1'b0 == ap_block_pp0_stage3_subdone)) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage3;
            end
        end
        ap_ST_fsm_state12 : begin
            ap_NS_fsm = ap_ST_fsm_state13;
        end
        ap_ST_fsm_state13 : begin
            if (((tmp_fu_415_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state13))) begin
                ap_NS_fsm = ap_ST_fsm_state13;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state14;
            end
        end
        ap_ST_fsm_state14 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign accum_out_address0 = zext_ln57_2_fu_444_p1;

assign accum_out_address1 = zext_ln57_fu_423_p1;

assign accum_out_d0 = ((icmp_ln69_4_fu_477_p2[0:0] == 1'b1) ? psum_5_06_reg_204 : select_ln69_3_fu_469_p3);

assign accum_out_d1 = ap_phi_mux_phi_ln69_phi_fu_290_p8;

assign add_ln49_fu_387_p2 = (x_reg_168 + 8'd8);

assign add_ln57_fu_432_p2 = (q_reg_276 + 4'd2);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_pp0_stage1 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_pp0_stage2 = ap_CS_fsm[32'd3];

assign ap_CS_fsm_pp0_stage3 = ap_CS_fsm[32'd4];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state12 = ap_CS_fsm[32'd5];

assign ap_CS_fsm_state13 = ap_CS_fsm[32'd6];

assign ap_CS_fsm_state14 = ap_CS_fsm[32'd7];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1_subdone = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage2 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage2_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage2_subdone = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage3 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage3_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage3_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((ap_done_reg == 1'b1) | (ap_start == 1'b0));
end

assign ap_block_state10_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state11_pp0_stage1_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage1_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage2_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage3_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage1_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage2_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state9_pp0_stage3_iter1 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_condition_514 = (~(trunc_ln57_fu_428_p1 == 3'd0) & ~(trunc_ln57_fu_428_p1 == 3'd4) & ~(trunc_ln57_fu_428_p1 == 3'd2));
end

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign ap_phi_mux_psum_2_03_phi_fu_244_p4 = grp_fu_305_p2;

assign ap_phi_mux_psum_3_04_phi_fu_232_p4 = grp_fu_310_p2;

assign ap_phi_mux_psum_4_05_phi_fu_220_p4 = grp_fu_305_p2;

assign ap_phi_mux_psum_5_06_phi_fu_208_p4 = grp_fu_310_p2;

assign ap_phi_mux_psum_6_07_phi_fu_196_p4 = grp_fu_305_p2;

assign ap_phi_mux_psum_7_08_phi_fu_184_p4 = grp_fu_310_p2;

assign icmp_ln49_fu_321_p2 = ((ap_phi_mux_x_phi_fu_172_p4 < 8'd144) ? 1'b1 : 1'b0);

assign icmp_ln69_3_fu_463_p2 = ((or_ln57_fu_438_p2 == 3'd3) ? 1'b1 : 1'b0);

assign icmp_ln69_4_fu_477_p2 = ((or_ln57_fu_438_p2 == 3'd5) ? 1'b1 : 1'b0);

assign icmp_ln69_fu_449_p2 = ((or_ln57_fu_438_p2 == 3'd1) ? 1'b1 : 1'b0);

assign or_ln53_10_fu_376_p2 = (x_reg_168 | 8'd5);

assign or_ln53_11_fu_393_p2 = (x_reg_168 | 8'd6);

assign or_ln53_12_fu_404_p2 = (x_reg_168 | 8'd7);

assign or_ln53_7_fu_343_p2 = (x_reg_168 | 8'd2);

assign or_ln53_8_fu_354_p2 = (x_reg_168 | 8'd3);

assign or_ln53_9_fu_365_p2 = (x_reg_168 | 8'd4);

assign or_ln53_fu_332_p2 = (ap_phi_mux_x_phi_fu_172_p4 | 8'd1);

assign or_ln57_fu_438_p2 = (trunc_ln57_fu_428_p1 | 3'd1);

assign select_ln69_3_fu_469_p3 = ((icmp_ln69_3_fu_463_p2[0:0] == 1'b1) ? psum_3_04_reg_228 : select_ln69_fu_455_p3);

assign select_ln69_fu_455_p3 = ((icmp_ln69_fu_449_p2[0:0] == 1'b1) ? psum_1_02_reg_252 : psum_7_08_reg_180);

assign tmp_fu_415_p3 = q_reg_276[32'd3];

assign trunc_ln57_fu_428_p1 = q_reg_276[2:0];

assign zext_ln49_fu_327_p1 = ap_phi_mux_x_phi_fu_172_p4;

assign zext_ln53_10_fu_382_p1 = or_ln53_10_fu_376_p2;

assign zext_ln53_11_fu_399_p1 = or_ln53_11_fu_393_p2;

assign zext_ln53_12_fu_410_p1 = or_ln53_12_fu_404_p2;

assign zext_ln53_7_fu_349_p1 = or_ln53_7_fu_343_p2;

assign zext_ln53_8_fu_360_p1 = or_ln53_8_fu_354_p2;

assign zext_ln53_9_fu_371_p1 = or_ln53_9_fu_365_p2;

assign zext_ln53_fu_338_p1 = or_ln53_fu_332_p2;

assign zext_ln57_2_fu_444_p1 = or_ln57_fu_438_p2;

assign zext_ln57_fu_423_p1 = q_reg_276;

endmodule //td_fused_top_tdf5_accum_1
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf5_accum_2 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        accum_in_10,
        accum_in_10_ap_vld,
        accum_in_address0,
        accum_in_ce0,
        accum_in_q0
);

parameter    ap_ST_fsm_state1 = 7'd1;
parameter    ap_ST_fsm_state2 = 7'd2;
parameter    ap_ST_fsm_state3 = 7'd4;
parameter    ap_ST_fsm_state4 = 7'd8;
parameter    ap_ST_fsm_state5 = 7'd16;
parameter    ap_ST_fsm_state6 = 7'd32;
parameter    ap_ST_fsm_state7 = 7'd64;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [15:0] accum_in_10;
output   accum_in_10_ap_vld;
output  [2:0] accum_in_address0;
output   accum_in_ce0;
input  [15:0] accum_in_q0;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg[15:0] accum_in_10;
reg accum_in_10_ap_vld;
reg accum_in_ce0;

reg    ap_done_reg;
  reg   [6:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
wire   [3:0] add_ln81_fu_74_p2;
reg   [3:0] add_ln81_reg_91;
wire    ap_CS_fsm_state2;
wire   [0:0] icmp_ln81_fu_85_p2;
wire    ap_CS_fsm_state3;
wire   [15:0] grp_fu_68_p2;
wire    ap_CS_fsm_state7;
reg   [3:0] i_1_1_reg_44;
reg    ap_block_state1;
reg   [15:0] sum_01_reg_55;
wire   [63:0] zext_ln81_fu_80_p1;
reg   [15:0] accum_in_10_preg;
reg   [6:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 7'd1;
#0 accum_in_10_preg = 16'd0;
end

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U301(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(sum_01_reg_55),
    .din1(accum_in_q0),
    .dout(grp_fu_68_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        accum_in_10_preg <= 16'd0;
    end else begin
        if (((icmp_ln81_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
            accum_in_10_preg <= sum_01_reg_55;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if (((icmp_ln81_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        i_1_1_reg_44 <= 4'd0;
    end else if ((1'b1 == ap_CS_fsm_state7)) begin
        i_1_1_reg_44 <= add_ln81_reg_91;
    end
end

always @ (posedge ap_clk) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        sum_01_reg_55 <= 16'd0;
    end else if ((1'b1 == ap_CS_fsm_state7)) begin
        sum_01_reg_55 <= grp_fu_68_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        add_ln81_reg_91 <= add_ln81_fu_74_p2;
    end
end

always @ (*) begin
    if (((icmp_ln81_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        accum_in_10 = sum_01_reg_55;
    end else begin
        accum_in_10 = accum_in_10_preg;
    end
end

always @ (*) begin
    if (((icmp_ln81_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        accum_in_10_ap_vld = 1'b1;
    end else begin
        accum_in_10_ap_vld = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        accum_in_ce0 = 1'b1;
    end else begin
        accum_in_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln81_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln81_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_state2 : begin
            if (((icmp_ln81_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end
        end
        ap_ST_fsm_state3 : begin
            ap_NS_fsm = ap_ST_fsm_state4;
        end
        ap_ST_fsm_state4 : begin
            ap_NS_fsm = ap_ST_fsm_state5;
        end
        ap_ST_fsm_state5 : begin
            ap_NS_fsm = ap_ST_fsm_state6;
        end
        ap_ST_fsm_state6 : begin
            ap_NS_fsm = ap_ST_fsm_state7;
        end
        ap_ST_fsm_state7 : begin
            ap_NS_fsm = ap_ST_fsm_state2;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign accum_in_address0 = zext_ln81_fu_80_p1;

assign add_ln81_fu_74_p2 = (i_1_1_reg_44 + 4'd1);

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state7 = ap_CS_fsm[32'd6];

always @ (*) begin
    ap_block_state1 = ((ap_done_reg == 1'b1) | (ap_start == 1'b0));
end

assign icmp_ln81_fu_85_p2 = ((i_1_1_reg_44 == 4'd8) ? 1'b1 : 1'b0);

assign zext_ln81_fu_80_p1 = i_1_1_reg_44;

endmodule //td_fused_top_tdf5_accum_2
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf5_adjust (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        sums_read,
        adjustments_address0,
        adjustments_ce0,
        adjustments_q0,
        input_indices_23_dout,
        input_indices_23_empty_n,
        input_indices_23_read,
        ap_return
);

parameter    ap_ST_fsm_state1 = 17'd1;
parameter    ap_ST_fsm_state2 = 17'd2;
parameter    ap_ST_fsm_state3 = 17'd4;
parameter    ap_ST_fsm_state4 = 17'd8;
parameter    ap_ST_fsm_state5 = 17'd16;
parameter    ap_ST_fsm_state6 = 17'd32;
parameter    ap_ST_fsm_state7 = 17'd64;
parameter    ap_ST_fsm_state8 = 17'd128;
parameter    ap_ST_fsm_state9 = 17'd256;
parameter    ap_ST_fsm_state10 = 17'd512;
parameter    ap_ST_fsm_state11 = 17'd1024;
parameter    ap_ST_fsm_state12 = 17'd2048;
parameter    ap_ST_fsm_state13 = 17'd4096;
parameter    ap_ST_fsm_state14 = 17'd8192;
parameter    ap_ST_fsm_state15 = 17'd16384;
parameter    ap_ST_fsm_state16 = 17'd32768;
parameter    ap_ST_fsm_state17 = 17'd65536;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
input  [15:0] sums_read;
output  [6:0] adjustments_address0;
output   adjustments_ce0;
input  [47:0] adjustments_q0;
input  [6:0] input_indices_23_dout;
input   input_indices_23_empty_n;
output   input_indices_23_read;
output  [15:0] ap_return;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg adjustments_ce0;
reg input_indices_23_read;

reg    ap_done_reg;
  reg   [16:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    input_indices_23_blk_n;
wire    ap_CS_fsm_state4;
reg   [15:0] tmp_42_i_i_reg_167;
reg   [15:0] tmp_43_i_i_reg_172;
wire   [15:0] grp_fu_81_p2;
reg   [15:0] sub_i_i_i_reg_177;
wire    ap_CS_fsm_state8;
wire    ap_CS_fsm_state9;
wire   [15:0] grp_fu_86_p2;
reg   [15:0] mul_i_i_i_reg_187;
wire    ap_CS_fsm_state12;
wire    ap_CS_fsm_state13;
wire   [63:0] zext_ln220_fu_90_p1;
reg    ap_block_state1;
wire    ap_CS_fsm_state2;
wire    ap_CS_fsm_state3;
wire   [15:0] grp_fu_77_p1;
wire   [15:0] grp_fu_81_p1;
wire   [15:0] grp_fu_86_p1;
wire   [15:0] trunc_ln220_fu_95_p1;
wire   [15:0] grp_fu_77_p2;
wire    ap_CS_fsm_state17;
wire   [15:0] bitcast_ln648_fu_132_p1;
wire   [0:0] tmp_fu_136_p3;
reg   [16:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 17'd1;
end

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U305(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(mul_i_i_i_reg_187),
    .din1(grp_fu_77_p1),
    .dout(grp_fu_77_p2)
);

td_fused_top_hsub_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hsub_16ns_16ns_16_5_full_dsp_1_U306(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(sums_read),
    .din1(grp_fu_81_p1),
    .dout(grp_fu_81_p2)
);

td_fused_top_hmul_16ns_16ns_16_4_max_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hmul_16ns_16ns_16_4_max_dsp_1_U307(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(sub_i_i_i_reg_177),
    .din1(grp_fu_86_p1),
    .dout(grp_fu_86_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state17)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state12)) begin
        mul_i_i_i_reg_187 <= grp_fu_86_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state8)) begin
        sub_i_i_i_reg_177 <= grp_fu_81_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        tmp_42_i_i_reg_167 <= {{adjustments_q0[31:16]}};
        tmp_43_i_i_reg_172 <= {{adjustments_q0[47:32]}};
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state2) | (~((input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1)))) begin
        adjustments_ce0 = 1'b1;
    end else begin
        adjustments_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state17)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state17)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        input_indices_23_blk_n = input_indices_23_empty_n;
    end else begin
        input_indices_23_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        input_indices_23_read = 1'b1;
    end else begin
        input_indices_23_read = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_state2 : begin
            ap_NS_fsm = ap_ST_fsm_state3;
        end
        ap_ST_fsm_state3 : begin
            ap_NS_fsm = ap_ST_fsm_state4;
        end
        ap_ST_fsm_state4 : begin
            ap_NS_fsm = ap_ST_fsm_state5;
        end
        ap_ST_fsm_state5 : begin
            ap_NS_fsm = ap_ST_fsm_state6;
        end
        ap_ST_fsm_state6 : begin
            ap_NS_fsm = ap_ST_fsm_state7;
        end
        ap_ST_fsm_state7 : begin
            ap_NS_fsm = ap_ST_fsm_state8;
        end
        ap_ST_fsm_state8 : begin
            ap_NS_fsm = ap_ST_fsm_state9;
        end
        ap_ST_fsm_state9 : begin
            ap_NS_fsm = ap_ST_fsm_state10;
        end
        ap_ST_fsm_state10 : begin
            ap_NS_fsm = ap_ST_fsm_state11;
        end
        ap_ST_fsm_state11 : begin
            ap_NS_fsm = ap_ST_fsm_state12;
        end
        ap_ST_fsm_state12 : begin
            ap_NS_fsm = ap_ST_fsm_state13;
        end
        ap_ST_fsm_state13 : begin
            ap_NS_fsm = ap_ST_fsm_state14;
        end
        ap_ST_fsm_state14 : begin
            ap_NS_fsm = ap_ST_fsm_state15;
        end
        ap_ST_fsm_state15 : begin
            ap_NS_fsm = ap_ST_fsm_state16;
        end
        ap_ST_fsm_state16 : begin
            ap_NS_fsm = ap_ST_fsm_state17;
        end
        ap_ST_fsm_state17 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign adjustments_address0 = zext_ln220_fu_90_p1;

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state12 = ap_CS_fsm[32'd11];

assign ap_CS_fsm_state13 = ap_CS_fsm[32'd12];

assign ap_CS_fsm_state17 = ap_CS_fsm[32'd16];

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

assign ap_CS_fsm_state8 = ap_CS_fsm[32'd7];

assign ap_CS_fsm_state9 = ap_CS_fsm[32'd8];

always @ (*) begin
    ap_block_state1 = ((input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0));
end

assign ap_return = ((tmp_fu_136_p3[0:0] == 1'b1) ? 16'd0 : grp_fu_77_p2);

assign bitcast_ln648_fu_132_p1 = grp_fu_77_p2;

assign grp_fu_77_p1 = tmp_43_i_i_reg_172;

assign grp_fu_81_p1 = trunc_ln220_fu_95_p1;

assign grp_fu_86_p1 = tmp_42_i_i_reg_167;

assign tmp_fu_136_p3 = bitcast_ln648_fu_132_p1[32'd15];

assign trunc_ln220_fu_95_p1 = adjustments_q0[15:0];

assign zext_ln220_fu_90_p1 = input_indices_23_dout;

endmodule //td_fused_top_tdf5_adjust
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf5_dot_product (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        ifmap_vec_address0,
        ifmap_vec_ce0,
        ifmap_vec_q0,
        weight_vecs_0_address0,
        weight_vecs_0_ce0,
        weight_vecs_0_q0,
        products_0_address0,
        products_0_ce0,
        products_0_we0,
        products_0_d0
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state10 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [7:0] ifmap_vec_address0;
output   ifmap_vec_ce0;
input  [15:0] ifmap_vec_q0;
output  [7:0] weight_vecs_0_address0;
output   weight_vecs_0_ce0;
input  [15:0] weight_vecs_0_q0;
output  [7:0] products_0_address0;
output   products_0_ce0;
output   products_0_we0;
output  [15:0] products_0_d0;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg ifmap_vec_ce0;
reg weight_vecs_0_ce0;
reg products_0_ce0;
reg products_0_we0;

reg    ap_done_reg;
  reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg   [7:0] indvar_flatten17_reg_97;
reg   [6:0] indvar_flatten_reg_108;
reg   [1:0] jj_reg_119;
reg   [4:0] ic_reg_131;
reg   [1:0] ii_reg_142;
wire   [7:0] add_ln147_3_fu_157_p2;
wire    ap_CS_fsm_pp0_stage0;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
wire    ap_block_state4_pp0_stage0_iter2;
wire    ap_block_state5_pp0_stage0_iter3;
wire    ap_block_state6_pp0_stage0_iter4;
wire    ap_block_state7_pp0_stage0_iter5;
wire    ap_block_state8_pp0_stage0_iter6;
wire    ap_block_state9_pp0_stage0_iter7;
wire    ap_block_pp0_stage0_11001;
wire   [0:0] icmp_ln147_fu_163_p2;
reg   [0:0] icmp_ln147_reg_408;
reg   [0:0] icmp_ln147_reg_408_pp0_iter1_reg;
reg   [0:0] icmp_ln147_reg_408_pp0_iter2_reg;
reg   [0:0] icmp_ln147_reg_408_pp0_iter3_reg;
reg   [0:0] icmp_ln147_reg_408_pp0_iter4_reg;
reg   [0:0] icmp_ln147_reg_408_pp0_iter5_reg;
reg   [0:0] icmp_ln147_reg_408_pp0_iter6_reg;
wire   [0:0] icmp_ln148_fu_169_p2;
reg   [0:0] icmp_ln148_reg_412;
wire   [0:0] and_ln147_fu_195_p2;
reg   [0:0] and_ln147_reg_419;
wire   [1:0] add_ln148_fu_201_p2;
reg   [1:0] add_ln148_reg_424;
wire   [4:0] select_ln148_fu_213_p3;
reg   [4:0] select_ln148_reg_429;
wire   [1:0] select_ln148_7_fu_221_p3;
reg   [1:0] select_ln148_7_reg_434;
wire   [3:0] trunc_ln150_fu_229_p1;
reg   [3:0] trunc_ln150_reg_440;
reg   [3:0] trunc_ln150_reg_440_pp0_iter1_reg;
reg   [3:0] trunc_ln150_reg_440_pp0_iter2_reg;
reg   [3:0] trunc_ln150_reg_440_pp0_iter3_reg;
reg   [3:0] trunc_ln150_reg_440_pp0_iter4_reg;
reg   [3:0] trunc_ln150_reg_440_pp0_iter5_reg;
reg   [3:0] trunc_ln150_reg_440_pp0_iter6_reg;
wire   [4:0] add_ln149_fu_233_p2;
wire   [6:0] select_ln148_9_fu_245_p3;
wire   [1:0] select_ln147_8_fu_287_p3;
reg   [1:0] select_ln147_8_reg_455;
reg    ap_enable_reg_pp0_iter1;
wire   [3:0] select_ln148_8_fu_370_p3;
reg   [3:0] select_ln148_8_reg_460;
reg   [3:0] select_ln148_8_reg_460_pp0_iter2_reg;
reg   [3:0] select_ln148_8_reg_460_pp0_iter3_reg;
reg   [3:0] select_ln148_8_reg_460_pp0_iter4_reg;
reg   [3:0] select_ln148_8_reg_460_pp0_iter5_reg;
reg   [3:0] select_ln148_8_reg_460_pp0_iter6_reg;
reg   [15:0] ifmap_vec_load_reg_475;
reg   [15:0] weight_vecs_0_load_reg_480;
wire   [15:0] grp_fu_153_p2;
reg   [15:0] mul_reg_485;
reg    ap_block_state1;
wire    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_flush_enable;
reg    ap_enable_reg_pp0_iter2;
reg    ap_condition_pp0_exit_iter1_state3;
reg    ap_enable_reg_pp0_iter3;
reg    ap_enable_reg_pp0_iter4;
reg    ap_enable_reg_pp0_iter5;
reg    ap_enable_reg_pp0_iter6;
reg    ap_enable_reg_pp0_iter7;
reg   [1:0] ap_phi_mux_jj_phi_fu_123_p4;
wire    ap_block_pp0_stage0;
reg   [1:0] ap_phi_mux_ii_phi_fu_146_p4;
wire   [63:0] p_cast25_fu_386_p1;
wire   [63:0] idxprom30_fu_398_p1;
wire   [0:0] icmp_ln149_fu_189_p2;
wire   [0:0] xor_ln147_fu_183_p2;
wire   [1:0] select_ln147_fu_175_p3;
wire   [0:0] or_ln148_fu_207_p2;
wire   [6:0] add_ln148_3_fu_239_p2;
wire   [3:0] shl_ln_fu_257_p3;
wire   [3:0] zext_ln150_fu_253_p1;
wire   [3:0] sub_ln150_fu_265_p2;
wire   [3:0] zext_ln150_3_fu_271_p1;
wire   [1:0] add_ln147_fu_281_p2;
wire   [3:0] tmp_fu_298_p3;
wire   [3:0] select_ln147_10_cast_fu_294_p1;
wire   [3:0] shl_ln150_mid1_fu_316_p3;
wire   [3:0] zext_ln150_6_fu_312_p1;
wire   [3:0] sub_ln150_3_fu_324_p2;
wire   [3:0] add_ln150_fu_275_p2;
wire   [3:0] empty_88_fu_306_p2;
wire   [3:0] select_ln148_9_cast_fu_344_p1;
wire   [3:0] empty_89_fu_347_p2;
wire   [3:0] select_ln147_9_fu_330_p3;
wire   [3:0] zext_ln150_7_fu_361_p1;
wire   [3:0] add_ln150_3_fu_364_p2;
wire   [3:0] select_ln147_10_fu_337_p3;
wire   [7:0] tmp_78_cast_fu_353_p3;
wire   [7:0] select_ln148_cast_fu_377_p1;
wire   [7:0] empty_90_fu_380_p2;
wire   [7:0] p_fu_392_p3;
wire    ap_CS_fsm_state10;
reg   [2:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
#0 ap_enable_reg_pp0_iter4 = 1'b0;
#0 ap_enable_reg_pp0_iter5 = 1'b0;
#0 ap_enable_reg_pp0_iter6 = 1'b0;
#0 ap_enable_reg_pp0_iter7 = 1'b0;
end

td_fused_top_hmul_16ns_16ns_16_4_max_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hmul_16ns_16ns_16_4_max_dsp_1_U293(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(ifmap_vec_load_reg_475),
    .din1(weight_vecs_0_load_reg_480),
    .dout(grp_fu_153_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state10)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if ((1'b1 == ap_condition_pp0_flush_enable)) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            if ((1'b1 == ap_condition_pp0_exit_iter1_state3)) begin
                ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter0;
            end else if ((1'b1 == 1'b1)) begin
                ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
            end
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter4 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter5 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter5 <= ap_enable_reg_pp0_iter4;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter6 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter6 <= ap_enable_reg_pp0_iter5;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter7 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter7 <= ap_enable_reg_pp0_iter6;
        end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter7 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_fu_163_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ic_reg_131 <= add_ln149_fu_233_p2;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ic_reg_131 <= 5'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_reg_408_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        ii_reg_142 <= select_ln147_8_reg_455;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ii_reg_142 <= 2'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_fu_163_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        indvar_flatten17_reg_97 <= add_ln147_3_fu_157_p2;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indvar_flatten17_reg_97 <= 8'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_fu_163_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        indvar_flatten_reg_108 <= select_ln148_9_fu_245_p3;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indvar_flatten_reg_108 <= 7'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_reg_408 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        jj_reg_119 <= select_ln148_7_reg_434;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        jj_reg_119 <= 2'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_fu_163_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        add_ln148_reg_424 <= add_ln148_fu_201_p2;
        and_ln147_reg_419 <= and_ln147_fu_195_p2;
        icmp_ln148_reg_412 <= icmp_ln148_fu_169_p2;
        select_ln148_reg_429 <= select_ln148_fu_213_p3;
        trunc_ln150_reg_440 <= trunc_ln150_fu_229_p1;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln147_reg_408 <= icmp_ln147_fu_163_p2;
        icmp_ln147_reg_408_pp0_iter1_reg <= icmp_ln147_reg_408;
        trunc_ln150_reg_440_pp0_iter1_reg <= trunc_ln150_reg_440;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        icmp_ln147_reg_408_pp0_iter2_reg <= icmp_ln147_reg_408_pp0_iter1_reg;
        icmp_ln147_reg_408_pp0_iter3_reg <= icmp_ln147_reg_408_pp0_iter2_reg;
        icmp_ln147_reg_408_pp0_iter4_reg <= icmp_ln147_reg_408_pp0_iter3_reg;
        icmp_ln147_reg_408_pp0_iter5_reg <= icmp_ln147_reg_408_pp0_iter4_reg;
        icmp_ln147_reg_408_pp0_iter6_reg <= icmp_ln147_reg_408_pp0_iter5_reg;
        select_ln148_8_reg_460_pp0_iter2_reg <= select_ln148_8_reg_460;
        select_ln148_8_reg_460_pp0_iter3_reg <= select_ln148_8_reg_460_pp0_iter2_reg;
        select_ln148_8_reg_460_pp0_iter4_reg <= select_ln148_8_reg_460_pp0_iter3_reg;
        select_ln148_8_reg_460_pp0_iter5_reg <= select_ln148_8_reg_460_pp0_iter4_reg;
        select_ln148_8_reg_460_pp0_iter6_reg <= select_ln148_8_reg_460_pp0_iter5_reg;
        trunc_ln150_reg_440_pp0_iter2_reg <= trunc_ln150_reg_440_pp0_iter1_reg;
        trunc_ln150_reg_440_pp0_iter3_reg <= trunc_ln150_reg_440_pp0_iter2_reg;
        trunc_ln150_reg_440_pp0_iter4_reg <= trunc_ln150_reg_440_pp0_iter3_reg;
        trunc_ln150_reg_440_pp0_iter5_reg <= trunc_ln150_reg_440_pp0_iter4_reg;
        trunc_ln150_reg_440_pp0_iter6_reg <= trunc_ln150_reg_440_pp0_iter5_reg;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_reg_408_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        ifmap_vec_load_reg_475 <= ifmap_vec_q0;
        weight_vecs_0_load_reg_480 <= weight_vecs_0_q0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_reg_408_pp0_iter5_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        mul_reg_485 <= grp_fu_153_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_reg_408 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        select_ln147_8_reg_455 <= select_ln147_8_fu_287_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_fu_163_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        select_ln148_7_reg_434 <= select_ln148_7_fu_221_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_reg_408 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        select_ln148_8_reg_460 <= select_ln148_8_fu_370_p3;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_condition_pp0_exit_iter1_state3 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter1_state3 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln147_fu_163_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_condition_pp0_flush_enable = 1'b1;
    end else begin
        ap_condition_pp0_flush_enable = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state10)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter7 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln147_reg_408_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        ap_phi_mux_ii_phi_fu_146_p4 = select_ln147_8_reg_455;
    end else begin
        ap_phi_mux_ii_phi_fu_146_p4 = ii_reg_142;
    end
end

always @ (*) begin
    if (((icmp_ln147_reg_408 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_jj_phi_fu_123_p4 = select_ln148_7_reg_434;
    end else begin
        ap_phi_mux_jj_phi_fu_123_p4 = jj_reg_119;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state10)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ifmap_vec_ce0 = 1'b1;
    end else begin
        ifmap_vec_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter7 == 1'b1))) begin
        products_0_ce0 = 1'b1;
    end else begin
        products_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln147_reg_408_pp0_iter6_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter7 == 1'b1))) begin
        products_0_we0 = 1'b1;
    end else begin
        products_0_we0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        weight_vecs_0_ce0 = 1'b1;
    end else begin
        weight_vecs_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((~((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b1)) & ~((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter7 == 1'b1) & (ap_enable_reg_pp0_iter6 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if ((((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter7 == 1'b1) & (ap_enable_reg_pp0_iter6 == 1'b0)) | ((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b1)))) begin
                ap_NS_fsm = ap_ST_fsm_state10;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state10 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln147_3_fu_157_p2 = (indvar_flatten17_reg_97 + 8'd1);

assign add_ln147_fu_281_p2 = (ap_phi_mux_ii_phi_fu_146_p4 + 2'd1);

assign add_ln148_3_fu_239_p2 = (indvar_flatten_reg_108 + 7'd1);

assign add_ln148_fu_201_p2 = (select_ln147_fu_175_p3 + 2'd1);

assign add_ln149_fu_233_p2 = (select_ln148_fu_213_p3 + 5'd1);

assign add_ln150_3_fu_364_p2 = (select_ln147_9_fu_330_p3 + zext_ln150_7_fu_361_p1);

assign add_ln150_fu_275_p2 = (sub_ln150_fu_265_p2 + zext_ln150_3_fu_271_p1);

assign and_ln147_fu_195_p2 = (xor_ln147_fu_183_p2 & icmp_ln149_fu_189_p2);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state10 = ap_CS_fsm[32'd2];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (ap_done_reg == 1'b1));
end

assign ap_block_state2_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter4 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage0_iter5 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage0_iter6 = ~(1'b1 == 1'b1);

assign ap_block_state9_pp0_stage0_iter7 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign empty_88_fu_306_p2 = (tmp_fu_298_p3 - select_ln147_10_cast_fu_294_p1);

assign empty_89_fu_347_p2 = (empty_88_fu_306_p2 + select_ln148_9_cast_fu_344_p1);

assign empty_90_fu_380_p2 = (tmp_78_cast_fu_353_p3 + select_ln148_cast_fu_377_p1);

assign icmp_ln147_fu_163_p2 = ((indvar_flatten17_reg_97 == 8'd144) ? 1'b1 : 1'b0);

assign icmp_ln148_fu_169_p2 = ((indvar_flatten_reg_108 == 7'd48) ? 1'b1 : 1'b0);

assign icmp_ln149_fu_189_p2 = ((ic_reg_131 == 5'd16) ? 1'b1 : 1'b0);

assign idxprom30_fu_398_p1 = p_fu_392_p3;

assign ifmap_vec_address0 = p_cast25_fu_386_p1;

assign or_ln148_fu_207_p2 = (icmp_ln148_fu_169_p2 | and_ln147_fu_195_p2);

assign p_cast25_fu_386_p1 = empty_90_fu_380_p2;

assign p_fu_392_p3 = {{select_ln148_8_reg_460_pp0_iter6_reg}, {trunc_ln150_reg_440_pp0_iter6_reg}};

assign products_0_address0 = idxprom30_fu_398_p1;

assign products_0_d0 = mul_reg_485;

assign select_ln147_10_cast_fu_294_p1 = select_ln147_8_fu_287_p3;

assign select_ln147_10_fu_337_p3 = ((icmp_ln148_reg_412[0:0] == 1'b1) ? sub_ln150_3_fu_324_p2 : add_ln150_fu_275_p2);

assign select_ln147_8_fu_287_p3 = ((icmp_ln148_reg_412[0:0] == 1'b1) ? add_ln147_fu_281_p2 : ap_phi_mux_ii_phi_fu_146_p4);

assign select_ln147_9_fu_330_p3 = ((icmp_ln148_reg_412[0:0] == 1'b1) ? sub_ln150_3_fu_324_p2 : sub_ln150_fu_265_p2);

assign select_ln147_fu_175_p3 = ((icmp_ln148_fu_169_p2[0:0] == 1'b1) ? 2'd0 : ap_phi_mux_jj_phi_fu_123_p4);

assign select_ln148_7_fu_221_p3 = ((and_ln147_fu_195_p2[0:0] == 1'b1) ? add_ln148_fu_201_p2 : select_ln147_fu_175_p3);

assign select_ln148_8_fu_370_p3 = ((and_ln147_reg_419[0:0] == 1'b1) ? add_ln150_3_fu_364_p2 : select_ln147_10_fu_337_p3);

assign select_ln148_9_cast_fu_344_p1 = select_ln148_7_reg_434;

assign select_ln148_9_fu_245_p3 = ((icmp_ln148_fu_169_p2[0:0] == 1'b1) ? 7'd1 : add_ln148_3_fu_239_p2);

assign select_ln148_cast_fu_377_p1 = select_ln148_reg_429;

assign select_ln148_fu_213_p3 = ((or_ln148_fu_207_p2[0:0] == 1'b1) ? 5'd0 : ic_reg_131);

assign shl_ln150_mid1_fu_316_p3 = {{add_ln147_fu_281_p2}, {2'd0}};

assign shl_ln_fu_257_p3 = {{ap_phi_mux_ii_phi_fu_146_p4}, {2'd0}};

assign sub_ln150_3_fu_324_p2 = (shl_ln150_mid1_fu_316_p3 - zext_ln150_6_fu_312_p1);

assign sub_ln150_fu_265_p2 = (shl_ln_fu_257_p3 - zext_ln150_fu_253_p1);

assign tmp_78_cast_fu_353_p3 = {{empty_89_fu_347_p2}, {4'd0}};

assign tmp_fu_298_p3 = {{select_ln147_8_fu_287_p3}, {2'd0}};

assign trunc_ln150_fu_229_p1 = select_ln148_fu_213_p3[3:0];

assign weight_vecs_0_address0 = p_cast25_fu_386_p1;

assign xor_ln147_fu_183_p2 = (icmp_ln148_fu_169_p2 ^ 1'd1);

assign zext_ln150_3_fu_271_p1 = jj_reg_119;

assign zext_ln150_6_fu_312_p1 = add_ln147_fu_281_p2;

assign zext_ln150_7_fu_361_p1 = add_ln148_reg_424;

assign zext_ln150_fu_253_p1 = ap_phi_mux_ii_phi_fu_146_p4;

endmodule //td_fused_top_tdf5_dot_product
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf5_get_next_ijk (
        ap_clk,
        ap_rst,
        ap_start,
        start_full_n,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        start_out,
        start_write,
        input_indices_2_out_din,
        input_indices_2_out_full_n,
        input_indices_2_out_write,
        input_indices_2_out1_din,
        input_indices_2_out1_full_n,
        input_indices_2_out1_write,
        output_indices_0_din,
        output_indices_0_full_n,
        output_indices_0_write,
        output_indices_1_din,
        output_indices_1_full_n,
        output_indices_1_write,
        resetMaximum_din,
        resetMaximum_full_n,
        resetMaximum_write,
        storeOutput_din,
        storeOutput_full_n,
        storeOutput_write,
        ap_return_0,
        ap_return_1
);

parameter    ap_ST_fsm_state1 = 1'd1;

input   ap_clk;
input   ap_rst;
input   ap_start;
input   start_full_n;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output   start_out;
output   start_write;
output  [6:0] input_indices_2_out_din;
input   input_indices_2_out_full_n;
output   input_indices_2_out_write;
output  [6:0] input_indices_2_out1_din;
input   input_indices_2_out1_full_n;
output   input_indices_2_out1_write;
output  [4:0] output_indices_0_din;
input   output_indices_0_full_n;
output   output_indices_0_write;
output  [9:0] output_indices_1_din;
input   output_indices_1_full_n;
output   output_indices_1_write;
output   resetMaximum_din;
input   resetMaximum_full_n;
output   resetMaximum_write;
output   storeOutput_din;
input   storeOutput_full_n;
output   storeOutput_write;
output  [15:0] ap_return_0;
output  [15:0] ap_return_1;

reg ap_done;
reg ap_idle;
reg start_write;
reg input_indices_2_out_write;
reg input_indices_2_out1_write;
reg output_indices_0_write;
reg output_indices_1_write;
reg resetMaximum_write;
reg storeOutput_write;

reg    real_start;
reg    start_once_reg;
reg    ap_done_reg;
  reg   [0:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    internal_ap_ready;
reg   [1:0] i_p_1;
reg   [1:0] j_p_1;
reg   [15:0] i_3;
reg   [15:0] j_3;
reg   [15:0] k_3;
reg   [15:0] i_out_1;
reg   [15:0] j_out_1;
reg    input_indices_2_out_blk_n;
reg    input_indices_2_out1_blk_n;
reg    output_indices_0_blk_n;
reg    output_indices_1_blk_n;
reg    resetMaximum_blk_n;
reg    storeOutput_blk_n;
wire   [1:0] select_ln142_fu_338_p3;
reg    ap_block_state1;
wire   [0:0] or_ln142_fu_312_p2;
wire   [1:0] select_ln142_5_fu_346_p3;
wire   [15:0] select_ln147_fu_278_p3;
wire   [0:0] and_ln142_2_fu_306_p2;
wire   [15:0] select_ln142_6_fu_360_p3;
wire   [0:0] and_ln132_fu_354_p2;
wire   [15:0] select_ln142_7_fu_388_p3;
wire   [0:0] and_ln135_fu_294_p2;
wire   [15:0] select_ln147_2_fu_286_p3;
wire   [15:0] select_ln142_8_fu_396_p3;
wire   [6:0] trunc_ln128_fu_182_p1;
wire   [1:0] or_ln124_fu_126_p2;
wire   [0:0] icmp_ln125_fu_139_p2;
wire   [0:0] icmp_ln125_2_fu_145_p2;
wire   [15:0] zext_ln126_fu_114_p1;
wire   [15:0] zext_ln127_fu_122_p1;
wire   [1:0] add_ln131_fu_206_p2;
wire   [1:0] add_ln134_fu_218_p2;
wire   [15:0] add_ln137_fu_230_p2;
wire   [15:0] add_ln141_fu_248_p2;
wire   [15:0] add_ln146_fu_266_p2;
wire   [0:0] icmp_ln147_fu_272_p2;
wire   [15:0] add_ln145_fu_260_p2;
wire   [0:0] icmp_ln132_fu_212_p2;
wire   [0:0] icmp_ln135_fu_224_p2;
wire   [0:0] icmp_ln138_fu_236_p2;
wire   [0:0] icmp_ln142_fu_254_p2;
wire   [0:0] and_ln142_fu_300_p2;
wire   [0:0] xor_ln135_fu_318_p2;
wire   [0:0] and_ln135_2_fu_324_p2;
wire   [1:0] select_ln135_fu_330_p3;
wire   [15:0] add_ln140_fu_242_p2;
wire   [0:0] xor_ln138_fu_368_p2;
wire   [0:0] and_ln138_fu_374_p2;
wire   [15:0] select_ln138_fu_380_p3;
wire   [15:0] add_ln126_fu_162_p2;
wire   [15:0] add_ln127_fu_172_p2;
reg   [0:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 start_once_reg = 1'b0;
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 1'd1;
#0 i_p_1 = 2'd0;
#0 j_p_1 = 2'd0;
#0 i_3 = 16'd0;
#0 j_3 = 16'd0;
#0 k_3 = 16'd0;
#0 i_out_1 = 16'd0;
#0 j_out_1 = 16'd0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        start_once_reg <= 1'b0;
    end else begin
        if (((real_start == 1'b1) & (internal_ap_ready == 1'b0))) begin
            start_once_reg <= 1'b1;
        end else if ((internal_ap_ready == 1'b1)) begin
            start_once_reg <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1) & (1'd1 == and_ln142_2_fu_306_p2))) begin
        i_3 <= select_ln147_fu_278_p3;
        i_out_1 <= select_ln147_2_fu_286_p3;
    end
end

always @ (posedge ap_clk) begin
    if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (or_ln142_fu_312_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1))) begin
        i_p_1 <= select_ln142_fu_338_p3;
    end
end

always @ (posedge ap_clk) begin
    if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1) & (1'd1 == and_ln132_fu_354_p2))) begin
        j_3 <= select_ln142_6_fu_360_p3;
        j_out_1 <= select_ln142_8_fu_396_p3;
    end
end

always @ (posedge ap_clk) begin
    if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        j_p_1 <= select_ln142_5_fu_346_p3;
    end
end

always @ (posedge ap_clk) begin
    if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1) & (1'd1 == and_ln135_fu_294_p2))) begin
        k_3 <= select_ln142_7_fu_388_p3;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((real_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        input_indices_2_out1_blk_n = input_indices_2_out1_full_n;
    end else begin
        input_indices_2_out1_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        input_indices_2_out1_write = 1'b1;
    end else begin
        input_indices_2_out1_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        input_indices_2_out_blk_n = input_indices_2_out_full_n;
    end else begin
        input_indices_2_out_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        input_indices_2_out_write = 1'b1;
    end else begin
        input_indices_2_out_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        internal_ap_ready = 1'b1;
    end else begin
        internal_ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        output_indices_0_blk_n = output_indices_0_full_n;
    end else begin
        output_indices_0_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        output_indices_0_write = 1'b1;
    end else begin
        output_indices_0_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        output_indices_1_blk_n = output_indices_1_full_n;
    end else begin
        output_indices_1_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        output_indices_1_write = 1'b1;
    end else begin
        output_indices_1_write = 1'b0;
    end
end

always @ (*) begin
    if (((start_full_n == 1'b0) & (start_once_reg == 1'b0))) begin
        real_start = 1'b0;
    end else begin
        real_start = ap_start;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        resetMaximum_blk_n = resetMaximum_full_n;
    end else begin
        resetMaximum_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        resetMaximum_write = 1'b1;
    end else begin
        resetMaximum_write = 1'b0;
    end
end

always @ (*) begin
    if (((real_start == 1'b1) & (start_once_reg == 1'b0))) begin
        start_write = 1'b1;
    end else begin
        start_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        storeOutput_blk_n = storeOutput_full_n;
    end else begin
        storeOutput_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        storeOutput_write = 1'b1;
    end else begin
        storeOutput_write = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln126_fu_162_p2 = (i_3 + zext_ln126_fu_114_p1);

assign add_ln127_fu_172_p2 = (j_3 + zext_ln127_fu_122_p1);

assign add_ln131_fu_206_p2 = (j_p_1 + 2'd1);

assign add_ln134_fu_218_p2 = (i_p_1 + 2'd1);

assign add_ln137_fu_230_p2 = (k_3 + 16'd1);

assign add_ln140_fu_242_p2 = (j_3 + 16'd2);

assign add_ln141_fu_248_p2 = (j_out_1 + 16'd1);

assign add_ln145_fu_260_p2 = (i_3 + 16'd2);

assign add_ln146_fu_266_p2 = (i_out_1 + 16'd1);

assign and_ln132_fu_354_p2 = (icmp_ln138_fu_236_p2 & and_ln135_fu_294_p2);

assign and_ln135_2_fu_324_p2 = (xor_ln135_fu_318_p2 & icmp_ln132_fu_212_p2);

assign and_ln135_fu_294_p2 = (icmp_ln135_fu_224_p2 & icmp_ln132_fu_212_p2);

assign and_ln138_fu_374_p2 = (xor_ln138_fu_368_p2 & and_ln135_fu_294_p2);

assign and_ln142_2_fu_306_p2 = (and_ln142_fu_300_p2 & and_ln135_fu_294_p2);

assign and_ln142_fu_300_p2 = (icmp_ln142_fu_254_p2 & icmp_ln138_fu_236_p2);

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

always @ (*) begin
    ap_block_state1 = ((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1));
end

assign ap_ready = internal_ap_ready;

assign ap_return_0 = add_ln126_fu_162_p2;

assign ap_return_1 = add_ln127_fu_172_p2;

assign icmp_ln125_2_fu_145_p2 = ((j_p_1 == 2'd1) ? 1'b1 : 1'b0);

assign icmp_ln125_fu_139_p2 = ((i_p_1 == 2'd1) ? 1'b1 : 1'b0);

assign icmp_ln132_fu_212_p2 = ((add_ln131_fu_206_p2 == 2'd2) ? 1'b1 : 1'b0);

assign icmp_ln135_fu_224_p2 = ((add_ln134_fu_218_p2 == 2'd2) ? 1'b1 : 1'b0);

assign icmp_ln138_fu_236_p2 = ((add_ln137_fu_230_p2 == 16'd128) ? 1'b1 : 1'b0);

assign icmp_ln142_fu_254_p2 = ((add_ln141_fu_248_p2 == 16'd28) ? 1'b1 : 1'b0);

assign icmp_ln147_fu_272_p2 = ((add_ln146_fu_266_p2 == 16'd28) ? 1'b1 : 1'b0);

assign input_indices_2_out1_din = trunc_ln128_fu_182_p1;

assign input_indices_2_out_din = trunc_ln128_fu_182_p1;

assign or_ln124_fu_126_p2 = (j_p_1 | i_p_1);

assign or_ln142_fu_312_p2 = (icmp_ln132_fu_212_p2 | and_ln142_2_fu_306_p2);

assign output_indices_0_din = i_out_1[4:0];

assign output_indices_1_din = j_out_1[9:0];

assign resetMaximum_din = ((or_ln124_fu_126_p2 == 2'd0) ? 1'b1 : 1'b0);

assign select_ln135_fu_330_p3 = ((and_ln135_2_fu_324_p2[0:0] == 1'b1) ? add_ln134_fu_218_p2 : 2'd0);

assign select_ln138_fu_380_p3 = ((and_ln138_fu_374_p2[0:0] == 1'b1) ? add_ln137_fu_230_p2 : 16'd0);

assign select_ln142_5_fu_346_p3 = ((or_ln142_fu_312_p2[0:0] == 1'b1) ? 2'd0 : add_ln131_fu_206_p2);

assign select_ln142_6_fu_360_p3 = ((and_ln142_2_fu_306_p2[0:0] == 1'b1) ? 16'd0 : add_ln140_fu_242_p2);

assign select_ln142_7_fu_388_p3 = ((and_ln142_2_fu_306_p2[0:0] == 1'b1) ? 16'd0 : select_ln138_fu_380_p3);

assign select_ln142_8_fu_396_p3 = ((and_ln142_2_fu_306_p2[0:0] == 1'b1) ? 16'd0 : add_ln141_fu_248_p2);

assign select_ln142_fu_338_p3 = ((and_ln142_2_fu_306_p2[0:0] == 1'b1) ? 2'd0 : select_ln135_fu_330_p3);

assign select_ln147_2_fu_286_p3 = ((icmp_ln147_fu_272_p2[0:0] == 1'b1) ? 16'd0 : add_ln146_fu_266_p2);

assign select_ln147_fu_278_p3 = ((icmp_ln147_fu_272_p2[0:0] == 1'b1) ? 16'd0 : add_ln145_fu_260_p2);

assign start_out = real_start;

assign storeOutput_din = (icmp_ln125_fu_139_p2 & icmp_ln125_2_fu_145_p2);

assign trunc_ln128_fu_182_p1 = k_3[6:0];

assign xor_ln135_fu_318_p2 = (icmp_ln135_fu_224_p2 ^ 1'd1);

assign xor_ln138_fu_368_p2 = (icmp_ln138_fu_236_p2 ^ 1'd1);

assign zext_ln126_fu_114_p1 = i_p_1;

assign zext_ln127_fu_122_p1 = j_p_1;

endmodule //td_fused_top_tdf5_get_next_ijk
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf5_poolOutputs (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        output_indices_04_dout,
        output_indices_04_empty_n,
        output_indices_04_read,
        output_indices_15_dout,
        output_indices_15_empty_n,
        output_indices_15_read,
        resetMaximum6_dout,
        resetMaximum6_empty_n,
        resetMaximum6_read,
        storeOutput7_dout,
        storeOutput7_empty_n,
        storeOutput7_read,
        p_read,
        out_data_address1,
        out_data_ce1,
        out_data_we1,
        out_data_d1
);

parameter    ap_ST_fsm_state1 = 4'd1;
parameter    ap_ST_fsm_state2 = 4'd2;
parameter    ap_ST_fsm_state3 = 4'd4;
parameter    ap_ST_fsm_state4 = 4'd8;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
input  [4:0] output_indices_04_dout;
input   output_indices_04_empty_n;
output   output_indices_04_read;
input  [9:0] output_indices_15_dout;
input   output_indices_15_empty_n;
output   output_indices_15_read;
input  [0:0] resetMaximum6_dout;
input   resetMaximum6_empty_n;
output   resetMaximum6_read;
input  [0:0] storeOutput7_dout;
input   storeOutput7_empty_n;
output   storeOutput7_read;
input  [15:0] p_read;
output  [14:0] out_data_address1;
output   out_data_ce1;
output   out_data_we1;
output  [63:0] out_data_d1;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg output_indices_04_read;
reg output_indices_15_read;
reg resetMaximum6_read;
reg storeOutput7_read;

reg    ap_done_reg;
  reg   [3:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg   [15:0] max_vals_5_0;
reg    output_indices_04_blk_n;
wire    ap_CS_fsm_state2;
reg    output_indices_15_blk_n;
reg    resetMaximum6_blk_n;
reg    storeOutput7_blk_n;
reg   [4:0] output_indices_04_read_reg_147;
reg   [9:0] output_indices_15_read_reg_152;
wire   [0:0] storeOutput7_read_read_fu_82_p2;
reg   [0:0] storeOutput7_read_reg_157;
wire    grp_tdf5_writeOutputs_unaligned_fu_88_ap_start;
wire    grp_tdf5_writeOutputs_unaligned_fu_88_ap_done;
wire    grp_tdf5_writeOutputs_unaligned_fu_88_ap_idle;
wire    grp_tdf5_writeOutputs_unaligned_fu_88_ap_ready;
wire   [14:0] grp_tdf5_writeOutputs_unaligned_fu_88_out_data_address1;
wire    grp_tdf5_writeOutputs_unaligned_fu_88_out_data_ce1;
wire    grp_tdf5_writeOutputs_unaligned_fu_88_out_data_we1;
wire   [63:0] grp_tdf5_writeOutputs_unaligned_fu_88_out_data_d1;
reg    grp_tdf5_writeOutputs_unaligned_fu_88_ap_start_reg;
wire    ap_CS_fsm_state3;
wire    ap_CS_fsm_state4;
reg    ap_block_state4_on_subcall_done;
wire   [15:0] select_ln24_fu_126_p3;
reg    ap_block_state2;
reg    ap_block_state1;
wire   [0:0] grp_fu_110_p2;
wire   [0:0] or_ln24_fu_120_p2;
reg    grp_fu_110_ce;
reg   [3:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 4'd1;
#0 max_vals_5_0 = 16'd0;
#0 grp_tdf5_writeOutputs_unaligned_fu_88_ap_start_reg = 1'b0;
end

td_fused_top_tdf5_writeOutputs_unaligned grp_tdf5_writeOutputs_unaligned_fu_88(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(grp_tdf5_writeOutputs_unaligned_fu_88_ap_start),
    .ap_done(grp_tdf5_writeOutputs_unaligned_fu_88_ap_done),
    .ap_idle(grp_tdf5_writeOutputs_unaligned_fu_88_ap_idle),
    .ap_ready(grp_tdf5_writeOutputs_unaligned_fu_88_ap_ready),
    .i(output_indices_04_read_reg_147),
    .j(output_indices_15_read_reg_152),
    .out_data_address1(grp_tdf5_writeOutputs_unaligned_fu_88_out_data_address1),
    .out_data_ce1(grp_tdf5_writeOutputs_unaligned_fu_88_out_data_ce1),
    .out_data_we1(grp_tdf5_writeOutputs_unaligned_fu_88_out_data_we1),
    .out_data_d1(grp_tdf5_writeOutputs_unaligned_fu_88_out_data_d1),
    .max_vals_5_0(max_vals_5_0)
);

td_fused_top_hcmp_16ns_16ns_1_2_no_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 1 ))
hcmp_16ns_16ns_1_2_no_dsp_1_U315(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(grp_fu_110_ce),
    .din0(max_vals_5_0),
    .din1(p_read),
    .opcode(5'd4),
    .dout(grp_fu_110_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_state4) & (1'b0 == ap_block_state4_on_subcall_done))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        grp_tdf5_writeOutputs_unaligned_fu_88_ap_start_reg <= 1'b0;
    end else begin
        if ((1'b1 == ap_CS_fsm_state3)) begin
            grp_tdf5_writeOutputs_unaligned_fu_88_ap_start_reg <= 1'b1;
        end else if ((grp_tdf5_writeOutputs_unaligned_fu_88_ap_ready == 1'b1)) begin
            grp_tdf5_writeOutputs_unaligned_fu_88_ap_start_reg <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((~((storeOutput7_empty_n == 1'b0) | (resetMaximum6_empty_n == 1'b0) | (output_indices_15_empty_n == 1'b0) | (output_indices_04_empty_n == 1'b0)) & (1'b1 == ap_CS_fsm_state2))) begin
        max_vals_5_0 <= select_ln24_fu_126_p3;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        output_indices_04_read_reg_147 <= output_indices_04_dout;
        output_indices_15_read_reg_152 <= output_indices_15_dout;
        storeOutput7_read_reg_157 <= storeOutput7_dout;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state4) & (1'b0 == ap_block_state4_on_subcall_done))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state4) & (1'b0 == ap_block_state4_on_subcall_done))) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1)) | (~((storeOutput7_empty_n == 1'b0) | (resetMaximum6_empty_n == 1'b0) | (output_indices_15_empty_n == 1'b0) | (output_indices_04_empty_n == 1'b0)) & (1'b1 == ap_CS_fsm_state2)))) begin
        grp_fu_110_ce = 1'b1;
    end else begin
        grp_fu_110_ce = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        output_indices_04_blk_n = output_indices_04_empty_n;
    end else begin
        output_indices_04_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((storeOutput7_empty_n == 1'b0) | (resetMaximum6_empty_n == 1'b0) | (output_indices_15_empty_n == 1'b0) | (output_indices_04_empty_n == 1'b0)) & (1'b1 == ap_CS_fsm_state2))) begin
        output_indices_04_read = 1'b1;
    end else begin
        output_indices_04_read = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        output_indices_15_blk_n = output_indices_15_empty_n;
    end else begin
        output_indices_15_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((storeOutput7_empty_n == 1'b0) | (resetMaximum6_empty_n == 1'b0) | (output_indices_15_empty_n == 1'b0) | (output_indices_04_empty_n == 1'b0)) & (1'b1 == ap_CS_fsm_state2))) begin
        output_indices_15_read = 1'b1;
    end else begin
        output_indices_15_read = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        resetMaximum6_blk_n = resetMaximum6_empty_n;
    end else begin
        resetMaximum6_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((storeOutput7_empty_n == 1'b0) | (resetMaximum6_empty_n == 1'b0) | (output_indices_15_empty_n == 1'b0) | (output_indices_04_empty_n == 1'b0)) & (1'b1 == ap_CS_fsm_state2))) begin
        resetMaximum6_read = 1'b1;
    end else begin
        resetMaximum6_read = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        storeOutput7_blk_n = storeOutput7_empty_n;
    end else begin
        storeOutput7_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((storeOutput7_empty_n == 1'b0) | (resetMaximum6_empty_n == 1'b0) | (output_indices_15_empty_n == 1'b0) | (output_indices_04_empty_n == 1'b0)) & (1'b1 == ap_CS_fsm_state2))) begin
        storeOutput7_read = 1'b1;
    end else begin
        storeOutput7_read = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_state2 : begin
            if ((~((storeOutput7_empty_n == 1'b0) | (resetMaximum6_empty_n == 1'b0) | (output_indices_15_empty_n == 1'b0) | (output_indices_04_empty_n == 1'b0)) & (storeOutput7_read_read_fu_82_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state2))) begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end else if ((~((storeOutput7_empty_n == 1'b0) | (resetMaximum6_empty_n == 1'b0) | (output_indices_15_empty_n == 1'b0) | (output_indices_04_empty_n == 1'b0)) & (storeOutput7_read_read_fu_82_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end
        end
        ap_ST_fsm_state3 : begin
            ap_NS_fsm = ap_ST_fsm_state4;
        end
        ap_ST_fsm_state4 : begin
            if (((1'b1 == ap_CS_fsm_state4) & (1'b0 == ap_block_state4_on_subcall_done))) begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (ap_done_reg == 1'b1));
end

always @ (*) begin
    ap_block_state2 = ((storeOutput7_empty_n == 1'b0) | (resetMaximum6_empty_n == 1'b0) | (output_indices_15_empty_n == 1'b0) | (output_indices_04_empty_n == 1'b0));
end

always @ (*) begin
    ap_block_state4_on_subcall_done = ((grp_tdf5_writeOutputs_unaligned_fu_88_ap_done == 1'b0) & (storeOutput7_read_reg_157 == 1'd1));
end

assign grp_tdf5_writeOutputs_unaligned_fu_88_ap_start = grp_tdf5_writeOutputs_unaligned_fu_88_ap_start_reg;

assign or_ln24_fu_120_p2 = (resetMaximum6_dout | grp_fu_110_p2);

assign out_data_address1 = grp_tdf5_writeOutputs_unaligned_fu_88_out_data_address1;

assign out_data_ce1 = grp_tdf5_writeOutputs_unaligned_fu_88_out_data_ce1;

assign out_data_d1 = grp_tdf5_writeOutputs_unaligned_fu_88_out_data_d1;

assign out_data_we1 = grp_tdf5_writeOutputs_unaligned_fu_88_out_data_we1;

assign select_ln24_fu_126_p3 = ((or_ln24_fu_120_p2[0:0] == 1'b1) ? p_read : max_vals_5_0);

assign storeOutput7_read_read_fu_82_p2 = storeOutput7_dout;

endmodule //td_fused_top_tdf5_poolOutputs
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf5_readFilters40 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        filter_data_address0,
        filter_data_ce0,
        filter_data_q0,
        input_indices_23_dout,
        input_indices_23_empty_n,
        input_indices_23_read,
        weight_vecs_0_address0,
        weight_vecs_0_ce0,
        weight_vecs_0_we0,
        weight_vecs_0_d0
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state7 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [14:0] filter_data_address0;
output   filter_data_ce0;
input  [15:0] filter_data_q0;
input  [6:0] input_indices_23_dout;
input   input_indices_23_empty_n;
output   input_indices_23_read;
output  [7:0] weight_vecs_0_address0;
output   weight_vecs_0_ce0;
output   weight_vecs_0_we0;
output  [15:0] weight_vecs_0_d0;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg filter_data_ce0;
reg input_indices_23_read;
reg weight_vecs_0_ce0;
reg weight_vecs_0_we0;

reg    ap_done_reg;
  reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    input_indices_23_blk_n;
reg   [7:0] indvar_flatten13_reg_123;
reg   [1:0] ii_reg_134;
reg   [6:0] indvar_flatten_reg_145;
reg   [1:0] jj_reg_156;
reg   [4:0] kk_reg_167;
wire   [10:0] sext_ln47_fu_200_p1;
reg   [10:0] sext_ln47_reg_408;
wire   [7:0] add_ln47_3_fu_204_p2;
wire    ap_CS_fsm_pp0_stage0;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
wire    ap_block_state4_pp0_stage0_iter2;
wire    ap_block_state5_pp0_stage0_iter3;
wire    ap_block_state6_pp0_stage0_iter4;
wire    ap_block_pp0_stage0_11001;
wire   [0:0] icmp_ln47_fu_210_p2;
reg   [0:0] icmp_ln47_reg_418;
reg   [0:0] icmp_ln47_reg_418_pp0_iter1_reg;
reg   [0:0] icmp_ln47_reg_418_pp0_iter2_reg;
reg   [0:0] icmp_ln47_reg_418_pp0_iter3_reg;
wire   [0:0] icmp_ln48_fu_222_p2;
reg   [0:0] icmp_ln48_reg_422;
wire   [1:0] select_ln47_3_fu_228_p3;
reg   [1:0] select_ln47_3_reg_429;
wire   [6:0] select_ln48_6_fu_242_p3;
wire   [1:0] select_ln48_5_fu_329_p3;
reg   [1:0] select_ln48_5_reg_442;
reg    ap_enable_reg_pp0_iter1;
wire   [7:0] add_ln55_12_fu_392_p2;
reg   [7:0] add_ln55_12_reg_452;
reg   [7:0] add_ln55_12_reg_452_pp0_iter2_reg;
reg   [7:0] add_ln55_12_reg_452_pp0_iter3_reg;
wire   [4:0] add_ln49_fu_398_p2;
reg    ap_block_state1;
wire    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_flush_enable;
reg    ap_enable_reg_pp0_iter2;
reg    ap_condition_pp0_exit_iter1_state3;
reg    ap_enable_reg_pp0_iter3;
reg    ap_enable_reg_pp0_iter4;
reg   [1:0] ap_phi_mux_ii_phi_fu_138_p4;
wire    ap_block_pp0_stage0;
reg   [1:0] ap_phi_mux_jj_phi_fu_160_p4;
wire   [63:0] zext_ln55_28_fu_387_p1;
wire   [63:0] zext_ln55_29_fu_404_p1;
wire   [8:0] tmp_fu_182_p3;
wire   [9:0] zext_ln55_21_fu_190_p1;
wire   [9:0] zext_ln55_fu_178_p1;
wire   [9:0] sub_ln55_fu_194_p2;
wire   [1:0] add_ln47_fu_216_p2;
wire   [6:0] add_ln48_3_fu_236_p2;
wire   [10:0] zext_ln55_23_fu_260_p1;
wire   [10:0] add_ln55_fu_263_p2;
wire   [10:0] shl_ln55_fu_268_p2;
wire   [3:0] tmp_s_fu_280_p3;
wire   [3:0] zext_ln55_22_fu_257_p1;
wire   [0:0] icmp_ln49_fu_298_p2;
wire   [0:0] xor_ln47_fu_293_p2;
wire   [1:0] select_ln47_fu_250_p3;
wire   [0:0] and_ln47_fu_304_p2;
wire   [0:0] or_ln48_fu_316_p2;
wire   [1:0] add_ln48_fu_310_p2;
wire   [10:0] sub_ln55_5_fu_274_p2;
wire   [10:0] zext_ln55_25_fu_341_p1;
wire   [10:0] add_ln55_9_fu_345_p2;
wire   [3:0] sub_ln55_6_fu_287_p2;
wire   [3:0] zext_ln55_24_fu_337_p1;
wire   [3:0] add_ln55_10_fu_359_p2;
wire   [4:0] select_ln48_fu_321_p3;
wire   [14:0] tmp_74_cast_fu_351_p3;
wire   [14:0] zext_ln55_27_fu_377_p1;
wire   [14:0] add_ln55_11_fu_381_p2;
wire   [7:0] tmp_76_cast_fu_365_p3;
wire   [7:0] zext_ln55_26_fu_373_p1;
wire    ap_CS_fsm_state7;
reg   [2:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
#0 ap_enable_reg_pp0_iter4 = 1'b0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state7)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if ((1'b1 == ap_condition_pp0_flush_enable)) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((~((ap_start == 1'b0) | (input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            if ((1'b1 == ap_condition_pp0_exit_iter1_state3)) begin
                ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter0;
            end else if ((1'b1 == 1'b1)) begin
                ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
            end
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter4 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
        end else if ((~((ap_start == 1'b0) | (input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter4 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln47_reg_418 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ii_reg_134 <= select_ln47_3_reg_429;
    end else if ((~((ap_start == 1'b0) | (input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ii_reg_134 <= 2'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_fu_210_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        indvar_flatten13_reg_123 <= add_ln47_3_fu_204_p2;
    end else if ((~((ap_start == 1'b0) | (input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indvar_flatten13_reg_123 <= 8'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_fu_210_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        indvar_flatten_reg_145 <= select_ln48_6_fu_242_p3;
    end else if ((~((ap_start == 1'b0) | (input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indvar_flatten_reg_145 <= 7'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_reg_418_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        jj_reg_156 <= select_ln48_5_reg_442;
    end else if ((~((ap_start == 1'b0) | (input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        jj_reg_156 <= 2'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln47_reg_418 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        kk_reg_167 <= add_ln49_fu_398_p2;
    end else if ((~((ap_start == 1'b0) | (input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        kk_reg_167 <= 5'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_reg_418 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        add_ln55_12_reg_452 <= add_ln55_12_fu_392_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        add_ln55_12_reg_452_pp0_iter2_reg <= add_ln55_12_reg_452;
        add_ln55_12_reg_452_pp0_iter3_reg <= add_ln55_12_reg_452_pp0_iter2_reg;
        icmp_ln47_reg_418_pp0_iter2_reg <= icmp_ln47_reg_418_pp0_iter1_reg;
        icmp_ln47_reg_418_pp0_iter3_reg <= icmp_ln47_reg_418_pp0_iter2_reg;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln47_reg_418 <= icmp_ln47_fu_210_p2;
        icmp_ln47_reg_418_pp0_iter1_reg <= icmp_ln47_reg_418;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_fu_210_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln48_reg_422 <= icmp_ln48_fu_222_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_fu_210_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        select_ln47_3_reg_429 <= select_ln47_3_fu_228_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln47_reg_418 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        select_ln48_5_reg_442 <= select_ln48_5_fu_329_p3;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state1)) begin
        sext_ln47_reg_408 <= sext_ln47_fu_200_p1;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_condition_pp0_exit_iter1_state3 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter1_state3 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln47_fu_210_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_condition_pp0_flush_enable = 1'b1;
    end else begin
        ap_condition_pp0_flush_enable = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state7)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln47_reg_418 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_phi_mux_ii_phi_fu_138_p4 = select_ln47_3_reg_429;
    end else begin
        ap_phi_mux_ii_phi_fu_138_p4 = ii_reg_134;
    end
end

always @ (*) begin
    if (((icmp_ln47_reg_418_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        ap_phi_mux_jj_phi_fu_160_p4 = select_ln48_5_reg_442;
    end else begin
        ap_phi_mux_jj_phi_fu_160_p4 = jj_reg_156;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state7)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter3 == 1'b1)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter4 == 1'b1)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1)))) begin
        filter_data_ce0 = 1'b1;
    end else begin
        filter_data_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        input_indices_23_blk_n = input_indices_23_empty_n;
    end else begin
        input_indices_23_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        input_indices_23_read = 1'b1;
    end else begin
        input_indices_23_read = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter4 == 1'b1))) begin
        weight_vecs_0_ce0 = 1'b1;
    end else begin
        weight_vecs_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln47_reg_418_pp0_iter3_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter4 == 1'b1))) begin
        weight_vecs_0_we0 = 1'b1;
    end else begin
        weight_vecs_0_we0 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_start == 1'b0) | (input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((~((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b0)) & ~((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter4 == 1'b1) & (ap_enable_reg_pp0_iter3 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if ((((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b0)) | ((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter4 == 1'b1) & (ap_enable_reg_pp0_iter3 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_state7;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state7 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln47_3_fu_204_p2 = (indvar_flatten13_reg_123 + 8'd1);

assign add_ln47_fu_216_p2 = (ap_phi_mux_ii_phi_fu_138_p4 + 2'd1);

assign add_ln48_3_fu_236_p2 = (indvar_flatten_reg_145 + 7'd1);

assign add_ln48_fu_310_p2 = (select_ln47_fu_250_p3 + 2'd1);

assign add_ln49_fu_398_p2 = (select_ln48_fu_321_p3 + 5'd1);

assign add_ln55_10_fu_359_p2 = (sub_ln55_6_fu_287_p2 + zext_ln55_24_fu_337_p1);

assign add_ln55_11_fu_381_p2 = (tmp_74_cast_fu_351_p3 + zext_ln55_27_fu_377_p1);

assign add_ln55_12_fu_392_p2 = (tmp_76_cast_fu_365_p3 + zext_ln55_26_fu_373_p1);

assign add_ln55_9_fu_345_p2 = (sub_ln55_5_fu_274_p2 + zext_ln55_25_fu_341_p1);

assign add_ln55_fu_263_p2 = ((sext_ln47_reg_408) + (zext_ln55_23_fu_260_p1));

assign and_ln47_fu_304_p2 = (xor_ln47_fu_293_p2 & icmp_ln49_fu_298_p2);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state7 = ap_CS_fsm[32'd2];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1));
end

assign ap_block_state2_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter4 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign filter_data_address0 = zext_ln55_28_fu_387_p1;

assign icmp_ln47_fu_210_p2 = ((indvar_flatten13_reg_123 == 8'd144) ? 1'b1 : 1'b0);

assign icmp_ln48_fu_222_p2 = ((indvar_flatten_reg_145 == 7'd48) ? 1'b1 : 1'b0);

assign icmp_ln49_fu_298_p2 = ((kk_reg_167 == 5'd16) ? 1'b1 : 1'b0);

assign or_ln48_fu_316_p2 = (icmp_ln48_reg_422 | and_ln47_fu_304_p2);

assign select_ln47_3_fu_228_p3 = ((icmp_ln48_fu_222_p2[0:0] == 1'b1) ? add_ln47_fu_216_p2 : ap_phi_mux_ii_phi_fu_138_p4);

assign select_ln47_fu_250_p3 = ((icmp_ln48_reg_422[0:0] == 1'b1) ? 2'd0 : ap_phi_mux_jj_phi_fu_160_p4);

assign select_ln48_5_fu_329_p3 = ((and_ln47_fu_304_p2[0:0] == 1'b1) ? add_ln48_fu_310_p2 : select_ln47_fu_250_p3);

assign select_ln48_6_fu_242_p3 = ((icmp_ln48_fu_222_p2[0:0] == 1'b1) ? 7'd1 : add_ln48_3_fu_236_p2);

assign select_ln48_fu_321_p3 = ((or_ln48_fu_316_p2[0:0] == 1'b1) ? 5'd0 : kk_reg_167);

assign sext_ln47_fu_200_p1 = (sub_ln55_fu_194_p2);

assign shl_ln55_fu_268_p2 = add_ln55_fu_263_p2 << 11'd2;

assign sub_ln55_5_fu_274_p2 = (shl_ln55_fu_268_p2 - add_ln55_fu_263_p2);

assign sub_ln55_6_fu_287_p2 = (tmp_s_fu_280_p3 - zext_ln55_22_fu_257_p1);

assign sub_ln55_fu_194_p2 = (zext_ln55_21_fu_190_p1 - zext_ln55_fu_178_p1);

assign tmp_74_cast_fu_351_p3 = {{add_ln55_9_fu_345_p2}, {4'd0}};

assign tmp_76_cast_fu_365_p3 = {{add_ln55_10_fu_359_p2}, {4'd0}};

assign tmp_fu_182_p3 = {{input_indices_23_dout}, {2'd0}};

assign tmp_s_fu_280_p3 = {{select_ln47_3_reg_429}, {2'd0}};

assign weight_vecs_0_address0 = zext_ln55_29_fu_404_p1;

assign weight_vecs_0_d0 = filter_data_q0;

assign xor_ln47_fu_293_p2 = (icmp_ln48_reg_422 ^ 1'd1);

assign zext_ln55_21_fu_190_p1 = tmp_fu_182_p3;

assign zext_ln55_22_fu_257_p1 = select_ln47_3_reg_429;

assign zext_ln55_23_fu_260_p1 = select_ln47_3_reg_429;

assign zext_ln55_24_fu_337_p1 = select_ln48_5_fu_329_p3;

assign zext_ln55_25_fu_341_p1 = select_ln48_5_fu_329_p3;

assign zext_ln55_26_fu_373_p1 = select_ln48_fu_321_p3;

assign zext_ln55_27_fu_377_p1 = select_ln48_fu_321_p3;

assign zext_ln55_28_fu_387_p1 = add_ln55_11_fu_381_p2;

assign zext_ln55_29_fu_404_p1 = add_ln55_12_reg_452_pp0_iter3_reg;

assign zext_ln55_fu_178_p1 = input_indices_23_dout;

endmodule //td_fused_top_tdf5_readFilters40
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf5_readInputs41 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        in_data_address0,
        in_data_ce0,
        in_data_q0,
        i_15,
        j_15,
        ifmap_vec_address0,
        ifmap_vec_ce0,
        ifmap_vec_we0,
        ifmap_vec_d0,
        ifmap_vec_address1,
        ifmap_vec_ce1,
        ifmap_vec_we1,
        ifmap_vec_d1
);

parameter    ap_ST_fsm_state1 = 4'd1;
parameter    ap_ST_fsm_pp0_stage0 = 4'd2;
parameter    ap_ST_fsm_pp0_stage1 = 4'd4;
parameter    ap_ST_fsm_state8 = 4'd8;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [13:0] in_data_address0;
output   in_data_ce0;
input  [63:0] in_data_q0;
input  [15:0] i_15;
input  [15:0] j_15;
output  [7:0] ifmap_vec_address0;
output   ifmap_vec_ce0;
output   ifmap_vec_we0;
output  [15:0] ifmap_vec_d0;
output  [7:0] ifmap_vec_address1;
output   ifmap_vec_ce1;
output   ifmap_vec_we1;
output  [15:0] ifmap_vec_d1;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg in_data_ce0;
reg[7:0] ifmap_vec_address0;
reg ifmap_vec_ce0;
reg ifmap_vec_we0;
reg[15:0] ifmap_vec_d0;
reg[7:0] ifmap_vec_address1;
reg ifmap_vec_ce1;
reg ifmap_vec_we1;
reg[15:0] ifmap_vec_d1;

reg    ap_done_reg;
  reg   [3:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg   [5:0] indvar_flatten47_reg_194;
reg   [1:0] ii_reg_206;
reg   [4:0] indvar_flatten_reg_218;
reg   [1:0] jj_reg_229;
reg   [4:0] kk_0_i_reg_241;
wire   [17:0] p_cast_i_fu_270_p1;
reg   [17:0] p_cast_i_reg_931;
wire   [11:0] trunc_ln22_fu_274_p1;
reg   [11:0] trunc_ln22_reg_937;
wire   [17:0] sext_ln22_fu_284_p1;
reg   [17:0] sext_ln22_reg_943;
wire   [5:0] p_cast_fu_288_p2;
reg   [5:0] p_cast_reg_949;
wire   [0:0] or_ln23_11_fu_308_p2;
reg   [0:0] or_ln23_11_reg_955;
wire   [11:0] p_mid137_fu_314_p2;
reg   [11:0] p_mid137_reg_960;
wire   [5:0] p_cast5_i_fu_333_p2;
reg   [5:0] p_cast5_i_reg_965;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state4_pp0_stage0_iter1;
wire    ap_block_state6_pp0_stage0_iter2;
wire    ap_block_pp0_stage0_11001;
wire   [0:0] is_padding_fu_373_p2;
reg   [0:0] is_padding_reg_971;
wire   [0:0] icmp_ln19_fu_379_p2;
reg   [0:0] icmp_ln19_reg_978;
reg   [0:0] icmp_ln19_reg_978_pp0_iter1_reg;
reg   [0:0] icmp_ln19_reg_978_pp0_iter2_reg;
wire   [1:0] add_ln19_fu_385_p2;
reg   [1:0] add_ln19_reg_982;
wire   [0:0] icmp_ln20_fu_391_p2;
reg   [0:0] icmp_ln20_reg_987;
wire   [1:0] select_ln19_fu_397_p3;
reg   [1:0] select_ln19_reg_999;
wire   [5:0] p_cast5_i_mid1_fu_418_p2;
reg   [5:0] p_cast5_i_mid1_reg_1004;
wire   [0:0] or_ln23_13_fu_437_p2;
reg   [0:0] or_ln23_13_reg_1010;
wire   [1:0] add_ln20_fu_442_p2;
reg   [1:0] add_ln20_reg_1017;
wire   [0:0] or_ln23_15_fu_477_p2;
reg   [0:0] or_ln23_15_reg_1023;
wire   [4:0] add_ln20_3_fu_483_p2;
reg   [4:0] add_ln20_3_reg_1030;
wire   [5:0] add_ln19_3_fu_489_p2;
reg   [5:0] add_ln19_3_reg_1035;
wire    ap_CS_fsm_pp0_stage1;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_state3_pp0_stage1_iter0;
wire    ap_block_state5_pp0_stage1_iter1;
wire    ap_block_state7_pp0_stage1_iter2;
wire    ap_block_pp0_stage1_11001;
wire   [1:0] select_ln19_13_fu_527_p3;
reg   [1:0] select_ln19_13_reg_1040;
wire   [4:0] select_ln20_fu_591_p3;
reg   [4:0] select_ln20_reg_1047;
wire   [1:0] select_ln20_11_fu_599_p3;
reg   [1:0] select_ln20_11_reg_1053;
wire   [0:0] select_ln20_12_fu_608_p3;
reg   [0:0] select_ln20_12_reg_1059;
reg   [0:0] select_ln20_12_reg_1059_pp0_iter1_reg;
wire   [3:0] empty_87_fu_704_p1;
reg   [3:0] empty_87_reg_1067;
reg   [3:0] empty_87_reg_1067_pp0_iter1_reg;
wire   [4:0] select_ln20_15_fu_731_p3;
reg   [4:0] select_ln20_15_reg_1079;
wire   [4:0] add_ln25_fu_737_p2;
reg   [4:0] add_ln25_reg_1084;
reg    ap_enable_reg_pp0_iter1;
wire   [5:0] add_ln33_fu_769_p2;
reg   [5:0] add_ln33_reg_1089;
wire   [7:0] add_ln33_3_fu_790_p2;
reg   [7:0] add_ln33_3_reg_1096;
wire   [15:0] select_ln33_14_fu_869_p3;
reg   [15:0] select_ln33_14_reg_1101;
wire   [15:0] select_ln33_15_fu_890_p3;
reg   [15:0] select_ln33_15_reg_1106;
reg    ap_block_state1;
wire    ap_block_pp0_stage1_subdone;
reg    ap_condition_pp0_exit_iter0_state3;
reg    ap_enable_reg_pp0_iter2;
reg   [5:0] ap_phi_mux_indvar_flatten47_phi_fu_198_p4;
wire    ap_block_pp0_stage0;
reg   [1:0] ap_phi_mux_ii_phi_fu_210_p4;
reg   [4:0] ap_phi_mux_indvar_flatten_phi_fu_222_p4;
reg   [1:0] ap_phi_mux_jj_phi_fu_233_p4;
reg   [4:0] ap_phi_mux_kk_0_i_phi_fu_245_p4;
wire    ap_block_pp0_stage1;
wire   [63:0] sext_ln32_fu_726_p1;
wire   [63:0] zext_ln33_13_fu_796_p1;
wire   [63:0] sext_ln33_fu_828_p1;
wire   [63:0] sext_ln33_5_fu_909_p1;
wire   [63:0] sext_ln33_6_fu_926_p1;
wire   [15:0] select_ln33_fu_808_p3;
wire   [15:0] select_ln33_13_fu_847_p3;
wire   [16:0] zext_ln19_fu_256_p1;
wire   [16:0] empty_82_fu_264_p2;
wire   [16:0] j_cast_i_fu_252_p1;
wire   [16:0] add_ln22_fu_278_p2;
wire   [5:0] empty_fu_260_p1;
wire   [0:0] tmp_fu_294_p3;
wire   [0:0] icmp_ln24_fu_302_p2;
wire   [17:0] ii_cast_i_fu_320_p1;
wire   [5:0] ii_cast_fu_324_p1;
wire   [17:0] empty_83_fu_328_p2;
wire   [17:0] zext_ln20_fu_344_p1;
wire   [17:0] add_ln22_3_fu_348_p2;
wire   [0:0] tmp_20_fu_353_p3;
wire   [0:0] icmp_ln24_3_fu_361_p2;
wire   [0:0] or_ln23_fu_367_p2;
wire   [0:0] empty_84_fu_338_p2;
wire   [17:0] ii_cast_i_mid1_fu_405_p1;
wire   [5:0] ii_cast_mid1_fu_409_p1;
wire   [17:0] p_mid111_fu_413_p2;
wire   [0:0] p_mid113_fu_423_p2;
wire   [17:0] zext_ln20_3_fu_448_p1;
wire   [17:0] add_ln22_4_fu_452_p2;
wire   [0:0] tmp_21_fu_457_p3;
wire   [0:0] icmp_ln24_4_fu_465_p2;
wire   [0:0] or_ln23_14_fu_471_p2;
wire   [0:0] select_ln19_15_fu_429_p3;
wire   [2:0] zext_ln22_fu_495_p1;
wire   [2:0] tmp2_fu_505_p2;
wire   [11:0] tmp2_cast_fu_511_p1;
wire   [11:0] empty_85_fu_515_p2;
wire   [5:0] row_coord_int_mid131_fu_543_p3;
wire   [5:0] row_coord_int_fu_499_p3;
wire   [11:0] col_coord_int_mid139_fu_549_p3;
wire   [11:0] col_coord_int_fu_520_p3;
wire   [0:0] icmp_ln25_fu_574_p2;
wire   [0:0] xor_ln19_fu_569_p2;
wire   [0:0] and_ln19_fu_580_p2;
wire   [0:0] or_ln20_fu_586_p2;
wire   [0:0] select_ln19_16_fu_538_p3;
wire   [5:0] select_ln19_14_fu_533_p3;
wire   [2:0] zext_ln22_3_fu_605_p1;
wire   [2:0] tmp2_mid1_fu_622_p2;
wire   [11:0] tmp2_cast_mid1_fu_628_p1;
wire   [11:0] p_mid1_fu_632_p2;
wire   [5:0] row_coord_int_mid1_fu_615_p3;
wire   [5:0] select_ln19_17_fu_555_p3;
wire   [5:0] select_ln20_13_fu_644_p3;
wire   [11:0] tmp_4_fu_652_p3;
wire   [8:0] tmp_5_fu_664_p3;
wire   [12:0] zext_ln32_fu_660_p1;
wire   [12:0] zext_ln32_16_fu_672_p1;
wire   [12:0] sub_ln32_fu_676_p2;
wire   [11:0] col_coord_int_mid1_fu_637_p3;
wire   [11:0] select_ln19_18_fu_562_p3;
wire   [11:0] select_ln20_14_fu_686_p3;
wire   [13:0] sext_ln20_fu_682_p1;
wire   [13:0] zext_ln32_17_fu_694_p1;
wire   [13:0] add_ln32_fu_698_p2;
wire   [1:0] lshr_ln_fu_708_p4;
wire   [15:0] tmp_22_fu_718_p3;
wire   [3:0] tmp_s_fu_745_p3;
wire   [4:0] zext_ln33_10_fu_752_p1;
wire   [4:0] zext_ln33_fu_742_p1;
wire   [4:0] sub_ln33_fu_756_p2;
wire   [5:0] sub_ln33_cast_fu_762_p1;
wire   [5:0] zext_ln33_11_fu_766_p1;
wire   [3:0] trunc_ln33_fu_775_p1;
wire   [7:0] tmp_63_cast_fu_779_p3;
wire   [7:0] zext_ln33_12_fu_787_p1;
wire   [15:0] trunc_ln32_fu_800_p1;
wire   [15:0] bitcast_ln32_fu_804_p1;
wire   [3:0] or_ln25_fu_816_p2;
wire   [9:0] tmp_23_fu_821_p3;
wire   [15:0] tmp_39_i_fu_833_p4;
wire   [15:0] bitcast_ln32_13_fu_843_p1;
wire   [15:0] tmp_40_i_fu_855_p4;
wire   [15:0] bitcast_ln32_14_fu_865_p1;
wire   [15:0] tmp_41_i_fu_876_p4;
wire   [15:0] bitcast_ln32_15_fu_886_p1;
wire   [3:0] or_ln25_9_fu_897_p2;
wire   [9:0] tmp_24_fu_902_p3;
wire   [3:0] or_ln25_10_fu_914_p2;
wire   [9:0] tmp_25_fu_919_p3;
wire    ap_CS_fsm_state8;
reg   [3:0] ap_NS_fsm;
wire    ap_block_pp0_stage0_subdone;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 4'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_condition_pp0_exit_iter0_state3) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            if ((1'b1 == ap_condition_pp0_exit_iter0_state3)) begin
                ap_enable_reg_pp0_iter1 <= (1'b1 ^ ap_condition_pp0_exit_iter0_state3);
            end else if ((1'b1 == 1'b1)) begin
                ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
            end
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter2 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln19_reg_978 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ii_reg_206 <= select_ln19_13_reg_1040;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ii_reg_206 <= 2'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln19_reg_978 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        indvar_flatten47_reg_194 <= add_ln19_3_reg_1035;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indvar_flatten47_reg_194 <= 6'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln19_reg_978 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        indvar_flatten_reg_218 <= select_ln20_15_reg_1079;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indvar_flatten_reg_218 <= 5'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln19_reg_978 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        jj_reg_229 <= select_ln20_11_reg_1053;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        jj_reg_229 <= 2'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln19_reg_978_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        kk_0_i_reg_241 <= add_ln25_reg_1084;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        kk_0_i_reg_241 <= 5'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
        add_ln19_3_reg_1035 <= add_ln19_3_fu_489_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln19_fu_379_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        add_ln19_reg_982 <= add_ln19_fu_385_p2;
        add_ln20_3_reg_1030 <= add_ln20_3_fu_483_p2;
        add_ln20_reg_1017 <= add_ln20_fu_442_p2;
        icmp_ln20_reg_987 <= icmp_ln20_fu_391_p2;
        or_ln23_13_reg_1010 <= or_ln23_13_fu_437_p2;
        or_ln23_15_reg_1023 <= or_ln23_15_fu_477_p2;
        p_cast5_i_mid1_reg_1004 <= p_cast5_i_mid1_fu_418_p2;
        select_ln19_reg_999 <= select_ln19_fu_397_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln19_reg_978 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        add_ln25_reg_1084 <= add_ln25_fu_737_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln19_reg_978_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
        add_ln33_3_reg_1096 <= add_ln33_3_fu_790_p2;
        add_ln33_reg_1089 <= add_ln33_fu_769_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln19_reg_978 == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
        empty_87_reg_1067 <= empty_87_fu_704_p1;
        select_ln20_12_reg_1059 <= select_ln20_12_fu_608_p3;
        select_ln20_reg_1047 <= select_ln20_fu_591_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
        empty_87_reg_1067_pp0_iter1_reg <= empty_87_reg_1067;
        select_ln20_12_reg_1059_pp0_iter1_reg <= select_ln20_12_reg_1059;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln19_reg_978 <= icmp_ln19_fu_379_p2;
        icmp_ln19_reg_978_pp0_iter1_reg <= icmp_ln19_reg_978;
        icmp_ln19_reg_978_pp0_iter2_reg <= icmp_ln19_reg_978_pp0_iter1_reg;
        is_padding_reg_971 <= is_padding_fu_373_p2;
        p_cast5_i_reg_965 <= p_cast5_i_fu_333_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state1)) begin
        or_ln23_11_reg_955 <= or_ln23_11_fu_308_p2;
        p_cast_i_reg_931 <= p_cast_i_fu_270_p1;
        p_cast_reg_949 <= p_cast_fu_288_p2;
        p_mid137_reg_960 <= p_mid137_fu_314_p2;
        sext_ln22_reg_943 <= sext_ln22_fu_284_p1;
        trunc_ln22_reg_937 <= trunc_ln22_fu_274_p1;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln19_reg_978 == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
        select_ln19_13_reg_1040 <= select_ln19_13_fu_527_p3;
        select_ln20_11_reg_1053 <= select_ln20_11_fu_599_p3;
        select_ln20_15_reg_1079 <= select_ln20_15_fu_731_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln19_reg_978_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        select_ln33_14_reg_1101 <= select_ln33_14_fu_869_p3;
        select_ln33_15_reg_1106 <= select_ln33_15_fu_890_p3;
    end
end

always @ (*) begin
    if ((icmp_ln19_reg_978 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state3 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state3 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state8)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln19_reg_978 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_ii_phi_fu_210_p4 = select_ln19_13_reg_1040;
    end else begin
        ap_phi_mux_ii_phi_fu_210_p4 = ii_reg_206;
    end
end

always @ (*) begin
    if (((icmp_ln19_reg_978 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_indvar_flatten47_phi_fu_198_p4 = add_ln19_3_reg_1035;
    end else begin
        ap_phi_mux_indvar_flatten47_phi_fu_198_p4 = indvar_flatten47_reg_194;
    end
end

always @ (*) begin
    if (((icmp_ln19_reg_978 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_indvar_flatten_phi_fu_222_p4 = select_ln20_15_reg_1079;
    end else begin
        ap_phi_mux_indvar_flatten_phi_fu_222_p4 = indvar_flatten_reg_218;
    end
end

always @ (*) begin
    if (((icmp_ln19_reg_978 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_jj_phi_fu_233_p4 = select_ln20_11_reg_1053;
    end else begin
        ap_phi_mux_jj_phi_fu_233_p4 = jj_reg_229;
    end
end

always @ (*) begin
    if (((icmp_ln19_reg_978_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_kk_0_i_phi_fu_245_p4 = add_ln25_reg_1084;
    end else begin
        ap_phi_mux_kk_0_i_phi_fu_245_p4 = kk_0_i_reg_241;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state8)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((ap_enable_reg_pp0_iter2 == 1'b1)) begin
        if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            ifmap_vec_address0 = sext_ln33_6_fu_926_p1;
        end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ifmap_vec_address0 = sext_ln33_fu_828_p1;
        end else begin
            ifmap_vec_address0 = 'bx;
        end
    end else begin
        ifmap_vec_address0 = 'bx;
    end
end

always @ (*) begin
    if ((ap_enable_reg_pp0_iter2 == 1'b1)) begin
        if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            ifmap_vec_address1 = sext_ln33_5_fu_909_p1;
        end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ifmap_vec_address1 = zext_ln33_13_fu_796_p1;
        end else begin
            ifmap_vec_address1 = 'bx;
        end
    end else begin
        ifmap_vec_address1 = 'bx;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1)) | ((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter2 == 1'b1)))) begin
        ifmap_vec_ce0 = 1'b1;
    end else begin
        ifmap_vec_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1)) | ((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter2 == 1'b1)))) begin
        ifmap_vec_ce1 = 1'b1;
    end else begin
        ifmap_vec_ce1 = 1'b0;
    end
end

always @ (*) begin
    if ((ap_enable_reg_pp0_iter2 == 1'b1)) begin
        if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            ifmap_vec_d0 = select_ln33_15_reg_1106;
        end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ifmap_vec_d0 = select_ln33_13_fu_847_p3;
        end else begin
            ifmap_vec_d0 = 'bx;
        end
    end else begin
        ifmap_vec_d0 = 'bx;
    end
end

always @ (*) begin
    if ((ap_enable_reg_pp0_iter2 == 1'b1)) begin
        if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            ifmap_vec_d1 = select_ln33_14_reg_1101;
        end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ifmap_vec_d1 = select_ln33_fu_808_p3;
        end else begin
            ifmap_vec_d1 = 'bx;
        end
    end else begin
        ifmap_vec_d1 = 'bx;
    end
end

always @ (*) begin
    if ((((icmp_ln19_reg_978_pp0_iter2_reg == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter2 == 1'b1)) | ((icmp_ln19_reg_978_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1)))) begin
        ifmap_vec_we0 = 1'b1;
    end else begin
        ifmap_vec_we0 = 1'b0;
    end
end

always @ (*) begin
    if ((((icmp_ln19_reg_978_pp0_iter2_reg == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter2 == 1'b1)) | ((icmp_ln19_reg_978_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1)))) begin
        ifmap_vec_we1 = 1'b1;
    end else begin
        ifmap_vec_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1)) | ((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1)) | ((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1)) | ((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1)))) begin
        in_data_ce0 = 1'b1;
    end else begin
        in_data_ce0 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_pp0_stage1 : begin
            if ((~((icmp_ln19_reg_978 == 1'd1) & (1'b0 == ap_block_pp0_stage1_subdone) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1)) & ~((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter2 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0)) & (1'b0 == ap_block_pp0_stage1_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if ((((icmp_ln19_reg_978 == 1'd1) & (1'b0 == ap_block_pp0_stage1_subdone) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1)) | ((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter2 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_state8;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end
        end
        ap_ST_fsm_state8 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln19_3_fu_489_p2 = (indvar_flatten47_reg_194 + 6'd1);

assign add_ln19_fu_385_p2 = (ap_phi_mux_ii_phi_fu_210_p4 + 2'd1);

assign add_ln20_3_fu_483_p2 = (ap_phi_mux_indvar_flatten_phi_fu_222_p4 + 5'd1);

assign add_ln20_fu_442_p2 = (select_ln19_fu_397_p3 + 2'd1);

assign add_ln22_3_fu_348_p2 = ((sext_ln22_reg_943) + (zext_ln20_fu_344_p1));

assign add_ln22_4_fu_452_p2 = ((sext_ln22_reg_943) + (zext_ln20_3_fu_448_p1));

assign add_ln22_fu_278_p2 = ((j_cast_i_fu_252_p1) + (17'd131071));

assign add_ln25_fu_737_p2 = (select_ln20_reg_1047 + 5'd4);

assign add_ln32_fu_698_p2 = ((sext_ln20_fu_682_p1) + (zext_ln32_17_fu_694_p1));

assign add_ln33_3_fu_790_p2 = (tmp_63_cast_fu_779_p3 + zext_ln33_12_fu_787_p1);

assign add_ln33_fu_769_p2 = ((sub_ln33_cast_fu_762_p1) + (zext_ln33_11_fu_766_p1));

assign and_ln19_fu_580_p2 = (xor_ln19_fu_569_p2 & icmp_ln25_fu_574_p2);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_pp0_stage1 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state8 = ap_CS_fsm[32'd3];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (ap_done_reg == 1'b1));
end

assign ap_block_state2_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage1_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage1_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage1_iter2 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign bitcast_ln32_13_fu_843_p1 = tmp_39_i_fu_833_p4;

assign bitcast_ln32_14_fu_865_p1 = tmp_40_i_fu_855_p4;

assign bitcast_ln32_15_fu_886_p1 = tmp_41_i_fu_876_p4;

assign bitcast_ln32_fu_804_p1 = trunc_ln32_fu_800_p1;

assign col_coord_int_fu_520_p3 = ((is_padding_reg_971[0:0] == 1'b1) ? 12'd0 : empty_85_fu_515_p2);

assign col_coord_int_mid139_fu_549_p3 = ((or_ln23_13_reg_1010[0:0] == 1'b1) ? 12'd0 : p_mid137_reg_960);

assign col_coord_int_mid1_fu_637_p3 = ((or_ln23_15_reg_1023[0:0] == 1'b1) ? 12'd0 : p_mid1_fu_632_p2);

assign empty_82_fu_264_p2 = ((zext_ln19_fu_256_p1) + (17'd131071));

assign empty_83_fu_328_p2 = ((p_cast_i_reg_931) + (ii_cast_i_fu_320_p1));

assign empty_84_fu_338_p2 = ((empty_83_fu_328_p2 > 18'd55) ? 1'b1 : 1'b0);

assign empty_85_fu_515_p2 = ((tmp2_cast_fu_511_p1) + (trunc_ln22_reg_937));

assign empty_87_fu_704_p1 = select_ln20_fu_591_p3[3:0];

assign empty_fu_260_p1 = i_15[5:0];

assign icmp_ln19_fu_379_p2 = ((ap_phi_mux_indvar_flatten47_phi_fu_198_p4 == 6'd36) ? 1'b1 : 1'b0);

assign icmp_ln20_fu_391_p2 = ((ap_phi_mux_indvar_flatten_phi_fu_222_p4 == 5'd12) ? 1'b1 : 1'b0);

assign icmp_ln24_3_fu_361_p2 = (((add_ln22_3_fu_348_p2) > (18'd55)) ? 1'b1 : 1'b0);

assign icmp_ln24_4_fu_465_p2 = (((add_ln22_4_fu_452_p2) > (18'd55)) ? 1'b1 : 1'b0);

assign icmp_ln24_fu_302_p2 = (((add_ln22_fu_278_p2) > (17'd55)) ? 1'b1 : 1'b0);

assign icmp_ln25_fu_574_p2 = ((ap_phi_mux_kk_0_i_phi_fu_245_p4 == 5'd16) ? 1'b1 : 1'b0);

assign ii_cast_fu_324_p1 = ap_phi_mux_ii_phi_fu_210_p4;

assign ii_cast_i_fu_320_p1 = ap_phi_mux_ii_phi_fu_210_p4;

assign ii_cast_i_mid1_fu_405_p1 = add_ln19_fu_385_p2;

assign ii_cast_mid1_fu_409_p1 = add_ln19_fu_385_p2;

assign in_data_address0 = sext_ln32_fu_726_p1;

assign is_padding_fu_373_p2 = (or_ln23_fu_367_p2 | empty_84_fu_338_p2);

assign j_cast_i_fu_252_p1 = j_15;

assign lshr_ln_fu_708_p4 = {{select_ln20_fu_591_p3[3:2]}};

assign or_ln20_fu_586_p2 = (icmp_ln20_reg_987 | and_ln19_fu_580_p2);

assign or_ln23_11_fu_308_p2 = (tmp_fu_294_p3 | icmp_ln24_fu_302_p2);

assign or_ln23_13_fu_437_p2 = (p_mid113_fu_423_p2 | or_ln23_11_reg_955);

assign or_ln23_14_fu_471_p2 = (tmp_21_fu_457_p3 | icmp_ln24_4_fu_465_p2);

assign or_ln23_15_fu_477_p2 = (select_ln19_15_fu_429_p3 | or_ln23_14_fu_471_p2);

assign or_ln23_fu_367_p2 = (tmp_20_fu_353_p3 | icmp_ln24_3_fu_361_p2);

assign or_ln25_10_fu_914_p2 = (empty_87_reg_1067_pp0_iter1_reg | 4'd3);

assign or_ln25_9_fu_897_p2 = (empty_87_reg_1067_pp0_iter1_reg | 4'd2);

assign or_ln25_fu_816_p2 = (empty_87_reg_1067_pp0_iter1_reg | 4'd1);

assign p_cast5_i_fu_333_p2 = (p_cast_reg_949 + ii_cast_fu_324_p1);

assign p_cast5_i_mid1_fu_418_p2 = (p_cast_reg_949 + ii_cast_mid1_fu_409_p1);

assign p_cast_fu_288_p2 = ((empty_fu_260_p1) + (6'd63));

assign p_cast_i_fu_270_p1 = (empty_82_fu_264_p2);

assign p_mid111_fu_413_p2 = ((p_cast_i_reg_931) + (ii_cast_i_mid1_fu_405_p1));

assign p_mid113_fu_423_p2 = ((p_mid111_fu_413_p2 > 18'd55) ? 1'b1 : 1'b0);

assign p_mid137_fu_314_p2 = ((trunc_ln22_fu_274_p1) + (12'd4095));

assign p_mid1_fu_632_p2 = ((tmp2_cast_mid1_fu_628_p1) + (trunc_ln22_reg_937));

assign row_coord_int_fu_499_p3 = ((is_padding_reg_971[0:0] == 1'b1) ? 6'd0 : p_cast5_i_reg_965);

assign row_coord_int_mid131_fu_543_p3 = ((or_ln23_13_reg_1010[0:0] == 1'b1) ? 6'd0 : p_cast5_i_mid1_reg_1004);

assign row_coord_int_mid1_fu_615_p3 = ((or_ln23_15_reg_1023[0:0] == 1'b1) ? 6'd0 : select_ln19_14_fu_533_p3);

assign select_ln19_13_fu_527_p3 = ((icmp_ln20_reg_987[0:0] == 1'b1) ? add_ln19_reg_982 : ii_reg_206);

assign select_ln19_14_fu_533_p3 = ((icmp_ln20_reg_987[0:0] == 1'b1) ? p_cast5_i_mid1_reg_1004 : p_cast5_i_reg_965);

assign select_ln19_15_fu_429_p3 = ((icmp_ln20_fu_391_p2[0:0] == 1'b1) ? p_mid113_fu_423_p2 : empty_84_fu_338_p2);

assign select_ln19_16_fu_538_p3 = ((icmp_ln20_reg_987[0:0] == 1'b1) ? or_ln23_13_reg_1010 : is_padding_reg_971);

assign select_ln19_17_fu_555_p3 = ((icmp_ln20_reg_987[0:0] == 1'b1) ? row_coord_int_mid131_fu_543_p3 : row_coord_int_fu_499_p3);

assign select_ln19_18_fu_562_p3 = ((icmp_ln20_reg_987[0:0] == 1'b1) ? col_coord_int_mid139_fu_549_p3 : col_coord_int_fu_520_p3);

assign select_ln19_fu_397_p3 = ((icmp_ln20_fu_391_p2[0:0] == 1'b1) ? 2'd0 : ap_phi_mux_jj_phi_fu_233_p4);

assign select_ln20_11_fu_599_p3 = ((and_ln19_fu_580_p2[0:0] == 1'b1) ? add_ln20_reg_1017 : select_ln19_reg_999);

assign select_ln20_12_fu_608_p3 = ((and_ln19_fu_580_p2[0:0] == 1'b1) ? or_ln23_15_reg_1023 : select_ln19_16_fu_538_p3);

assign select_ln20_13_fu_644_p3 = ((and_ln19_fu_580_p2[0:0] == 1'b1) ? row_coord_int_mid1_fu_615_p3 : select_ln19_17_fu_555_p3);

assign select_ln20_14_fu_686_p3 = ((and_ln19_fu_580_p2[0:0] == 1'b1) ? col_coord_int_mid1_fu_637_p3 : select_ln19_18_fu_562_p3);

assign select_ln20_15_fu_731_p3 = ((icmp_ln20_reg_987[0:0] == 1'b1) ? 5'd1 : add_ln20_3_reg_1030);

assign select_ln20_fu_591_p3 = ((or_ln20_fu_586_p2[0:0] == 1'b1) ? 5'd0 : ap_phi_mux_kk_0_i_phi_fu_245_p4);

assign select_ln33_13_fu_847_p3 = ((select_ln20_12_reg_1059_pp0_iter1_reg[0:0] == 1'b1) ? 16'd0 : bitcast_ln32_13_fu_843_p1);

assign select_ln33_14_fu_869_p3 = ((select_ln20_12_reg_1059_pp0_iter1_reg[0:0] == 1'b1) ? 16'd0 : bitcast_ln32_14_fu_865_p1);

assign select_ln33_15_fu_890_p3 = ((select_ln20_12_reg_1059_pp0_iter1_reg[0:0] == 1'b1) ? 16'd0 : bitcast_ln32_15_fu_886_p1);

assign select_ln33_fu_808_p3 = ((select_ln20_12_reg_1059_pp0_iter1_reg[0:0] == 1'b1) ? 16'd0 : bitcast_ln32_fu_804_p1);

assign sext_ln20_fu_682_p1 = (sub_ln32_fu_676_p2);

assign sext_ln22_fu_284_p1 = add_ln22_fu_278_p2;

assign sext_ln32_fu_726_p1 = (tmp_22_fu_718_p3);

assign sext_ln33_5_fu_909_p1 = (tmp_24_fu_902_p3);

assign sext_ln33_6_fu_926_p1 = (tmp_25_fu_919_p3);

assign sext_ln33_fu_828_p1 = (tmp_23_fu_821_p3);

assign sub_ln32_fu_676_p2 = (zext_ln32_fu_660_p1 - zext_ln32_16_fu_672_p1);

assign sub_ln33_cast_fu_762_p1 = (sub_ln33_fu_756_p2);

assign sub_ln33_fu_756_p2 = (zext_ln33_10_fu_752_p1 - zext_ln33_fu_742_p1);

assign tmp2_cast_fu_511_p1 = (tmp2_fu_505_p2);

assign tmp2_cast_mid1_fu_628_p1 = (tmp2_mid1_fu_622_p2);

assign tmp2_fu_505_p2 = ((zext_ln22_fu_495_p1) + (3'd7));

assign tmp2_mid1_fu_622_p2 = ((zext_ln22_3_fu_605_p1) + (3'd7));

assign tmp_20_fu_353_p3 = add_ln22_3_fu_348_p2[32'd17];

assign tmp_21_fu_457_p3 = add_ln22_4_fu_452_p2[32'd17];

assign tmp_22_fu_718_p3 = {{add_ln32_fu_698_p2}, {lshr_ln_fu_708_p4}};

assign tmp_23_fu_821_p3 = {{add_ln33_reg_1089}, {or_ln25_fu_816_p2}};

assign tmp_24_fu_902_p3 = {{add_ln33_reg_1089}, {or_ln25_9_fu_897_p2}};

assign tmp_25_fu_919_p3 = {{add_ln33_reg_1089}, {or_ln25_10_fu_914_p2}};

assign tmp_39_i_fu_833_p4 = {{in_data_q0[31:16]}};

assign tmp_40_i_fu_855_p4 = {{in_data_q0[47:32]}};

assign tmp_41_i_fu_876_p4 = {{in_data_q0[63:48]}};

assign tmp_4_fu_652_p3 = {{select_ln20_13_fu_644_p3}, {6'd0}};

assign tmp_5_fu_664_p3 = {{select_ln20_13_fu_644_p3}, {3'd0}};

assign tmp_63_cast_fu_779_p3 = {{trunc_ln33_fu_775_p1}, {4'd0}};

assign tmp_fu_294_p3 = add_ln22_fu_278_p2[32'd16];

assign tmp_s_fu_745_p3 = {{select_ln19_13_reg_1040}, {2'd0}};

assign trunc_ln22_fu_274_p1 = j_15[11:0];

assign trunc_ln32_fu_800_p1 = in_data_q0[15:0];

assign trunc_ln33_fu_775_p1 = add_ln33_fu_769_p2[3:0];

assign xor_ln19_fu_569_p2 = (icmp_ln20_reg_987 ^ 1'd1);

assign zext_ln19_fu_256_p1 = i_15;

assign zext_ln20_3_fu_448_p1 = add_ln20_fu_442_p2;

assign zext_ln20_fu_344_p1 = ap_phi_mux_jj_phi_fu_233_p4;

assign zext_ln22_3_fu_605_p1 = add_ln20_reg_1017;

assign zext_ln22_fu_495_p1 = jj_reg_229;

assign zext_ln32_16_fu_672_p1 = tmp_5_fu_664_p3;

assign zext_ln32_17_fu_694_p1 = select_ln20_14_fu_686_p3;

assign zext_ln32_fu_660_p1 = tmp_4_fu_652_p3;

assign zext_ln33_10_fu_752_p1 = tmp_s_fu_745_p3;

assign zext_ln33_11_fu_766_p1 = select_ln20_11_reg_1053;

assign zext_ln33_12_fu_787_p1 = select_ln20_reg_1047;

assign zext_ln33_13_fu_796_p1 = add_ln33_3_reg_1096;

assign zext_ln33_fu_742_p1 = select_ln19_13_reg_1040;

endmodule //td_fused_top_tdf5_readInputs41
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf5_writeOutputs_unaligned (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        i,
        j,
        out_data_address1,
        out_data_ce1,
        out_data_we1,
        out_data_d1,
        max_vals_5_0
);

parameter    ap_ST_fsm_state1 = 2'd1;
parameter    ap_ST_fsm_state2 = 2'd2;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
input  [4:0] i;
input  [9:0] j;
output  [14:0] out_data_address1;
output   out_data_ce1;
output   out_data_we1;
output  [63:0] out_data_d1;
input  [15:0] max_vals_5_0;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg out_data_ce1;
reg out_data_we1;

  reg   [1:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg   [15:0] outputCount_5;
reg   [15:0] outputChanIdx_5;
reg   [15:0] outputRow_11_0;
reg   [15:0] outputRow_11_1;
reg   [15:0] outputRow_11_2;
reg   [15:0] outputRow_11_3;
wire   [15:0] add_ln87_fu_173_p2;
wire   [0:0] icmp_ln88_fu_179_p2;
reg   [0:0] icmp_ln88_reg_293;
reg   [15:0] ap_phi_mux_empty_phi_fu_90_p4;
reg   [15:0] empty_reg_87;
wire    ap_CS_fsm_state2;
wire   [63:0] zext_ln94_8_fu_207_p1;
wire   [15:0] select_ln97_fu_265_p3;
wire   [1:0] trunc_ln86_fu_145_p1;
reg   [15:0] ap_sig_allocacmp_outputRow_11_0_load;
reg   [15:0] ap_sig_allocacmp_outputRow_11_1_load;
reg   [15:0] ap_sig_allocacmp_outputRow_11_2_load;
reg   [15:0] ap_sig_allocacmp_outputRow_11_3_load;
wire   [6:0] tmp_s_fu_105_p3;
wire   [9:0] tmp_fu_97_p3;
wire   [9:0] zext_ln94_fu_113_p1;
wire   [9:0] sub_ln94_fu_117_p2;
wire   [9:0] add_ln94_fu_123_p2;
wire   [6:0] trunc_ln94_fu_193_p1;
wire   [14:0] tmp_60_cast_fu_129_p3;
wire   [14:0] zext_ln94_7_fu_197_p1;
wire   [14:0] add_ln94_4_fu_201_p2;
wire   [15:0] bitcast_ln94_12_fu_236_p1;
wire   [15:0] bitcast_ln94_11_fu_228_p1;
wire   [15:0] bitcast_ln94_10_fu_220_p1;
wire   [15:0] bitcast_ln94_fu_212_p1;
wire   [15:0] add_ln96_fu_253_p2;
wire   [0:0] icmp_ln97_fu_259_p2;
reg   [1:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_CS_fsm = 2'd1;
#0 outputCount_5 = 16'd0;
#0 outputChanIdx_5 = 16'd0;
#0 outputRow_11_0 = 16'd0;
#0 outputRow_11_1 = 16'd0;
#0 outputRow_11_2 = 16'd0;
#0 outputRow_11_3 = 16'd0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln88_reg_293 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        empty_reg_87 <= 16'd0;
    end else if (((ap_start == 1'b1) & (icmp_ln88_fu_179_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state1))) begin
        empty_reg_87 <= add_ln87_fu_173_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state1)) begin
        icmp_ln88_reg_293 <= icmp_ln88_fu_179_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_start == 1'b1) & (icmp_ln88_fu_179_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1))) begin
        outputChanIdx_5 <= select_ln97_fu_265_p3;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        outputCount_5 <= ap_phi_mux_empty_phi_fu_90_p4;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_start == 1'b1) & (trunc_ln86_fu_145_p1 == 2'd0) & (1'b1 == ap_CS_fsm_state1))) begin
        outputRow_11_0 <= max_vals_5_0;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_start == 1'b1) & (trunc_ln86_fu_145_p1 == 2'd1) & (1'b1 == ap_CS_fsm_state1))) begin
        outputRow_11_1 <= max_vals_5_0;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_start == 1'b1) & (trunc_ln86_fu_145_p1 == 2'd2) & (1'b1 == ap_CS_fsm_state1))) begin
        outputRow_11_2 <= max_vals_5_0;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_start == 1'b1) & (trunc_ln86_fu_145_p1 == 2'd3) & (1'b1 == ap_CS_fsm_state1))) begin
        outputRow_11_3 <= max_vals_5_0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state2) | ((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1)))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = 1'b0;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln88_reg_293 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        ap_phi_mux_empty_phi_fu_90_p4 = 16'd0;
    end else begin
        ap_phi_mux_empty_phi_fu_90_p4 = empty_reg_87;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((trunc_ln86_fu_145_p1 == 2'd0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_sig_allocacmp_outputRow_11_0_load = max_vals_5_0;
    end else begin
        ap_sig_allocacmp_outputRow_11_0_load = outputRow_11_0;
    end
end

always @ (*) begin
    if (((trunc_ln86_fu_145_p1 == 2'd1) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_sig_allocacmp_outputRow_11_1_load = max_vals_5_0;
    end else begin
        ap_sig_allocacmp_outputRow_11_1_load = outputRow_11_1;
    end
end

always @ (*) begin
    if (((trunc_ln86_fu_145_p1 == 2'd2) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_sig_allocacmp_outputRow_11_2_load = max_vals_5_0;
    end else begin
        ap_sig_allocacmp_outputRow_11_2_load = outputRow_11_2;
    end
end

always @ (*) begin
    if (((trunc_ln86_fu_145_p1 == 2'd3) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_sig_allocacmp_outputRow_11_3_load = max_vals_5_0;
    end else begin
        ap_sig_allocacmp_outputRow_11_3_load = outputRow_11_3;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state2) | ((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)))) begin
        out_data_ce1 = 1'b1;
    end else begin
        out_data_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_start == 1'b1) & (icmp_ln88_fu_179_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1))) begin
        out_data_we1 = 1'b1;
    end else begin
        out_data_we1 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_state2 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln87_fu_173_p2 = (outputCount_5 + 16'd1);

assign add_ln94_4_fu_201_p2 = (tmp_60_cast_fu_129_p3 + zext_ln94_7_fu_197_p1);

assign add_ln94_fu_123_p2 = (sub_ln94_fu_117_p2 + j);

assign add_ln96_fu_253_p2 = (outputChanIdx_5 + 16'd1);

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign bitcast_ln94_10_fu_220_p1 = ap_sig_allocacmp_outputRow_11_1_load;

assign bitcast_ln94_11_fu_228_p1 = ap_sig_allocacmp_outputRow_11_2_load;

assign bitcast_ln94_12_fu_236_p1 = ap_sig_allocacmp_outputRow_11_3_load;

assign bitcast_ln94_fu_212_p1 = ap_sig_allocacmp_outputRow_11_0_load;

assign icmp_ln88_fu_179_p2 = ((add_ln87_fu_173_p2 == 16'd4) ? 1'b1 : 1'b0);

assign icmp_ln97_fu_259_p2 = ((add_ln96_fu_253_p2 == 16'd32) ? 1'b1 : 1'b0);

assign out_data_address1 = zext_ln94_8_fu_207_p1;

assign out_data_d1 = {{{{bitcast_ln94_12_fu_236_p1}, {bitcast_ln94_11_fu_228_p1}}, {bitcast_ln94_10_fu_220_p1}}, {bitcast_ln94_fu_212_p1}};

assign select_ln97_fu_265_p3 = ((icmp_ln97_fu_259_p2[0:0] == 1'b1) ? 16'd0 : add_ln96_fu_253_p2);

assign sub_ln94_fu_117_p2 = (tmp_fu_97_p3 - zext_ln94_fu_113_p1);

assign tmp_60_cast_fu_129_p3 = {{add_ln94_fu_123_p2}, {5'd0}};

assign tmp_fu_97_p3 = {{i}, {5'd0}};

assign tmp_s_fu_105_p3 = {{i}, {2'd0}};

assign trunc_ln86_fu_145_p1 = outputCount_5[1:0];

assign trunc_ln94_fu_193_p1 = outputChanIdx_5[6:0];

assign zext_ln94_7_fu_197_p1 = trunc_ln94_fu_193_p1;

assign zext_ln94_8_fu_207_p1 = add_ln94_4_fu_201_p2;

assign zext_ln94_fu_113_p1 = tmp_s_fu_105_p3;

endmodule //td_fused_top_tdf5_writeOutputs_unaligned
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf6_19 (
        in_data_address0,
        in_data_ce0,
        in_data_d0,
        in_data_q0,
        in_data_we0,
        in_data_address1,
        in_data_ce1,
        in_data_d1,
        in_data_q1,
        in_data_we1,
        out_data_address0,
        out_data_ce0,
        out_data_d0,
        out_data_q0,
        out_data_we0,
        out_data_address1,
        out_data_ce1,
        out_data_d1,
        out_data_q1,
        out_data_we1,
        filter_data_address0,
        filter_data_ce0,
        filter_data_d0,
        filter_data_q0,
        filter_data_we0,
        filter_data_address1,
        filter_data_ce1,
        filter_data_d1,
        filter_data_q1,
        filter_data_we1,
        adjustments_address0,
        adjustments_ce0,
        adjustments_d0,
        adjustments_q0,
        adjustments_we0,
        adjustments_address1,
        adjustments_ce1,
        adjustments_d1,
        adjustments_q1,
        adjustments_we1,
        ap_clk,
        ap_rst,
        in_data_empty_n,
        in_data_read,
        out_data_full_n,
        out_data_write,
        ap_start,
        ap_done,
        ap_ready,
        ap_idle,
        ap_continue
);


output  [14:0] in_data_address0;
output   in_data_ce0;
output  [63:0] in_data_d0;
input  [63:0] in_data_q0;
output   in_data_we0;
output  [14:0] in_data_address1;
output   in_data_ce1;
output  [63:0] in_data_d1;
input  [63:0] in_data_q1;
output   in_data_we1;
output  [12:0] out_data_address0;
output   out_data_ce0;
output  [63:0] out_data_d0;
input  [63:0] out_data_q0;
output   out_data_we0;
output  [12:0] out_data_address1;
output   out_data_ce1;
output  [63:0] out_data_d1;
input  [63:0] out_data_q1;
output   out_data_we1;
output  [11:0] filter_data_address0;
output   filter_data_ce0;
output  [15:0] filter_data_d0;
input  [15:0] filter_data_q0;
output   filter_data_we0;
output  [11:0] filter_data_address1;
output   filter_data_ce1;
output  [15:0] filter_data_d1;
input  [15:0] filter_data_q1;
output   filter_data_we1;
output  [4:0] adjustments_address0;
output   adjustments_ce0;
output  [47:0] adjustments_d0;
input  [47:0] adjustments_q0;
output   adjustments_we0;
output  [4:0] adjustments_address1;
output   adjustments_ce1;
output  [47:0] adjustments_d1;
input  [47:0] adjustments_q1;
output   adjustments_we1;
input   ap_clk;
input   ap_rst;
input   in_data_empty_n;
output   in_data_read;
input   out_data_full_n;
output   out_data_write;
input   ap_start;
output   ap_done;
output   ap_ready;
output   ap_idle;
input   ap_continue;

reg ap_done;
reg ap_ready;
reg ap_idle;

wire   [14:0] dataflow_in_loop_TOP_LOOP37644_U0_in_data_address0;
wire    dataflow_in_loop_TOP_LOOP37644_U0_in_data_ce0;
wire   [63:0] dataflow_in_loop_TOP_LOOP37644_U0_in_data_d0;
wire    dataflow_in_loop_TOP_LOOP37644_U0_in_data_we0;
wire   [14:0] dataflow_in_loop_TOP_LOOP37644_U0_in_data_address1;
wire    dataflow_in_loop_TOP_LOOP37644_U0_in_data_ce1;
wire   [63:0] dataflow_in_loop_TOP_LOOP37644_U0_in_data_d1;
wire    dataflow_in_loop_TOP_LOOP37644_U0_in_data_we1;
wire   [11:0] dataflow_in_loop_TOP_LOOP37644_U0_filter_data_address0;
wire    dataflow_in_loop_TOP_LOOP37644_U0_filter_data_ce0;
wire   [15:0] dataflow_in_loop_TOP_LOOP37644_U0_filter_data_d0;
wire    dataflow_in_loop_TOP_LOOP37644_U0_filter_data_we0;
wire   [11:0] dataflow_in_loop_TOP_LOOP37644_U0_filter_data_address1;
wire    dataflow_in_loop_TOP_LOOP37644_U0_filter_data_ce1;
wire   [15:0] dataflow_in_loop_TOP_LOOP37644_U0_filter_data_d1;
wire    dataflow_in_loop_TOP_LOOP37644_U0_filter_data_we1;
wire   [4:0] dataflow_in_loop_TOP_LOOP37644_U0_adjustments_address0;
wire    dataflow_in_loop_TOP_LOOP37644_U0_adjustments_ce0;
wire   [47:0] dataflow_in_loop_TOP_LOOP37644_U0_adjustments_d0;
wire    dataflow_in_loop_TOP_LOOP37644_U0_adjustments_we0;
wire   [4:0] dataflow_in_loop_TOP_LOOP37644_U0_adjustments_address1;
wire    dataflow_in_loop_TOP_LOOP37644_U0_adjustments_ce1;
wire   [47:0] dataflow_in_loop_TOP_LOOP37644_U0_adjustments_d1;
wire    dataflow_in_loop_TOP_LOOP37644_U0_adjustments_we1;
wire   [12:0] dataflow_in_loop_TOP_LOOP37644_U0_out_data_address0;
wire    dataflow_in_loop_TOP_LOOP37644_U0_out_data_ce0;
wire   [63:0] dataflow_in_loop_TOP_LOOP37644_U0_out_data_d0;
wire    dataflow_in_loop_TOP_LOOP37644_U0_out_data_we0;
wire   [12:0] dataflow_in_loop_TOP_LOOP37644_U0_out_data_address1;
wire    dataflow_in_loop_TOP_LOOP37644_U0_out_data_ce1;
wire   [63:0] dataflow_in_loop_TOP_LOOP37644_U0_out_data_d1;
wire    dataflow_in_loop_TOP_LOOP37644_U0_out_data_we1;
wire    dataflow_in_loop_TOP_LOOP37644_U0_ap_start;
wire    dataflow_in_loop_TOP_LOOP37644_U0_in_data_read;
wire    dataflow_in_loop_TOP_LOOP37644_U0_out_data_write;
wire    dataflow_in_loop_TOP_LOOP37644_U0_ap_done;
wire    dataflow_in_loop_TOP_LOOP37644_U0_ap_ready;
wire    dataflow_in_loop_TOP_LOOP37644_U0_ap_idle;
reg    dataflow_in_loop_TOP_LOOP37644_U0_ap_continue;
wire    dataflow_in_loop_TOP_LOOP37644_U0_in_data_full_n;
wire    dataflow_in_loop_TOP_LOOP37644_U0_in_data_write;
wire    ap_sync_continue;
wire    ap_sync_done;
wire    ap_sync_ready;
reg   [14:0] loop_dataflow_input_count;
reg   [14:0] loop_dataflow_output_count;
wire   [14:0] bound_minus_1;
wire    dataflow_in_loop_TOP_LOOP37644_U0_start_full_n;
wire    dataflow_in_loop_TOP_LOOP37644_U0_start_write;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 loop_dataflow_input_count = 15'd0;
#0 loop_dataflow_output_count = 15'd0;
end

td_fused_top_dataflow_in_loop_TOP_LOOP37644 dataflow_in_loop_TOP_LOOP37644_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .in_data_address0(dataflow_in_loop_TOP_LOOP37644_U0_in_data_address0),
    .in_data_ce0(dataflow_in_loop_TOP_LOOP37644_U0_in_data_ce0),
    .in_data_d0(dataflow_in_loop_TOP_LOOP37644_U0_in_data_d0),
    .in_data_q0(in_data_q0),
    .in_data_we0(dataflow_in_loop_TOP_LOOP37644_U0_in_data_we0),
    .in_data_address1(dataflow_in_loop_TOP_LOOP37644_U0_in_data_address1),
    .in_data_ce1(dataflow_in_loop_TOP_LOOP37644_U0_in_data_ce1),
    .in_data_d1(dataflow_in_loop_TOP_LOOP37644_U0_in_data_d1),
    .in_data_q1(64'd0),
    .in_data_we1(dataflow_in_loop_TOP_LOOP37644_U0_in_data_we1),
    .filter_data_address0(dataflow_in_loop_TOP_LOOP37644_U0_filter_data_address0),
    .filter_data_ce0(dataflow_in_loop_TOP_LOOP37644_U0_filter_data_ce0),
    .filter_data_d0(dataflow_in_loop_TOP_LOOP37644_U0_filter_data_d0),
    .filter_data_q0(filter_data_q0),
    .filter_data_we0(dataflow_in_loop_TOP_LOOP37644_U0_filter_data_we0),
    .filter_data_address1(dataflow_in_loop_TOP_LOOP37644_U0_filter_data_address1),
    .filter_data_ce1(dataflow_in_loop_TOP_LOOP37644_U0_filter_data_ce1),
    .filter_data_d1(dataflow_in_loop_TOP_LOOP37644_U0_filter_data_d1),
    .filter_data_q1(16'd0),
    .filter_data_we1(dataflow_in_loop_TOP_LOOP37644_U0_filter_data_we1),
    .adjustments_address0(dataflow_in_loop_TOP_LOOP37644_U0_adjustments_address0),
    .adjustments_ce0(dataflow_in_loop_TOP_LOOP37644_U0_adjustments_ce0),
    .adjustments_d0(dataflow_in_loop_TOP_LOOP37644_U0_adjustments_d0),
    .adjustments_q0(adjustments_q0),
    .adjustments_we0(dataflow_in_loop_TOP_LOOP37644_U0_adjustments_we0),
    .adjustments_address1(dataflow_in_loop_TOP_LOOP37644_U0_adjustments_address1),
    .adjustments_ce1(dataflow_in_loop_TOP_LOOP37644_U0_adjustments_ce1),
    .adjustments_d1(dataflow_in_loop_TOP_LOOP37644_U0_adjustments_d1),
    .adjustments_q1(48'd0),
    .adjustments_we1(dataflow_in_loop_TOP_LOOP37644_U0_adjustments_we1),
    .out_data_address0(dataflow_in_loop_TOP_LOOP37644_U0_out_data_address0),
    .out_data_ce0(dataflow_in_loop_TOP_LOOP37644_U0_out_data_ce0),
    .out_data_d0(dataflow_in_loop_TOP_LOOP37644_U0_out_data_d0),
    .out_data_q0(64'd0),
    .out_data_we0(dataflow_in_loop_TOP_LOOP37644_U0_out_data_we0),
    .out_data_address1(dataflow_in_loop_TOP_LOOP37644_U0_out_data_address1),
    .out_data_ce1(dataflow_in_loop_TOP_LOOP37644_U0_out_data_ce1),
    .out_data_d1(dataflow_in_loop_TOP_LOOP37644_U0_out_data_d1),
    .out_data_q1(64'd0),
    .out_data_we1(dataflow_in_loop_TOP_LOOP37644_U0_out_data_we1),
    .ap_start(dataflow_in_loop_TOP_LOOP37644_U0_ap_start),
    .in_data_empty_n(1'b0),
    .in_data_read(dataflow_in_loop_TOP_LOOP37644_U0_in_data_read),
    .out_data_full_n(out_data_full_n),
    .out_data_write(dataflow_in_loop_TOP_LOOP37644_U0_out_data_write),
    .ap_done(dataflow_in_loop_TOP_LOOP37644_U0_ap_done),
    .ap_ready(dataflow_in_loop_TOP_LOOP37644_U0_ap_ready),
    .ap_idle(dataflow_in_loop_TOP_LOOP37644_U0_ap_idle),
    .ap_continue(dataflow_in_loop_TOP_LOOP37644_U0_ap_continue)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        loop_dataflow_input_count <= 15'd0;
    end else begin
        if ((~(loop_dataflow_input_count == bound_minus_1) & (dataflow_in_loop_TOP_LOOP37644_U0_ap_ready == 1'b1) & (ap_start == 1'b1))) begin
            loop_dataflow_input_count <= (loop_dataflow_input_count + 15'd1);
        end else if (((dataflow_in_loop_TOP_LOOP37644_U0_ap_ready == 1'b1) & (loop_dataflow_input_count == bound_minus_1) & (ap_start == 1'b1))) begin
            loop_dataflow_input_count <= 15'd0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        loop_dataflow_output_count <= 15'd0;
    end else begin
        if ((~(loop_dataflow_output_count == bound_minus_1) & (dataflow_in_loop_TOP_LOOP37644_U0_ap_done == 1'b1) & (dataflow_in_loop_TOP_LOOP37644_U0_ap_continue == 1'b1))) begin
            loop_dataflow_output_count <= (loop_dataflow_output_count + 15'd1);
        end else if (((dataflow_in_loop_TOP_LOOP37644_U0_ap_done == 1'b1) & (loop_dataflow_output_count == bound_minus_1) & (dataflow_in_loop_TOP_LOOP37644_U0_ap_continue == 1'b1))) begin
            loop_dataflow_output_count <= 15'd0;
        end
    end
end

always @ (*) begin
    if (((dataflow_in_loop_TOP_LOOP37644_U0_ap_done == 1'b1) & (loop_dataflow_output_count == bound_minus_1))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = 1'b0;
    end
end

always @ (*) begin
    if (((dataflow_in_loop_TOP_LOOP37644_U0_ap_idle == 1'b1) & (loop_dataflow_output_count == 15'd0) & (ap_start == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((dataflow_in_loop_TOP_LOOP37644_U0_ap_ready == 1'b1) & (loop_dataflow_input_count == bound_minus_1) & (ap_start == 1'b1))) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((~(loop_dataflow_output_count == bound_minus_1) | (ap_continue == 1'b1))) begin
        dataflow_in_loop_TOP_LOOP37644_U0_ap_continue = 1'b1;
    end else begin
        dataflow_in_loop_TOP_LOOP37644_U0_ap_continue = 1'b0;
    end
end

assign adjustments_address0 = dataflow_in_loop_TOP_LOOP37644_U0_adjustments_address0;

assign adjustments_address1 = 5'd0;

assign adjustments_ce0 = dataflow_in_loop_TOP_LOOP37644_U0_adjustments_ce0;

assign adjustments_ce1 = 1'b0;

assign adjustments_d0 = 48'd0;

assign adjustments_d1 = 48'd0;

assign adjustments_we0 = 1'b0;

assign adjustments_we1 = 1'b0;

assign ap_sync_continue = ap_continue;

assign ap_sync_done = dataflow_in_loop_TOP_LOOP37644_U0_ap_done;

assign ap_sync_ready = dataflow_in_loop_TOP_LOOP37644_U0_ap_ready;

assign bound_minus_1 = (15'd25088 - 15'd1);

assign dataflow_in_loop_TOP_LOOP37644_U0_ap_start = ap_start;

assign dataflow_in_loop_TOP_LOOP37644_U0_in_data_full_n = in_data_empty_n;

assign dataflow_in_loop_TOP_LOOP37644_U0_in_data_write = 1'b0;

assign dataflow_in_loop_TOP_LOOP37644_U0_start_full_n = 1'b1;

assign dataflow_in_loop_TOP_LOOP37644_U0_start_write = 1'b0;

assign filter_data_address0 = dataflow_in_loop_TOP_LOOP37644_U0_filter_data_address0;

assign filter_data_address1 = 12'd0;

assign filter_data_ce0 = dataflow_in_loop_TOP_LOOP37644_U0_filter_data_ce0;

assign filter_data_ce1 = 1'b0;

assign filter_data_d0 = 16'd0;

assign filter_data_d1 = 16'd0;

assign filter_data_we0 = 1'b0;

assign filter_data_we1 = 1'b0;

assign in_data_address0 = dataflow_in_loop_TOP_LOOP37644_U0_in_data_address0;

assign in_data_address1 = 15'd0;

assign in_data_ce0 = dataflow_in_loop_TOP_LOOP37644_U0_in_data_ce0;

assign in_data_ce1 = 1'b0;

assign in_data_d0 = 64'd0;

assign in_data_d1 = 64'd0;

assign in_data_read = dataflow_in_loop_TOP_LOOP37644_U0_in_data_write;

assign in_data_we0 = 1'b0;

assign in_data_we1 = 1'b0;

assign out_data_address0 = 13'd0;

assign out_data_address1 = dataflow_in_loop_TOP_LOOP37644_U0_out_data_address1;

assign out_data_ce0 = 1'b0;

assign out_data_ce1 = dataflow_in_loop_TOP_LOOP37644_U0_out_data_ce1;

assign out_data_d0 = 64'd0;

assign out_data_d1 = dataflow_in_loop_TOP_LOOP37644_U0_out_data_d1;

assign out_data_we0 = 1'b0;

assign out_data_we1 = dataflow_in_loop_TOP_LOOP37644_U0_out_data_we1;

assign out_data_write = dataflow_in_loop_TOP_LOOP37644_U0_out_data_write;

endmodule //td_fused_top_tdf6_19
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf6_accum_1 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        accum_in_0_address0,
        accum_in_0_ce0,
        accum_in_0_q0,
        accum_in_0_address1,
        accum_in_0_ce1,
        accum_in_0_q1,
        accum_out_address0,
        accum_out_ce0,
        accum_out_we0,
        accum_out_d0,
        accum_out_address1,
        accum_out_ce1,
        accum_out_we1,
        accum_out_d1
);

parameter    ap_ST_fsm_state1 = 8'd1;
parameter    ap_ST_fsm_pp0_stage0 = 8'd2;
parameter    ap_ST_fsm_pp0_stage1 = 8'd4;
parameter    ap_ST_fsm_pp0_stage2 = 8'd8;
parameter    ap_ST_fsm_pp0_stage3 = 8'd16;
parameter    ap_ST_fsm_state12 = 8'd32;
parameter    ap_ST_fsm_state13 = 8'd64;
parameter    ap_ST_fsm_state14 = 8'd128;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [6:0] accum_in_0_address0;
output   accum_in_0_ce0;
input  [15:0] accum_in_0_q0;
output  [6:0] accum_in_0_address1;
output   accum_in_0_ce1;
input  [15:0] accum_in_0_q1;
output  [2:0] accum_out_address0;
output   accum_out_ce0;
output   accum_out_we0;
output  [15:0] accum_out_d0;
output  [2:0] accum_out_address1;
output   accum_out_ce1;
output   accum_out_we1;
output  [15:0] accum_out_d1;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg[6:0] accum_in_0_address0;
reg accum_in_0_ce0;
reg[6:0] accum_in_0_address1;
reg accum_in_0_ce1;
reg accum_out_ce0;
reg accum_out_we0;
reg accum_out_ce1;
reg accum_out_we1;

reg    ap_done_reg;
  reg   [7:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg   [7:0] x_reg_170;
reg   [15:0] psum_7_08_reg_182;
reg   [15:0] psum_6_07_reg_194;
reg   [15:0] psum_5_06_reg_206;
reg   [15:0] psum_4_05_reg_218;
reg   [15:0] psum_3_04_reg_230;
reg   [15:0] psum_2_03_reg_242;
reg   [15:0] psum_1_02_reg_254;
reg   [15:0] psum_0_01_reg_266;
wire   [0:0] tmp_fu_323_p3;
reg   [0:0] tmp_reg_494;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state6_pp0_stage0_iter1;
wire    ap_block_state10_pp0_stage0_iter2;
wire    ap_block_pp0_stage0_11001;
reg   [0:0] tmp_reg_494_pp0_iter1_reg;
reg   [0:0] tmp_reg_494_pp0_iter2_reg;
wire   [6:0] trunc_ln25_fu_336_p1;
reg   [6:0] trunc_ln25_reg_498;
reg   [15:0] accum_in_0_load_reg_518;
wire    ap_CS_fsm_pp0_stage1;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_state3_pp0_stage1_iter0;
wire    ap_block_state7_pp0_stage1_iter1;
wire    ap_block_state11_pp0_stage1_iter2;
wire    ap_block_pp0_stage1_11001;
reg   [15:0] accum_in_0_load_22_reg_523;
reg   [15:0] accum_in_0_load_23_reg_538;
wire    ap_CS_fsm_pp0_stage2;
wire    ap_block_state4_pp0_stage2_iter0;
wire    ap_block_state8_pp0_stage2_iter1;
wire    ap_block_pp0_stage2_11001;
reg   [15:0] accum_in_0_load_24_reg_543;
wire   [7:0] add_ln25_fu_391_p2;
reg   [7:0] add_ln25_reg_558;
wire    ap_CS_fsm_pp0_stage3;
wire    ap_block_state5_pp0_stage3_iter0;
wire    ap_block_state9_pp0_stage3_iter1;
wire    ap_block_pp0_stage3_11001;
reg   [15:0] accum_in_0_load_25_reg_563;
reg   [15:0] accum_in_0_load_26_reg_568;
reg   [15:0] accum_in_0_load_27_reg_583;
reg    ap_enable_reg_pp0_iter1;
reg   [15:0] accum_in_0_load_28_reg_588;
wire   [15:0] grp_fu_307_p2;
wire   [15:0] grp_fu_312_p2;
reg    ap_enable_reg_pp0_iter2;
wire   [3:0] add_ln33_fu_434_p2;
wire    ap_CS_fsm_state13;
wire   [0:0] tmp_19_fu_417_p3;
reg    ap_block_state1;
wire    ap_block_pp0_stage2_subdone;
reg    ap_condition_pp0_exit_iter0_state4;
wire    ap_block_pp0_stage3_subdone;
wire    ap_block_pp0_stage1_subdone;
reg   [7:0] ap_phi_mux_x_phi_fu_174_p4;
wire    ap_block_pp0_stage0;
wire   [15:0] ap_phi_mux_psum_7_08_phi_fu_186_p4;
wire    ap_block_pp0_stage1;
wire   [15:0] ap_phi_mux_psum_6_07_phi_fu_198_p4;
wire   [15:0] ap_phi_mux_psum_5_06_phi_fu_210_p4;
wire   [15:0] ap_phi_mux_psum_4_05_phi_fu_222_p4;
wire   [15:0] ap_phi_mux_psum_3_04_phi_fu_234_p4;
wire    ap_block_pp0_stage3;
wire   [15:0] ap_phi_mux_psum_2_03_phi_fu_246_p4;
wire    ap_block_pp0_stage2;
reg   [3:0] q_reg_278;
wire    ap_CS_fsm_state12;
reg   [15:0] ap_phi_mux_phi_ln45_phi_fu_292_p8;
wire   [2:0] trunc_ln33_fu_430_p1;
wire   [63:0] zext_ln25_fu_331_p1;
wire   [63:0] zext_ln29_fu_346_p1;
wire   [63:0] zext_ln29_7_fu_356_p1;
wire   [63:0] zext_ln29_8_fu_366_p1;
wire   [63:0] zext_ln29_9_fu_376_p1;
wire   [63:0] zext_ln29_10_fu_386_p1;
wire   [63:0] zext_ln29_11_fu_402_p1;
wire   [63:0] zext_ln29_12_fu_412_p1;
wire   [63:0] zext_ln33_fu_425_p1;
wire   [63:0] zext_ln33_2_fu_446_p1;
reg   [15:0] grp_fu_307_p0;
reg   [15:0] grp_fu_307_p1;
reg   [15:0] grp_fu_312_p0;
reg   [15:0] grp_fu_312_p1;
wire   [6:0] or_ln29_fu_340_p2;
wire   [6:0] or_ln29_7_fu_351_p2;
wire   [6:0] or_ln29_8_fu_361_p2;
wire   [6:0] or_ln29_9_fu_371_p2;
wire   [6:0] or_ln29_10_fu_381_p2;
wire   [6:0] or_ln29_11_fu_397_p2;
wire   [6:0] or_ln29_12_fu_407_p2;
wire   [2:0] or_ln33_fu_440_p2;
wire   [0:0] icmp_ln45_fu_451_p2;
wire   [0:0] icmp_ln45_3_fu_465_p2;
wire   [15:0] select_ln45_fu_457_p3;
wire   [0:0] icmp_ln45_4_fu_479_p2;
wire   [15:0] select_ln45_3_fu_471_p3;
wire    ap_CS_fsm_state14;
reg   [7:0] ap_NS_fsm;
wire    ap_block_pp0_stage0_subdone;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
reg    ap_condition_517;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 8'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
end

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U363(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(grp_fu_307_p0),
    .din1(grp_fu_307_p1),
    .dout(grp_fu_307_p2)
);

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U364(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(grp_fu_312_p0),
    .din1(grp_fu_312_p1),
    .dout(grp_fu_312_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state14)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage2_subdone) & (1'b1 == ap_condition_pp0_exit_iter0_state4) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage3_subdone) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b0)) | ((1'b0 == ap_block_pp0_stage3_subdone) & (1'b1 == ap_CS_fsm_pp0_stage3)))) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end else if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter2 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state12)) begin
        q_reg_278 <= 4'd0;
    end else if (((tmp_19_fu_417_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state13))) begin
        q_reg_278 <= add_ln33_fu_434_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (tmp_reg_494 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        x_reg_170 <= add_ln25_reg_558;
    end else if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        x_reg_170 <= 8'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage1_11001) & (tmp_reg_494 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
        accum_in_0_load_22_reg_523 <= accum_in_0_q0;
        accum_in_0_load_reg_518 <= accum_in_0_q1;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage2_11001) & (tmp_reg_494 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage2) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
        accum_in_0_load_23_reg_538 <= accum_in_0_q1;
        accum_in_0_load_24_reg_543 <= accum_in_0_q0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage3_11001) & (tmp_reg_494 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage3) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
        accum_in_0_load_25_reg_563 <= accum_in_0_q1;
        accum_in_0_load_26_reg_568 <= accum_in_0_q0;
        add_ln25_reg_558 <= add_ln25_fu_391_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (tmp_reg_494 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        accum_in_0_load_27_reg_583 <= accum_in_0_q1;
        accum_in_0_load_28_reg_588 <= accum_in_0_q0;
    end
end

always @ (posedge ap_clk) begin
    if (((tmp_reg_494_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage2_11001) & (1'b1 == ap_CS_fsm_pp0_stage2) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        psum_0_01_reg_266 <= grp_fu_307_p2;
        psum_1_02_reg_254 <= grp_fu_312_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((tmp_reg_494_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage3_11001) & (1'b1 == ap_CS_fsm_pp0_stage3) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        psum_2_03_reg_242 <= grp_fu_307_p2;
        psum_3_04_reg_230 <= grp_fu_312_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((tmp_reg_494_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        psum_4_05_reg_218 <= grp_fu_307_p2;
        psum_5_06_reg_206 <= grp_fu_312_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((tmp_reg_494_pp0_iter2_reg == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
        psum_6_07_reg_194 <= grp_fu_307_p2;
        psum_7_08_reg_182 <= grp_fu_312_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_reg_494 <= ap_phi_mux_x_phi_fu_174_p4[32'd7];
        tmp_reg_494_pp0_iter1_reg <= tmp_reg_494;
        tmp_reg_494_pp0_iter2_reg <= tmp_reg_494_pp0_iter1_reg;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (tmp_fu_323_p3 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        trunc_ln25_reg_498 <= trunc_ln25_fu_336_p1;
    end
end

always @ (*) begin
    if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
        if (((1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            accum_in_0_address0 = zext_ln29_12_fu_412_p1;
        end else if (((1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            accum_in_0_address0 = zext_ln29_10_fu_386_p1;
        end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            accum_in_0_address0 = zext_ln29_8_fu_366_p1;
        end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            accum_in_0_address0 = zext_ln29_fu_346_p1;
        end else begin
            accum_in_0_address0 = 'bx;
        end
    end else begin
        accum_in_0_address0 = 'bx;
    end
end

always @ (*) begin
    if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
        if (((1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            accum_in_0_address1 = zext_ln29_11_fu_402_p1;
        end else if (((1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            accum_in_0_address1 = zext_ln29_9_fu_376_p1;
        end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            accum_in_0_address1 = zext_ln29_7_fu_356_p1;
        end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            accum_in_0_address1 = zext_ln25_fu_331_p1;
        end else begin
            accum_in_0_address1 = 'bx;
        end
    end else begin
        accum_in_0_address1 = 'bx;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1)) | ((1'b0 == ap_block_pp0_stage3_11001) & (1'b1 == ap_CS_fsm_pp0_stage3) & (ap_enable_reg_pp0_iter0 == 1'b1)) | ((1'b0 == ap_block_pp0_stage2_11001) & (1'b1 == ap_CS_fsm_pp0_stage2) & (ap_enable_reg_pp0_iter0 == 1'b1)) | ((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1)))) begin
        accum_in_0_ce0 = 1'b1;
    end else begin
        accum_in_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1)) | ((1'b0 == ap_block_pp0_stage3_11001) & (1'b1 == ap_CS_fsm_pp0_stage3) & (ap_enable_reg_pp0_iter0 == 1'b1)) | ((1'b0 == ap_block_pp0_stage2_11001) & (1'b1 == ap_CS_fsm_pp0_stage2) & (ap_enable_reg_pp0_iter0 == 1'b1)) | ((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1)))) begin
        accum_in_0_ce1 = 1'b1;
    end else begin
        accum_in_0_ce1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state13)) begin
        accum_out_ce0 = 1'b1;
    end else begin
        accum_out_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state13)) begin
        accum_out_ce1 = 1'b1;
    end else begin
        accum_out_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((tmp_19_fu_417_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state13))) begin
        accum_out_we0 = 1'b1;
    end else begin
        accum_out_we0 = 1'b0;
    end
end

always @ (*) begin
    if (((tmp_19_fu_417_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state13))) begin
        accum_out_we1 = 1'b1;
    end else begin
        accum_out_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((tmp_reg_494 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state4 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state4 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state14)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((tmp_19_fu_417_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state13))) begin
        if ((trunc_ln33_fu_430_p1 == 3'd0)) begin
            ap_phi_mux_phi_ln45_phi_fu_292_p8 = psum_0_01_reg_266;
        end else if ((1'b1 == ap_condition_517)) begin
            ap_phi_mux_phi_ln45_phi_fu_292_p8 = psum_6_07_reg_194;
        end else if ((trunc_ln33_fu_430_p1 == 3'd4)) begin
            ap_phi_mux_phi_ln45_phi_fu_292_p8 = psum_4_05_reg_218;
        end else if ((trunc_ln33_fu_430_p1 == 3'd2)) begin
            ap_phi_mux_phi_ln45_phi_fu_292_p8 = psum_2_03_reg_242;
        end else begin
            ap_phi_mux_phi_ln45_phi_fu_292_p8 = 'bx;
        end
    end else begin
        ap_phi_mux_phi_ln45_phi_fu_292_p8 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0) & (tmp_reg_494 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_x_phi_fu_174_p4 = add_ln25_reg_558;
    end else begin
        ap_phi_mux_x_phi_fu_174_p4 = x_reg_170;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state14)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_307_p0 = ap_phi_mux_psum_6_07_phi_fu_198_p4;
    end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_307_p0 = ap_phi_mux_psum_4_05_phi_fu_222_p4;
    end else if (((1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
        grp_fu_307_p0 = ap_phi_mux_psum_2_03_phi_fu_246_p4;
    end else if (((1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
        grp_fu_307_p0 = grp_fu_307_p2;
    end else begin
        grp_fu_307_p0 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_307_p1 = accum_in_0_load_27_reg_583;
    end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_307_p1 = accum_in_0_load_25_reg_563;
    end else if (((1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
        grp_fu_307_p1 = accum_in_0_load_23_reg_538;
    end else if (((1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
        grp_fu_307_p1 = accum_in_0_load_reg_518;
    end else begin
        grp_fu_307_p1 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_312_p0 = ap_phi_mux_psum_7_08_phi_fu_186_p4;
    end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_312_p0 = ap_phi_mux_psum_5_06_phi_fu_210_p4;
    end else if (((1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
        grp_fu_312_p0 = ap_phi_mux_psum_3_04_phi_fu_234_p4;
    end else if (((1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
        grp_fu_312_p0 = grp_fu_312_p2;
    end else begin
        grp_fu_312_p0 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_312_p1 = accum_in_0_load_28_reg_588;
    end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_312_p1 = accum_in_0_load_26_reg_568;
    end else if (((1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
        grp_fu_312_p1 = accum_in_0_load_24_reg_543;
    end else if (((1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
        grp_fu_312_p1 = accum_in_0_load_22_reg_523;
    end else begin
        grp_fu_312_p1 = 'bx;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_pp0_stage1 : begin
            if ((~((1'b0 == ap_block_pp0_stage1_subdone) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b0)) & (1'b0 == ap_block_pp0_stage1_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage2;
            end else if (((1'b0 == ap_block_pp0_stage1_subdone) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
                ap_NS_fsm = ap_ST_fsm_state12;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end
        end
        ap_ST_fsm_pp0_stage2 : begin
            if ((~((1'b0 == ap_block_pp0_stage2_subdone) & (tmp_reg_494 == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1)) & (1'b0 == ap_block_pp0_stage2_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage3;
            end else if (((1'b0 == ap_block_pp0_stage2_subdone) & (tmp_reg_494 == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
                ap_NS_fsm = ap_ST_fsm_state12;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage2;
            end
        end
        ap_ST_fsm_pp0_stage3 : begin
            if ((1'b0 == ap_block_pp0_stage3_subdone)) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage3;
            end
        end
        ap_ST_fsm_state12 : begin
            ap_NS_fsm = ap_ST_fsm_state13;
        end
        ap_ST_fsm_state13 : begin
            if (((tmp_19_fu_417_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state13))) begin
                ap_NS_fsm = ap_ST_fsm_state13;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state14;
            end
        end
        ap_ST_fsm_state14 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign accum_out_address0 = zext_ln33_2_fu_446_p1;

assign accum_out_address1 = zext_ln33_fu_425_p1;

assign accum_out_d0 = ((icmp_ln45_4_fu_479_p2[0:0] == 1'b1) ? psum_5_06_reg_206 : select_ln45_3_fu_471_p3);

assign accum_out_d1 = ap_phi_mux_phi_ln45_phi_fu_292_p8;

assign add_ln25_fu_391_p2 = (x_reg_170 + 8'd8);

assign add_ln33_fu_434_p2 = (q_reg_278 + 4'd2);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_pp0_stage1 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_pp0_stage2 = ap_CS_fsm[32'd3];

assign ap_CS_fsm_pp0_stage3 = ap_CS_fsm[32'd4];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state12 = ap_CS_fsm[32'd5];

assign ap_CS_fsm_state13 = ap_CS_fsm[32'd6];

assign ap_CS_fsm_state14 = ap_CS_fsm[32'd7];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1_subdone = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage2 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage2_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage2_subdone = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage3 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage3_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage3_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((ap_done_reg == 1'b1) | (ap_start == 1'b0));
end

assign ap_block_state10_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state11_pp0_stage1_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage1_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage2_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage3_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage1_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage2_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state9_pp0_stage3_iter1 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_condition_517 = (~(trunc_ln33_fu_430_p1 == 3'd0) & ~(trunc_ln33_fu_430_p1 == 3'd4) & ~(trunc_ln33_fu_430_p1 == 3'd2));
end

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign ap_phi_mux_psum_2_03_phi_fu_246_p4 = grp_fu_307_p2;

assign ap_phi_mux_psum_3_04_phi_fu_234_p4 = grp_fu_312_p2;

assign ap_phi_mux_psum_4_05_phi_fu_222_p4 = grp_fu_307_p2;

assign ap_phi_mux_psum_5_06_phi_fu_210_p4 = grp_fu_312_p2;

assign ap_phi_mux_psum_6_07_phi_fu_198_p4 = grp_fu_307_p2;

assign ap_phi_mux_psum_7_08_phi_fu_186_p4 = grp_fu_312_p2;

assign icmp_ln45_3_fu_465_p2 = ((or_ln33_fu_440_p2 == 3'd3) ? 1'b1 : 1'b0);

assign icmp_ln45_4_fu_479_p2 = ((or_ln33_fu_440_p2 == 3'd5) ? 1'b1 : 1'b0);

assign icmp_ln45_fu_451_p2 = ((or_ln33_fu_440_p2 == 3'd1) ? 1'b1 : 1'b0);

assign or_ln29_10_fu_381_p2 = (trunc_ln25_reg_498 | 7'd5);

assign or_ln29_11_fu_397_p2 = (trunc_ln25_reg_498 | 7'd6);

assign or_ln29_12_fu_407_p2 = (trunc_ln25_reg_498 | 7'd7);

assign or_ln29_7_fu_351_p2 = (trunc_ln25_reg_498 | 7'd2);

assign or_ln29_8_fu_361_p2 = (trunc_ln25_reg_498 | 7'd3);

assign or_ln29_9_fu_371_p2 = (trunc_ln25_reg_498 | 7'd4);

assign or_ln29_fu_340_p2 = (trunc_ln25_fu_336_p1 | 7'd1);

assign or_ln33_fu_440_p2 = (trunc_ln33_fu_430_p1 | 3'd1);

assign select_ln45_3_fu_471_p3 = ((icmp_ln45_3_fu_465_p2[0:0] == 1'b1) ? psum_3_04_reg_230 : select_ln45_fu_457_p3);

assign select_ln45_fu_457_p3 = ((icmp_ln45_fu_451_p2[0:0] == 1'b1) ? psum_1_02_reg_254 : psum_7_08_reg_182);

assign tmp_19_fu_417_p3 = q_reg_278[32'd3];

assign tmp_fu_323_p3 = ap_phi_mux_x_phi_fu_174_p4[32'd7];

assign trunc_ln25_fu_336_p1 = ap_phi_mux_x_phi_fu_174_p4[6:0];

assign trunc_ln33_fu_430_p1 = q_reg_278[2:0];

assign zext_ln25_fu_331_p1 = ap_phi_mux_x_phi_fu_174_p4;

assign zext_ln29_10_fu_386_p1 = or_ln29_10_fu_381_p2;

assign zext_ln29_11_fu_402_p1 = or_ln29_11_fu_397_p2;

assign zext_ln29_12_fu_412_p1 = or_ln29_12_fu_407_p2;

assign zext_ln29_7_fu_356_p1 = or_ln29_7_fu_351_p2;

assign zext_ln29_8_fu_366_p1 = or_ln29_8_fu_361_p2;

assign zext_ln29_9_fu_376_p1 = or_ln29_9_fu_371_p2;

assign zext_ln29_fu_346_p1 = or_ln29_fu_340_p2;

assign zext_ln33_2_fu_446_p1 = or_ln33_fu_440_p2;

assign zext_ln33_fu_425_p1 = q_reg_278;

endmodule //td_fused_top_tdf6_accum_1
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf6_accum_2 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        accum_in_8,
        accum_in_8_ap_vld,
        accum_in_address0,
        accum_in_ce0,
        accum_in_q0
);

parameter    ap_ST_fsm_state1 = 7'd1;
parameter    ap_ST_fsm_state2 = 7'd2;
parameter    ap_ST_fsm_state3 = 7'd4;
parameter    ap_ST_fsm_state4 = 7'd8;
parameter    ap_ST_fsm_state5 = 7'd16;
parameter    ap_ST_fsm_state6 = 7'd32;
parameter    ap_ST_fsm_state7 = 7'd64;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [15:0] accum_in_8;
output   accum_in_8_ap_vld;
output  [2:0] accum_in_address0;
output   accum_in_ce0;
input  [15:0] accum_in_q0;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg[15:0] accum_in_8;
reg accum_in_8_ap_vld;
reg accum_in_ce0;

reg    ap_done_reg;
  reg   [6:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
wire   [3:0] add_ln57_fu_74_p2;
reg   [3:0] add_ln57_reg_91;
wire    ap_CS_fsm_state2;
wire   [0:0] icmp_ln57_fu_85_p2;
wire    ap_CS_fsm_state3;
wire   [15:0] grp_fu_68_p2;
wire    ap_CS_fsm_state7;
reg   [3:0] i_1_1_reg_44;
reg    ap_block_state1;
reg   [15:0] sum_01_reg_55;
wire   [63:0] zext_ln57_fu_80_p1;
reg   [15:0] accum_in_8_preg;
reg   [6:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 7'd1;
#0 accum_in_8_preg = 16'd0;
end

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U367(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(sum_01_reg_55),
    .din1(accum_in_q0),
    .dout(grp_fu_68_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        accum_in_8_preg <= 16'd0;
    end else begin
        if (((icmp_ln57_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
            accum_in_8_preg <= sum_01_reg_55;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if (((icmp_ln57_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        i_1_1_reg_44 <= 4'd0;
    end else if ((1'b1 == ap_CS_fsm_state7)) begin
        i_1_1_reg_44 <= add_ln57_reg_91;
    end
end

always @ (posedge ap_clk) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        sum_01_reg_55 <= 16'd0;
    end else if ((1'b1 == ap_CS_fsm_state7)) begin
        sum_01_reg_55 <= grp_fu_68_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        add_ln57_reg_91 <= add_ln57_fu_74_p2;
    end
end

always @ (*) begin
    if (((icmp_ln57_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        accum_in_8 = sum_01_reg_55;
    end else begin
        accum_in_8 = accum_in_8_preg;
    end
end

always @ (*) begin
    if (((icmp_ln57_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        accum_in_8_ap_vld = 1'b1;
    end else begin
        accum_in_8_ap_vld = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        accum_in_ce0 = 1'b1;
    end else begin
        accum_in_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln57_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln57_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_state2 : begin
            if (((icmp_ln57_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end
        end
        ap_ST_fsm_state3 : begin
            ap_NS_fsm = ap_ST_fsm_state4;
        end
        ap_ST_fsm_state4 : begin
            ap_NS_fsm = ap_ST_fsm_state5;
        end
        ap_ST_fsm_state5 : begin
            ap_NS_fsm = ap_ST_fsm_state6;
        end
        ap_ST_fsm_state6 : begin
            ap_NS_fsm = ap_ST_fsm_state7;
        end
        ap_ST_fsm_state7 : begin
            ap_NS_fsm = ap_ST_fsm_state2;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign accum_in_address0 = zext_ln57_fu_80_p1;

assign add_ln57_fu_74_p2 = (i_1_1_reg_44 + 4'd1);

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state7 = ap_CS_fsm[32'd6];

always @ (*) begin
    ap_block_state1 = ((ap_done_reg == 1'b1) | (ap_start == 1'b0));
end

assign icmp_ln57_fu_85_p2 = ((i_1_1_reg_44 == 4'd8) ? 1'b1 : 1'b0);

assign zext_ln57_fu_80_p1 = i_1_1_reg_44;

endmodule //td_fused_top_tdf6_accum_2
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf6_adjust (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        sums_read,
        adjustments_address0,
        adjustments_ce0,
        adjustments_q0,
        indices_23_dout,
        indices_23_empty_n,
        indices_23_read,
        ap_return
);

parameter    ap_ST_fsm_state1 = 17'd1;
parameter    ap_ST_fsm_state2 = 17'd2;
parameter    ap_ST_fsm_state3 = 17'd4;
parameter    ap_ST_fsm_state4 = 17'd8;
parameter    ap_ST_fsm_state5 = 17'd16;
parameter    ap_ST_fsm_state6 = 17'd32;
parameter    ap_ST_fsm_state7 = 17'd64;
parameter    ap_ST_fsm_state8 = 17'd128;
parameter    ap_ST_fsm_state9 = 17'd256;
parameter    ap_ST_fsm_state10 = 17'd512;
parameter    ap_ST_fsm_state11 = 17'd1024;
parameter    ap_ST_fsm_state12 = 17'd2048;
parameter    ap_ST_fsm_state13 = 17'd4096;
parameter    ap_ST_fsm_state14 = 17'd8192;
parameter    ap_ST_fsm_state15 = 17'd16384;
parameter    ap_ST_fsm_state16 = 17'd32768;
parameter    ap_ST_fsm_state17 = 17'd65536;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
input  [15:0] sums_read;
output  [4:0] adjustments_address0;
output   adjustments_ce0;
input  [47:0] adjustments_q0;
input  [4:0] indices_23_dout;
input   indices_23_empty_n;
output   indices_23_read;
output  [15:0] ap_return;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg adjustments_ce0;
reg indices_23_read;

reg    ap_done_reg;
  reg   [16:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    indices_23_blk_n;
wire    ap_CS_fsm_state4;
reg   [15:0] tmp_34_i_i_reg_167;
reg   [15:0] tmp_35_i_i_reg_172;
wire   [15:0] grp_fu_81_p2;
reg   [15:0] sub_i_i_i_reg_177;
wire    ap_CS_fsm_state8;
wire    ap_CS_fsm_state9;
wire   [15:0] grp_fu_86_p2;
reg   [15:0] mul_i_i_i_reg_187;
wire    ap_CS_fsm_state12;
wire    ap_CS_fsm_state13;
wire   [63:0] zext_ln220_fu_90_p1;
reg    ap_block_state1;
wire    ap_CS_fsm_state2;
wire    ap_CS_fsm_state3;
wire   [15:0] grp_fu_77_p1;
wire   [15:0] grp_fu_81_p1;
wire   [15:0] grp_fu_86_p1;
wire   [15:0] trunc_ln220_fu_95_p1;
wire   [15:0] grp_fu_77_p2;
wire    ap_CS_fsm_state17;
wire   [15:0] bitcast_ln648_fu_132_p1;
wire   [0:0] tmp_fu_136_p3;
reg   [16:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 17'd1;
end

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U371(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(mul_i_i_i_reg_187),
    .din1(grp_fu_77_p1),
    .dout(grp_fu_77_p2)
);

td_fused_top_hsub_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hsub_16ns_16ns_16_5_full_dsp_1_U372(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(sums_read),
    .din1(grp_fu_81_p1),
    .dout(grp_fu_81_p2)
);

td_fused_top_hmul_16ns_16ns_16_4_max_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hmul_16ns_16ns_16_4_max_dsp_1_U373(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(sub_i_i_i_reg_177),
    .din1(grp_fu_86_p1),
    .dout(grp_fu_86_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state17)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state12)) begin
        mul_i_i_i_reg_187 <= grp_fu_86_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state8)) begin
        sub_i_i_i_reg_177 <= grp_fu_81_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        tmp_34_i_i_reg_167 <= {{adjustments_q0[31:16]}};
        tmp_35_i_i_reg_172 <= {{adjustments_q0[47:32]}};
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state2) | (~((indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1)))) begin
        adjustments_ce0 = 1'b1;
    end else begin
        adjustments_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state17)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state17)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_23_blk_n = indices_23_empty_n;
    end else begin
        indices_23_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_23_read = 1'b1;
    end else begin
        indices_23_read = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_state2 : begin
            ap_NS_fsm = ap_ST_fsm_state3;
        end
        ap_ST_fsm_state3 : begin
            ap_NS_fsm = ap_ST_fsm_state4;
        end
        ap_ST_fsm_state4 : begin
            ap_NS_fsm = ap_ST_fsm_state5;
        end
        ap_ST_fsm_state5 : begin
            ap_NS_fsm = ap_ST_fsm_state6;
        end
        ap_ST_fsm_state6 : begin
            ap_NS_fsm = ap_ST_fsm_state7;
        end
        ap_ST_fsm_state7 : begin
            ap_NS_fsm = ap_ST_fsm_state8;
        end
        ap_ST_fsm_state8 : begin
            ap_NS_fsm = ap_ST_fsm_state9;
        end
        ap_ST_fsm_state9 : begin
            ap_NS_fsm = ap_ST_fsm_state10;
        end
        ap_ST_fsm_state10 : begin
            ap_NS_fsm = ap_ST_fsm_state11;
        end
        ap_ST_fsm_state11 : begin
            ap_NS_fsm = ap_ST_fsm_state12;
        end
        ap_ST_fsm_state12 : begin
            ap_NS_fsm = ap_ST_fsm_state13;
        end
        ap_ST_fsm_state13 : begin
            ap_NS_fsm = ap_ST_fsm_state14;
        end
        ap_ST_fsm_state14 : begin
            ap_NS_fsm = ap_ST_fsm_state15;
        end
        ap_ST_fsm_state15 : begin
            ap_NS_fsm = ap_ST_fsm_state16;
        end
        ap_ST_fsm_state16 : begin
            ap_NS_fsm = ap_ST_fsm_state17;
        end
        ap_ST_fsm_state17 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign adjustments_address0 = zext_ln220_fu_90_p1;

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state12 = ap_CS_fsm[32'd11];

assign ap_CS_fsm_state13 = ap_CS_fsm[32'd12];

assign ap_CS_fsm_state17 = ap_CS_fsm[32'd16];

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

assign ap_CS_fsm_state8 = ap_CS_fsm[32'd7];

assign ap_CS_fsm_state9 = ap_CS_fsm[32'd8];

always @ (*) begin
    ap_block_state1 = ((indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0));
end

assign ap_return = ((tmp_fu_136_p3[0:0] == 1'b1) ? 16'd0 : grp_fu_77_p2);

assign bitcast_ln648_fu_132_p1 = grp_fu_77_p2;

assign grp_fu_77_p1 = tmp_35_i_i_reg_172;

assign grp_fu_81_p1 = trunc_ln220_fu_95_p1;

assign grp_fu_86_p1 = tmp_34_i_i_reg_167;

assign tmp_fu_136_p3 = bitcast_ln648_fu_132_p1[32'd15];

assign trunc_ln220_fu_95_p1 = adjustments_q0[15:0];

assign zext_ln220_fu_90_p1 = indices_23_dout;

endmodule //td_fused_top_tdf6_adjust
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf6_dot_product (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        ifmap_vec_0_0_address0,
        ifmap_vec_0_0_ce0,
        ifmap_vec_0_0_q0,
        weight_vecs_0_0_0_address0,
        weight_vecs_0_0_0_ce0,
        weight_vecs_0_0_0_q0,
        products_0_address0,
        products_0_ce0,
        products_0_we0,
        products_0_d0
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state9 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [6:0] ifmap_vec_0_0_address0;
output   ifmap_vec_0_0_ce0;
input  [15:0] ifmap_vec_0_0_q0;
output  [6:0] weight_vecs_0_0_0_address0;
output   weight_vecs_0_0_0_ce0;
input  [15:0] weight_vecs_0_0_0_q0;
output  [6:0] products_0_address0;
output   products_0_ce0;
output   products_0_we0;
output  [15:0] products_0_d0;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg ifmap_vec_0_0_ce0;
reg weight_vecs_0_0_0_ce0;
reg products_0_ce0;
reg products_0_we0;

reg    ap_done_reg;
  reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg   [7:0] ic_0_0_reg_69;
wire   [7:0] add_ln149_fu_84_p2;
wire    ap_CS_fsm_pp0_stage0;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
wire    ap_block_state4_pp0_stage0_iter2;
wire    ap_block_state5_pp0_stage0_iter3;
wire    ap_block_state6_pp0_stage0_iter4;
wire    ap_block_state7_pp0_stage0_iter5;
wire    ap_block_state8_pp0_stage0_iter6;
wire    ap_block_pp0_stage0_11001;
wire   [0:0] icmp_ln149_fu_90_p2;
reg   [0:0] icmp_ln149_reg_107;
reg   [0:0] icmp_ln149_reg_107_pp0_iter1_reg;
reg   [0:0] icmp_ln149_reg_107_pp0_iter2_reg;
reg   [0:0] icmp_ln149_reg_107_pp0_iter3_reg;
reg   [0:0] icmp_ln149_reg_107_pp0_iter4_reg;
reg   [0:0] icmp_ln149_reg_107_pp0_iter5_reg;
wire   [63:0] idxprom17_0_0_fu_96_p1;
reg   [63:0] idxprom17_0_0_reg_111;
reg   [63:0] idxprom17_0_0_reg_111_pp0_iter1_reg;
reg   [63:0] idxprom17_0_0_reg_111_pp0_iter2_reg;
reg   [63:0] idxprom17_0_0_reg_111_pp0_iter3_reg;
reg   [63:0] idxprom17_0_0_reg_111_pp0_iter4_reg;
reg   [63:0] idxprom17_0_0_reg_111_pp0_iter5_reg;
reg   [15:0] ifmap_vec_0_0_load_reg_126;
reg   [15:0] weight_vecs_0_0_0_load_reg_131;
wire   [15:0] grp_fu_80_p2;
reg   [15:0] mul_reg_136;
reg    ap_block_state1;
wire    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_exit_iter0_state2;
reg    ap_enable_reg_pp0_iter1;
reg    ap_enable_reg_pp0_iter2;
reg    ap_enable_reg_pp0_iter3;
reg    ap_enable_reg_pp0_iter4;
reg    ap_enable_reg_pp0_iter5;
reg    ap_enable_reg_pp0_iter6;
wire    ap_block_pp0_stage0;
wire    ap_CS_fsm_state9;
reg   [2:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
#0 ap_enable_reg_pp0_iter4 = 1'b0;
#0 ap_enable_reg_pp0_iter5 = 1'b0;
#0 ap_enable_reg_pp0_iter6 = 1'b0;
end

td_fused_top_hmul_16ns_16ns_16_4_max_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hmul_16ns_16ns_16_4_max_dsp_1_U359(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(ifmap_vec_0_0_load_reg_126),
    .din1(weight_vecs_0_0_0_load_reg_131),
    .dout(grp_fu_80_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b1 == ap_condition_pp0_exit_iter0_state2))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            if ((1'b1 == ap_condition_pp0_exit_iter0_state2)) begin
                ap_enable_reg_pp0_iter1 <= (1'b1 ^ ap_condition_pp0_exit_iter0_state2);
            end else if ((1'b1 == 1'b1)) begin
                ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
            end
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter4 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter5 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter5 <= ap_enable_reg_pp0_iter4;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter6 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter6 <= ap_enable_reg_pp0_iter5;
        end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter6 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln149_fu_90_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ic_0_0_reg_69 <= add_ln149_fu_84_p2;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ic_0_0_reg_69 <= 8'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln149_reg_107 <= icmp_ln149_fu_90_p2;
        icmp_ln149_reg_107_pp0_iter1_reg <= icmp_ln149_reg_107;
        idxprom17_0_0_reg_111_pp0_iter1_reg[7 : 0] <= idxprom17_0_0_reg_111[7 : 0];
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        icmp_ln149_reg_107_pp0_iter2_reg <= icmp_ln149_reg_107_pp0_iter1_reg;
        icmp_ln149_reg_107_pp0_iter3_reg <= icmp_ln149_reg_107_pp0_iter2_reg;
        icmp_ln149_reg_107_pp0_iter4_reg <= icmp_ln149_reg_107_pp0_iter3_reg;
        icmp_ln149_reg_107_pp0_iter5_reg <= icmp_ln149_reg_107_pp0_iter4_reg;
        idxprom17_0_0_reg_111_pp0_iter2_reg[7 : 0] <= idxprom17_0_0_reg_111_pp0_iter1_reg[7 : 0];
        idxprom17_0_0_reg_111_pp0_iter3_reg[7 : 0] <= idxprom17_0_0_reg_111_pp0_iter2_reg[7 : 0];
        idxprom17_0_0_reg_111_pp0_iter4_reg[7 : 0] <= idxprom17_0_0_reg_111_pp0_iter3_reg[7 : 0];
        idxprom17_0_0_reg_111_pp0_iter5_reg[7 : 0] <= idxprom17_0_0_reg_111_pp0_iter4_reg[7 : 0];
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln149_fu_90_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        idxprom17_0_0_reg_111[7 : 0] <= idxprom17_0_0_fu_96_p1[7 : 0];
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln149_reg_107 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ifmap_vec_0_0_load_reg_126 <= ifmap_vec_0_0_q0;
        weight_vecs_0_0_0_load_reg_131 <= weight_vecs_0_0_0_q0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln149_reg_107_pp0_iter4_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        mul_reg_136 <= grp_fu_80_p2;
    end
end

always @ (*) begin
    if ((icmp_ln149_fu_90_p2 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state2 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state2 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state9)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state9)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ifmap_vec_0_0_ce0 = 1'b1;
    end else begin
        ifmap_vec_0_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter6 == 1'b1))) begin
        products_0_ce0 = 1'b1;
    end else begin
        products_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln149_reg_107_pp0_iter5_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter6 == 1'b1))) begin
        products_0_we0 = 1'b1;
    end else begin
        products_0_we0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        weight_vecs_0_0_0_ce0 = 1'b1;
    end else begin
        weight_vecs_0_0_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((~((icmp_ln149_fu_90_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0)) & ~((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter6 == 1'b1) & (ap_enable_reg_pp0_iter5 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if ((((icmp_ln149_fu_90_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0)) | ((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter6 == 1'b1) & (ap_enable_reg_pp0_iter5 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_state9;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state9 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln149_fu_84_p2 = (ic_0_0_reg_69 + 8'd1);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state9 = ap_CS_fsm[32'd2];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (ap_done_reg == 1'b1));
end

assign ap_block_state2_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter4 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage0_iter5 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage0_iter6 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign icmp_ln149_fu_90_p2 = ((ic_0_0_reg_69 == 8'd128) ? 1'b1 : 1'b0);

assign idxprom17_0_0_fu_96_p1 = ic_0_0_reg_69;

assign ifmap_vec_0_0_address0 = idxprom17_0_0_fu_96_p1;

assign products_0_address0 = idxprom17_0_0_reg_111_pp0_iter5_reg;

assign products_0_d0 = mul_reg_136;

assign weight_vecs_0_0_0_address0 = idxprom17_0_0_fu_96_p1;

always @ (posedge ap_clk) begin
    idxprom17_0_0_reg_111[63:8] <= 56'b00000000000000000000000000000000000000000000000000000000;
    idxprom17_0_0_reg_111_pp0_iter1_reg[63:8] <= 56'b00000000000000000000000000000000000000000000000000000000;
    idxprom17_0_0_reg_111_pp0_iter2_reg[63:8] <= 56'b00000000000000000000000000000000000000000000000000000000;
    idxprom17_0_0_reg_111_pp0_iter3_reg[63:8] <= 56'b00000000000000000000000000000000000000000000000000000000;
    idxprom17_0_0_reg_111_pp0_iter4_reg[63:8] <= 56'b00000000000000000000000000000000000000000000000000000000;
    idxprom17_0_0_reg_111_pp0_iter5_reg[63:8] <= 56'b00000000000000000000000000000000000000000000000000000000;
end

endmodule //td_fused_top_tdf6_dot_product
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_tdf6_filters_ram (addr0, ce0, q0, addr1, ce1, d1, we1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 12;
parameter MEM_SIZE = 4096;

input[AWIDTH-1:0] addr0;
input ce0;
output wire[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
input clk;

 reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];
wire [AWIDTH-1:0] addr0_t0; 
reg [AWIDTH-1:0] addr0_t1; 
reg [DWIDTH-1:0] q0_t0;
reg [DWIDTH-1:0] q0_t1;
wire [AWIDTH-1:0] addr1_t0; 
reg [AWIDTH-1:0] addr1_t1; 
wire [DWIDTH-1:0] d1_t0; 
wire we1_t0; 
reg [DWIDTH-1:0] d1_t1; 
reg we1_t1; 


assign addr0_t0 = addr0;
assign q0 = q0_t1;
assign addr1_t0 = addr1;
assign d1_t0 = d1;
assign we1_t0 = we1;

always @(posedge clk)  
begin
    if (ce0) 
    begin
        addr0_t1 <= addr0_t0; 
        q0_t1 <= q0_t0;
    end
    if (ce1) 
    begin
        addr1_t1 <= addr1_t0; 
        d1_t1 <= d1_t0;
        we1_t1 <= we1_t0;
    end
end


always @(posedge clk)  
begin 
    if (ce0) begin
        q0_t0 <= ram[addr0_t1];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1_t1) 
            ram[addr1_t1] <= d1_t1; 
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_tdf6_filters(
    reset,
    clk,
    address0,
    ce0,
    q0,
    address1,
    ce1,
    we1,
    d1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd4096;
parameter AddressWidth = 32'd12;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;



td_fused_top_tdf6_filters_ram td_fused_top_tdf6_filters_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 )
);

endmodule

// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf6_get_next_ijk (
        ap_clk,
        ap_rst,
        ap_start,
        start_full_n,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        start_out,
        start_write,
        indices_0_din,
        indices_0_full_n,
        indices_0_write,
        indices_1_din,
        indices_1_full_n,
        indices_1_write,
        indices_2_out_din,
        indices_2_out_full_n,
        indices_2_out_write,
        indices_2_out1_din,
        indices_2_out1_full_n,
        indices_2_out1_write
);

parameter    ap_ST_fsm_state1 = 1'd1;

input   ap_clk;
input   ap_rst;
input   ap_start;
input   start_full_n;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output   start_out;
output   start_write;
output  [15:0] indices_0_din;
input   indices_0_full_n;
output   indices_0_write;
output  [15:0] indices_1_din;
input   indices_1_full_n;
output   indices_1_write;
output  [4:0] indices_2_out_din;
input   indices_2_out_full_n;
output   indices_2_out_write;
output  [4:0] indices_2_out1_din;
input   indices_2_out1_full_n;
output   indices_2_out1_write;

reg ap_done;
reg ap_idle;
reg start_write;
reg indices_0_write;
reg indices_1_write;
reg indices_2_out_write;
reg indices_2_out1_write;

reg    real_start;
reg    start_once_reg;
reg    ap_done_reg;
  reg   [0:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    internal_ap_ready;
reg   [15:0] i_1;
reg   [15:0] j_1;
reg   [15:0] k_1;
reg    indices_0_blk_n;
reg    indices_1_blk_n;
reg    indices_2_out_blk_n;
reg    indices_2_out1_blk_n;
reg   [0:0] ap_phi_mux_j_17_flag_0_i_phi_fu_77_p6;
reg    ap_block_state1;
wire   [0:0] icmp_ln78_fu_141_p2;
wire   [0:0] icmp_ln81_fu_154_p2;
reg   [15:0] ap_phi_mux_j_17_new_0_i_phi_fu_91_p6;
wire   [15:0] add_ln80_fu_147_p2;
reg   [15:0] ap_phi_mux_k_17_new_0_i_phi_fu_104_p6;
wire   [15:0] add_ln77_fu_134_p2;
wire   [15:0] select_ln84_fu_172_p3;
wire   [4:0] trunc_ln76_fu_128_p1;
wire   [15:0] add_ln83_fu_160_p2;
wire   [0:0] icmp_ln84_fu_166_p2;
reg   [0:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 start_once_reg = 1'b0;
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 1'd1;
#0 i_1 = 16'd0;
#0 j_1 = 16'd0;
#0 k_1 = 16'd0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((~((real_start == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        start_once_reg <= 1'b0;
    end else begin
        if (((real_start == 1'b1) & (internal_ap_ready == 1'b0))) begin
            start_once_reg <= 1'b1;
        end else if ((internal_ap_ready == 1'b1)) begin
            start_once_reg <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((~((real_start == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (icmp_ln81_fu_154_p2 == 1'd1) & (icmp_ln78_fu_141_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1))) begin
        i_1 <= select_ln84_fu_172_p3;
    end
end

always @ (posedge ap_clk) begin
    if ((~((real_start == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (ap_phi_mux_j_17_flag_0_i_phi_fu_77_p6 == 1'd1) & (1'b1 == ap_CS_fsm_state1))) begin
        j_1 <= ap_phi_mux_j_17_new_0_i_phi_fu_91_p6;
    end
end

always @ (posedge ap_clk) begin
    if ((~((real_start == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        k_1 <= ap_phi_mux_k_17_new_0_i_phi_fu_104_p6;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((real_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln78_fu_141_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_phi_mux_j_17_flag_0_i_phi_fu_77_p6 = 1'd0;
    end else if ((((icmp_ln81_fu_154_p2 == 1'd0) & (icmp_ln78_fu_141_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1)) | ((icmp_ln81_fu_154_p2 == 1'd1) & (icmp_ln78_fu_141_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1)))) begin
        ap_phi_mux_j_17_flag_0_i_phi_fu_77_p6 = 1'd1;
    end else begin
        ap_phi_mux_j_17_flag_0_i_phi_fu_77_p6 = 'bx;
    end
end

always @ (*) begin
    if (((icmp_ln78_fu_141_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1))) begin
        if ((icmp_ln81_fu_154_p2 == 1'd0)) begin
            ap_phi_mux_j_17_new_0_i_phi_fu_91_p6 = add_ln80_fu_147_p2;
        end else if ((icmp_ln81_fu_154_p2 == 1'd1)) begin
            ap_phi_mux_j_17_new_0_i_phi_fu_91_p6 = 16'd0;
        end else begin
            ap_phi_mux_j_17_new_0_i_phi_fu_91_p6 = 'bx;
        end
    end else begin
        ap_phi_mux_j_17_new_0_i_phi_fu_91_p6 = 'bx;
    end
end

always @ (*) begin
    if (((icmp_ln78_fu_141_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_phi_mux_k_17_new_0_i_phi_fu_104_p6 = add_ln77_fu_134_p2;
    end else if ((((icmp_ln81_fu_154_p2 == 1'd0) & (icmp_ln78_fu_141_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1)) | ((icmp_ln81_fu_154_p2 == 1'd1) & (icmp_ln78_fu_141_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1)))) begin
        ap_phi_mux_k_17_new_0_i_phi_fu_104_p6 = 16'd0;
    end else begin
        ap_phi_mux_k_17_new_0_i_phi_fu_104_p6 = 'bx;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_0_blk_n = indices_0_full_n;
    end else begin
        indices_0_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_0_write = 1'b1;
    end else begin
        indices_0_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_1_blk_n = indices_1_full_n;
    end else begin
        indices_1_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_1_write = 1'b1;
    end else begin
        indices_1_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_2_out1_blk_n = indices_2_out1_full_n;
    end else begin
        indices_2_out1_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_2_out1_write = 1'b1;
    end else begin
        indices_2_out1_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_2_out_blk_n = indices_2_out_full_n;
    end else begin
        indices_2_out_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_2_out_write = 1'b1;
    end else begin
        indices_2_out_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        internal_ap_ready = 1'b1;
    end else begin
        internal_ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((start_full_n == 1'b0) & (start_once_reg == 1'b0))) begin
        real_start = 1'b0;
    end else begin
        real_start = ap_start;
    end
end

always @ (*) begin
    if (((real_start == 1'b1) & (start_once_reg == 1'b0))) begin
        start_write = 1'b1;
    end else begin
        start_write = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln77_fu_134_p2 = (k_1 + 16'd1);

assign add_ln80_fu_147_p2 = (j_1 + 16'd1);

assign add_ln83_fu_160_p2 = (i_1 + 16'd1);

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

always @ (*) begin
    ap_block_state1 = ((real_start == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1));
end

assign ap_ready = internal_ap_ready;

assign icmp_ln78_fu_141_p2 = ((add_ln77_fu_134_p2 == 16'd32) ? 1'b1 : 1'b0);

assign icmp_ln81_fu_154_p2 = ((add_ln80_fu_147_p2 == 16'd28) ? 1'b1 : 1'b0);

assign icmp_ln84_fu_166_p2 = ((add_ln83_fu_160_p2 == 16'd28) ? 1'b1 : 1'b0);

assign indices_0_din = i_1;

assign indices_1_din = j_1;

assign indices_2_out1_din = trunc_ln76_fu_128_p1;

assign indices_2_out_din = trunc_ln76_fu_128_p1;

assign select_ln84_fu_172_p3 = ((icmp_ln84_fu_166_p2[0:0] == 1'b1) ? 16'd0 : add_ln83_fu_160_p2);

assign start_out = real_start;

assign trunc_ln76_fu_128_p1 = k_1[4:0];

endmodule //td_fused_top_tdf6_get_next_ijk
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf6_readFilters46 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        filter_data_address0,
        filter_data_ce0,
        filter_data_q0,
        indices_23_dout,
        indices_23_empty_n,
        indices_23_read,
        weight_vecs_0_0_0_address0,
        weight_vecs_0_0_0_ce0,
        weight_vecs_0_0_0_we0,
        weight_vecs_0_0_0_d0
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state6 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [11:0] filter_data_address0;
output   filter_data_ce0;
input  [15:0] filter_data_q0;
input  [4:0] indices_23_dout;
input   indices_23_empty_n;
output   indices_23_read;
output  [6:0] weight_vecs_0_0_0_address0;
output   weight_vecs_0_0_0_ce0;
output   weight_vecs_0_0_0_we0;
output  [15:0] weight_vecs_0_0_0_d0;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg filter_data_ce0;
reg indices_23_read;
reg weight_vecs_0_0_0_ce0;
reg weight_vecs_0_0_0_we0;

reg    ap_done_reg;
  reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    indices_23_blk_n;
reg   [7:0] kk_0_0_i_i_reg_93;
reg   [7:0] kk_0_0_i_i_reg_93_pp0_iter1_reg;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
wire    ap_block_state4_pp0_stage0_iter2;
wire    ap_block_state5_pp0_stage0_iter3;
wire    ap_block_pp0_stage0_11001;
reg   [7:0] kk_0_0_i_i_reg_93_pp0_iter2_reg;
wire   [11:0] tmp_fu_105_p3;
reg   [11:0] tmp_reg_144;
wire   [7:0] add_ln49_fu_113_p2;
reg   [7:0] add_ln49_reg_149;
reg    ap_enable_reg_pp0_iter0;
wire   [0:0] icmp_ln49_fu_119_p2;
reg   [0:0] icmp_ln49_reg_154;
reg   [0:0] icmp_ln49_reg_154_pp0_iter1_reg;
reg   [0:0] icmp_ln49_reg_154_pp0_iter2_reg;
reg    ap_block_state1;
wire    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_exit_iter0_state2;
reg    ap_enable_reg_pp0_iter1;
reg    ap_enable_reg_pp0_iter2;
reg    ap_enable_reg_pp0_iter3;
reg   [7:0] ap_phi_mux_kk_0_0_i_i_phi_fu_97_p4;
wire    ap_block_pp0_stage0;
wire   [63:0] zext_ln55_20_fu_134_p1;
wire   [63:0] idxprom16_0_0_i_i_fu_139_p1;
wire   [11:0] zext_ln55_fu_125_p1;
wire   [11:0] add_ln55_fu_129_p2;
wire    ap_CS_fsm_state6;
reg   [2:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state6)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_condition_pp0_exit_iter0_state2) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            if ((1'b1 == ap_condition_pp0_exit_iter0_state2)) begin
                ap_enable_reg_pp0_iter1 <= (1'b1 ^ ap_condition_pp0_exit_iter0_state2);
            end else if ((1'b1 == 1'b1)) begin
                ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
            end
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end else if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter3 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln49_reg_154 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        kk_0_0_i_i_reg_93 <= add_ln49_reg_149;
    end else if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        kk_0_0_i_i_reg_93 <= 8'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        add_ln49_reg_149 <= add_ln49_fu_113_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln49_reg_154 <= icmp_ln49_fu_119_p2;
        icmp_ln49_reg_154_pp0_iter1_reg <= icmp_ln49_reg_154;
        kk_0_0_i_i_reg_93_pp0_iter1_reg <= kk_0_0_i_i_reg_93;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        icmp_ln49_reg_154_pp0_iter2_reg <= icmp_ln49_reg_154_pp0_iter1_reg;
        kk_0_0_i_i_reg_93_pp0_iter2_reg <= kk_0_0_i_i_reg_93_pp0_iter1_reg;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state1)) begin
        tmp_reg_144[11 : 7] <= tmp_fu_105_p3[11 : 7];
    end
end

always @ (*) begin
    if ((icmp_ln49_fu_119_p2 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state2 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state2 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state6)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln49_reg_154 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_kk_0_0_i_i_phi_fu_97_p4 = add_ln49_reg_149;
    end else begin
        ap_phi_mux_kk_0_0_i_i_phi_fu_97_p4 = kk_0_0_i_i_reg_93;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state6)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter3 == 1'b1)))) begin
        filter_data_ce0 = 1'b1;
    end else begin
        filter_data_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_23_blk_n = indices_23_empty_n;
    end else begin
        indices_23_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_23_read = 1'b1;
    end else begin
        indices_23_read = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter3 == 1'b1))) begin
        weight_vecs_0_0_0_ce0 = 1'b1;
    end else begin
        weight_vecs_0_0_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln49_reg_154_pp0_iter2_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter3 == 1'b1))) begin
        weight_vecs_0_0_0_we0 = 1'b1;
    end else begin
        weight_vecs_0_0_0_we0 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((~((icmp_ln49_fu_119_p2 == 1'd1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter1 == 1'b0)) & ~((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter3 == 1'b1) & (ap_enable_reg_pp0_iter2 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if ((((icmp_ln49_fu_119_p2 == 1'd1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter1 == 1'b0)) | ((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter3 == 1'b1) & (ap_enable_reg_pp0_iter2 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_state6;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state6 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln49_fu_113_p2 = (ap_phi_mux_kk_0_0_i_i_phi_fu_97_p4 + 8'd1);

assign add_ln55_fu_129_p2 = (tmp_reg_144 + zext_ln55_fu_125_p1);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state6 = ap_CS_fsm[32'd2];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1));
end

assign ap_block_state2_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign filter_data_address0 = zext_ln55_20_fu_134_p1;

assign icmp_ln49_fu_119_p2 = ((ap_phi_mux_kk_0_0_i_i_phi_fu_97_p4 == 8'd128) ? 1'b1 : 1'b0);

assign idxprom16_0_0_i_i_fu_139_p1 = kk_0_0_i_i_reg_93_pp0_iter2_reg;

assign tmp_fu_105_p3 = {{indices_23_dout}, {7'd0}};

assign weight_vecs_0_0_0_address0 = idxprom16_0_0_i_i_fu_139_p1;

assign weight_vecs_0_0_0_d0 = filter_data_q0;

assign zext_ln55_20_fu_134_p1 = add_ln55_fu_129_p2;

assign zext_ln55_fu_125_p1 = ap_phi_mux_kk_0_0_i_i_phi_fu_97_p4;

always @ (posedge ap_clk) begin
    tmp_reg_144[6:0] <= 7'b0000000;
end

endmodule //td_fused_top_tdf6_readFilters46
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf6_readInputs (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        in_data_address0,
        in_data_ce0,
        in_data_q0,
        indices_01_dout,
        indices_01_empty_n,
        indices_01_read,
        indices_12_dout,
        indices_12_empty_n,
        indices_12_read,
        ifmap_vec_0_0_address0,
        ifmap_vec_0_0_ce0,
        ifmap_vec_0_0_we0,
        ifmap_vec_0_0_d0,
        ifmap_vec_0_0_address1,
        ifmap_vec_0_0_ce1,
        ifmap_vec_0_0_we1,
        ifmap_vec_0_0_d1,
        indices_01_out_din,
        indices_01_out_full_n,
        indices_01_out_write,
        indices_12_out_din,
        indices_12_out_full_n,
        indices_12_out_write
);

parameter    ap_ST_fsm_state1 = 5'd1;
parameter    ap_ST_fsm_state2 = 5'd2;
parameter    ap_ST_fsm_pp0_stage0 = 5'd4;
parameter    ap_ST_fsm_pp0_stage1 = 5'd8;
parameter    ap_ST_fsm_state8 = 5'd16;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [14:0] in_data_address0;
output   in_data_ce0;
input  [63:0] in_data_q0;
input  [15:0] indices_01_dout;
input   indices_01_empty_n;
output   indices_01_read;
input  [15:0] indices_12_dout;
input   indices_12_empty_n;
output   indices_12_read;
output  [6:0] ifmap_vec_0_0_address0;
output   ifmap_vec_0_0_ce0;
output   ifmap_vec_0_0_we0;
output  [15:0] ifmap_vec_0_0_d0;
output  [6:0] ifmap_vec_0_0_address1;
output   ifmap_vec_0_0_ce1;
output   ifmap_vec_0_0_we1;
output  [15:0] ifmap_vec_0_0_d1;
output  [4:0] indices_01_out_din;
input   indices_01_out_full_n;
output   indices_01_out_write;
output  [9:0] indices_12_out_din;
input   indices_12_out_full_n;
output   indices_12_out_write;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg in_data_ce0;
reg indices_01_read;
reg indices_12_read;
reg[6:0] ifmap_vec_0_0_address0;
reg ifmap_vec_0_0_ce0;
reg ifmap_vec_0_0_we0;
reg[15:0] ifmap_vec_0_0_d0;
reg[6:0] ifmap_vec_0_0_address1;
reg ifmap_vec_0_0_ce1;
reg ifmap_vec_0_0_we1;
reg[15:0] ifmap_vec_0_0_d1;
reg indices_01_out_write;
reg indices_12_out_write;

reg    ap_done_reg;
  reg   [4:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    indices_01_blk_n;
reg    indices_12_blk_n;
reg    indices_01_out_blk_n;
reg    indices_12_out_blk_n;
reg   [7:0] kk_0_i_i_reg_180;
reg   [7:0] kk_0_i_i_reg_180_pp0_iter1_reg;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_block_state3_pp0_stage0_iter0;
wire    ap_block_state5_pp0_stage0_iter1;
wire    ap_block_state7_pp0_stage0_iter2;
wire    ap_block_pp0_stage0_11001;
wire   [4:0] trunc_ln135_fu_192_p1;
reg   [4:0] trunc_ln135_reg_434;
reg   [15:0] col_coord_reg_439;
wire   [0:0] is_padding_fu_214_p2;
reg   [0:0] is_padding_reg_444;
wire   [11:0] add_ln32_fu_274_p2;
reg   [11:0] add_ln32_reg_454;
wire    ap_CS_fsm_state2;
wire   [0:0] icmp_ln25_fu_280_p2;
reg   [0:0] icmp_ln25_reg_459;
reg   [0:0] icmp_ln25_reg_459_pp0_iter1_reg;
wire   [7:0] add_ln25_fu_308_p2;
reg   [7:0] add_ln25_reg_468;
wire    ap_CS_fsm_pp0_stage1;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_state4_pp0_stage1_iter0;
wire    ap_block_state6_pp0_stage1_iter1;
wire    ap_block_pp0_stage1_11001;
wire   [6:0] empty_80_fu_314_p1;
reg   [6:0] empty_80_reg_473;
wire   [15:0] select_ln33_11_fu_386_p3;
reg   [15:0] select_ln33_11_reg_479;
wire   [15:0] select_ln33_12_fu_407_p3;
reg   [15:0] select_ln33_12_reg_484;
wire    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_exit_iter0_state3;
reg    ap_enable_reg_pp0_iter1;
wire    ap_block_pp0_stage1_subdone;
reg    ap_enable_reg_pp0_iter2;
reg   [7:0] ap_phi_mux_kk_0_i_i_phi_fu_184_p4;
wire    ap_block_pp0_stage0;
wire   [63:0] sext_ln32_fu_303_p1;
wire   [63:0] zext_ln32_fu_318_p1;
wire    ap_block_pp0_stage1;
wire   [63:0] zext_ln32_10_fu_345_p1;
wire   [63:0] zext_ln32_11_fu_419_p1;
wire   [63:0] zext_ln32_12_fu_429_p1;
reg    ap_block_state1;
wire   [15:0] select_ln33_fu_331_p3;
wire   [15:0] select_ln33_10_fu_364_p3;
wire   [0:0] cmp7_i_i_fu_202_p2;
wire   [0:0] icmp_ln24_fu_208_p2;
wire   [4:0] empty_78_fu_220_p1;
wire   [4:0] row_coord_int_fu_223_p3;
wire   [9:0] tmp_fu_236_p3;
wire   [6:0] tmp_s_fu_248_p3;
wire   [10:0] zext_ln32_13_fu_244_p1;
wire   [10:0] zext_ln32_14_fu_256_p1;
wire   [10:0] sub_ln32_fu_260_p2;
wire   [4:0] col_coord_int_fu_229_p3;
wire   [11:0] sub_ln32_cast_fu_266_p1;
wire   [11:0] zext_ln32_15_fu_270_p1;
wire   [4:0] lshr_ln_fu_286_p4;
wire   [16:0] tmp_18_fu_296_p3;
wire   [15:0] trunc_ln32_fu_323_p1;
wire   [15:0] bitcast_ln32_fu_327_p1;
wire   [6:0] or_ln25_fu_339_p2;
wire   [15:0] tmp_31_i_i_fu_350_p4;
wire   [15:0] bitcast_ln32_10_fu_360_p1;
wire   [15:0] tmp_32_i_i_fu_372_p4;
wire   [15:0] bitcast_ln32_11_fu_382_p1;
wire   [15:0] tmp_33_i_i_fu_393_p4;
wire   [15:0] bitcast_ln32_12_fu_403_p1;
wire   [6:0] or_ln25_7_fu_414_p2;
wire   [6:0] or_ln25_8_fu_424_p2;
wire    ap_CS_fsm_state8;
reg   [4:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 5'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b1 == ap_condition_pp0_exit_iter0_state3))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1)) | ((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b0)))) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            ap_enable_reg_pp0_iter2 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln25_reg_459 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        kk_0_i_i_reg_180 <= add_ln25_reg_468;
    end else if ((1'b1 == ap_CS_fsm_state2)) begin
        kk_0_i_i_reg_180 <= 8'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln25_reg_459 == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
        add_ln25_reg_468 <= add_ln25_fu_308_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        add_ln32_reg_454 <= add_ln32_fu_274_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state1)) begin
        col_coord_reg_439 <= indices_12_dout;
        is_padding_reg_444 <= is_padding_fu_214_p2;
        trunc_ln135_reg_434 <= trunc_ln135_fu_192_p1;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln25_reg_459_pp0_iter1_reg == 1'd0))) begin
        empty_80_reg_473 <= empty_80_fu_314_p1;
        select_ln33_11_reg_479 <= select_ln33_11_fu_386_p3;
        select_ln33_12_reg_484 <= select_ln33_12_fu_407_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln25_reg_459 <= icmp_ln25_fu_280_p2;
        icmp_ln25_reg_459_pp0_iter1_reg <= icmp_ln25_reg_459;
        kk_0_i_i_reg_180_pp0_iter1_reg <= kk_0_i_i_reg_180;
    end
end

always @ (*) begin
    if ((icmp_ln25_fu_280_p2 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state3 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state3 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state8)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln25_reg_459 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_kk_0_i_i_phi_fu_184_p4 = add_ln25_reg_468;
    end else begin
        ap_phi_mux_kk_0_i_i_phi_fu_184_p4 = kk_0_i_i_reg_180;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state8)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        ifmap_vec_0_0_address0 = zext_ln32_12_fu_429_p1;
    end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ifmap_vec_0_0_address0 = zext_ln32_10_fu_345_p1;
    end else begin
        ifmap_vec_0_0_address0 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        ifmap_vec_0_0_address1 = zext_ln32_11_fu_419_p1;
    end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ifmap_vec_0_0_address1 = zext_ln32_fu_318_p1;
    end else begin
        ifmap_vec_0_0_address1 = 'bx;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1)) | ((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1)))) begin
        ifmap_vec_0_0_ce0 = 1'b1;
    end else begin
        ifmap_vec_0_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1)) | ((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1)))) begin
        ifmap_vec_0_0_ce1 = 1'b1;
    end else begin
        ifmap_vec_0_0_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        ifmap_vec_0_0_d0 = select_ln33_12_reg_484;
    end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ifmap_vec_0_0_d0 = select_ln33_10_fu_364_p3;
    end else begin
        ifmap_vec_0_0_d0 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        ifmap_vec_0_0_d1 = select_ln33_11_reg_479;
    end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ifmap_vec_0_0_d1 = select_ln33_fu_331_p3;
    end else begin
        ifmap_vec_0_0_d1 = 'bx;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1) & (icmp_ln25_reg_459_pp0_iter1_reg == 1'd0)) | ((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln25_reg_459_pp0_iter1_reg == 1'd0)))) begin
        ifmap_vec_0_0_we0 = 1'b1;
    end else begin
        ifmap_vec_0_0_we0 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1) & (icmp_ln25_reg_459_pp0_iter1_reg == 1'd0)) | ((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln25_reg_459_pp0_iter1_reg == 1'd0)))) begin
        ifmap_vec_0_0_we1 = 1'b1;
    end else begin
        ifmap_vec_0_0_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1)) | ((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1)) | ((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1)) | ((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1)))) begin
        in_data_ce0 = 1'b1;
    end else begin
        in_data_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_01_blk_n = indices_01_empty_n;
    end else begin
        indices_01_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_01_out_blk_n = indices_01_out_full_n;
    end else begin
        indices_01_out_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((indices_12_out_full_n == 1'b0) | (indices_01_out_full_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_01_out_write = 1'b1;
    end else begin
        indices_01_out_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((indices_12_out_full_n == 1'b0) | (indices_01_out_full_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_01_read = 1'b1;
    end else begin
        indices_01_read = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_12_blk_n = indices_12_empty_n;
    end else begin
        indices_12_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_12_out_blk_n = indices_12_out_full_n;
    end else begin
        indices_12_out_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((indices_12_out_full_n == 1'b0) | (indices_01_out_full_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_12_out_write = 1'b1;
    end else begin
        indices_12_out_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((indices_12_out_full_n == 1'b0) | (indices_01_out_full_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_12_read = 1'b1;
    end else begin
        indices_12_read = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((indices_12_out_full_n == 1'b0) | (indices_01_out_full_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_state2 : begin
            ap_NS_fsm = ap_ST_fsm_pp0_stage0;
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((~((icmp_ln25_fu_280_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1)) & ~((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0)) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end else if ((((icmp_ln25_fu_280_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1)) | ((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_state8;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_pp0_stage1 : begin
            if ((1'b0 == ap_block_pp0_stage1_subdone)) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end
        end
        ap_ST_fsm_state8 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln25_fu_308_p2 = (kk_0_i_i_reg_180 + 8'd4);

assign add_ln32_fu_274_p2 = ((sub_ln32_cast_fu_266_p1) + (zext_ln32_15_fu_270_p1));

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_pp0_stage1 = ap_CS_fsm[32'd3];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state8 = ap_CS_fsm[32'd4];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((indices_12_out_full_n == 1'b0) | (indices_01_out_full_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0));
end

assign ap_block_state3_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage1_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage1_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign bitcast_ln32_10_fu_360_p1 = tmp_31_i_i_fu_350_p4;

assign bitcast_ln32_11_fu_382_p1 = tmp_32_i_i_fu_372_p4;

assign bitcast_ln32_12_fu_403_p1 = tmp_33_i_i_fu_393_p4;

assign bitcast_ln32_fu_327_p1 = trunc_ln32_fu_323_p1;

assign cmp7_i_i_fu_202_p2 = ((indices_01_dout > 16'd27) ? 1'b1 : 1'b0);

assign col_coord_int_fu_229_p3 = ((is_padding_reg_444[0:0] == 1'b1) ? 5'd0 : empty_78_fu_220_p1);

assign empty_78_fu_220_p1 = col_coord_reg_439[4:0];

assign empty_80_fu_314_p1 = kk_0_i_i_reg_180_pp0_iter1_reg[6:0];

assign icmp_ln24_fu_208_p2 = ((indices_12_dout > 16'd27) ? 1'b1 : 1'b0);

assign icmp_ln25_fu_280_p2 = ((ap_phi_mux_kk_0_i_i_phi_fu_184_p4 == 8'd128) ? 1'b1 : 1'b0);

assign in_data_address0 = sext_ln32_fu_303_p1;

assign indices_01_out_din = indices_01_dout[4:0];

assign indices_12_out_din = indices_12_dout[9:0];

assign is_padding_fu_214_p2 = (icmp_ln24_fu_208_p2 | cmp7_i_i_fu_202_p2);

assign lshr_ln_fu_286_p4 = {{ap_phi_mux_kk_0_i_i_phi_fu_184_p4[6:2]}};

assign or_ln25_7_fu_414_p2 = (empty_80_reg_473 | 7'd2);

assign or_ln25_8_fu_424_p2 = (empty_80_reg_473 | 7'd3);

assign or_ln25_fu_339_p2 = (empty_80_fu_314_p1 | 7'd1);

assign row_coord_int_fu_223_p3 = ((is_padding_reg_444[0:0] == 1'b1) ? 5'd0 : trunc_ln135_reg_434);

assign select_ln33_10_fu_364_p3 = ((is_padding_reg_444[0:0] == 1'b1) ? 16'd0 : bitcast_ln32_10_fu_360_p1);

assign select_ln33_11_fu_386_p3 = ((is_padding_reg_444[0:0] == 1'b1) ? 16'd0 : bitcast_ln32_11_fu_382_p1);

assign select_ln33_12_fu_407_p3 = ((is_padding_reg_444[0:0] == 1'b1) ? 16'd0 : bitcast_ln32_12_fu_403_p1);

assign select_ln33_fu_331_p3 = ((is_padding_reg_444[0:0] == 1'b1) ? 16'd0 : bitcast_ln32_fu_327_p1);

assign sext_ln32_fu_303_p1 = (tmp_18_fu_296_p3);

assign sub_ln32_cast_fu_266_p1 = (sub_ln32_fu_260_p2);

assign sub_ln32_fu_260_p2 = (zext_ln32_13_fu_244_p1 - zext_ln32_14_fu_256_p1);

assign tmp_18_fu_296_p3 = {{add_ln32_reg_454}, {lshr_ln_fu_286_p4}};

assign tmp_31_i_i_fu_350_p4 = {{in_data_q0[31:16]}};

assign tmp_32_i_i_fu_372_p4 = {{in_data_q0[47:32]}};

assign tmp_33_i_i_fu_393_p4 = {{in_data_q0[63:48]}};

assign tmp_fu_236_p3 = {{row_coord_int_fu_223_p3}, {5'd0}};

assign tmp_s_fu_248_p3 = {{row_coord_int_fu_223_p3}, {2'd0}};

assign trunc_ln135_fu_192_p1 = indices_01_dout[4:0];

assign trunc_ln32_fu_323_p1 = in_data_q0[15:0];

assign zext_ln32_10_fu_345_p1 = or_ln25_fu_339_p2;

assign zext_ln32_11_fu_419_p1 = or_ln25_7_fu_414_p2;

assign zext_ln32_12_fu_429_p1 = or_ln25_8_fu_424_p2;

assign zext_ln32_13_fu_244_p1 = tmp_fu_236_p3;

assign zext_ln32_14_fu_256_p1 = tmp_s_fu_248_p3;

assign zext_ln32_15_fu_270_p1 = col_coord_int_fu_229_p3;

assign zext_ln32_fu_318_p1 = kk_0_i_i_reg_180_pp0_iter1_reg;

endmodule //td_fused_top_tdf6_readInputs
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf6_writeOutputs_unaligned (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        indices_01_dout,
        indices_01_empty_n,
        indices_01_read,
        indices_12_dout,
        indices_12_empty_n,
        indices_12_read,
        p_read,
        out_data_address1,
        out_data_ce1,
        out_data_we1,
        out_data_d1
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_state2 = 3'd2;
parameter    ap_ST_fsm_state3 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
input  [4:0] indices_01_dout;
input   indices_01_empty_n;
output   indices_01_read;
input  [9:0] indices_12_dout;
input   indices_12_empty_n;
output   indices_12_read;
input  [15:0] p_read;
output  [12:0] out_data_address1;
output   out_data_ce1;
output   out_data_we1;
output  [63:0] out_data_d1;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg indices_01_read;
reg indices_12_read;
reg out_data_ce1;
reg out_data_we1;

reg    ap_done_reg;
  reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg   [15:0] outputCount_4;
reg   [15:0] outputChanIdx_4;
reg   [15:0] outputRow_12_0;
reg   [15:0] outputRow_12_1;
reg   [15:0] outputRow_12_2;
reg   [15:0] outputRow_12_3;
reg    indices_01_blk_n;
reg    indices_12_blk_n;
wire   [9:0] add_ln94_fu_147_p2;
reg   [9:0] add_ln94_reg_304;
wire   [15:0] add_ln87_fu_192_p2;
wire    ap_CS_fsm_state2;
wire   [0:0] icmp_ln88_fu_198_p2;
reg   [0:0] icmp_ln88_reg_317;
reg   [15:0] ap_phi_mux_empty_phi_fu_114_p4;
reg   [15:0] empty_reg_111;
wire    ap_CS_fsm_state3;
wire   [63:0] zext_ln94_6_fu_226_p1;
wire   [15:0] select_ln97_fu_284_p3;
wire   [1:0] trunc_ln86_fu_164_p1;
reg   [15:0] ap_sig_allocacmp_outputRow_12_0_load;
reg   [15:0] ap_sig_allocacmp_outputRow_12_1_load;
reg   [15:0] ap_sig_allocacmp_outputRow_12_2_load;
reg   [15:0] ap_sig_allocacmp_outputRow_12_3_load;
reg    ap_block_state1;
wire   [6:0] tmp_s_fu_129_p3;
wire   [9:0] tmp_fu_121_p3;
wire   [9:0] zext_ln94_fu_137_p1;
wire   [9:0] sub_ln94_fu_141_p2;
wire   [4:0] trunc_ln94_fu_212_p1;
wire   [12:0] tmp_53_cast_fu_153_p3;
wire   [12:0] zext_ln94_5_fu_216_p1;
wire   [12:0] add_ln94_3_fu_220_p2;
wire   [15:0] bitcast_ln94_9_fu_255_p1;
wire   [15:0] bitcast_ln94_8_fu_247_p1;
wire   [15:0] bitcast_ln94_7_fu_239_p1;
wire   [15:0] bitcast_ln94_fu_231_p1;
wire   [15:0] add_ln96_fu_272_p2;
wire   [0:0] icmp_ln97_fu_278_p2;
reg   [2:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 3'd1;
#0 outputCount_4 = 16'd0;
#0 outputChanIdx_4 = 16'd0;
#0 outputRow_12_0 = 16'd0;
#0 outputRow_12_1 = 16'd0;
#0 outputRow_12_2 = 16'd0;
#0 outputRow_12_3 = 16'd0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state3)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln88_reg_317 == 1'd1) & (1'b1 == ap_CS_fsm_state3))) begin
        empty_reg_111 <= 16'd0;
    end else if (((icmp_ln88_fu_198_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state2))) begin
        empty_reg_111 <= add_ln87_fu_192_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state1)) begin
        add_ln94_reg_304 <= add_ln94_fu_147_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        icmp_ln88_reg_317 <= icmp_ln88_fu_198_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln88_fu_198_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        outputChanIdx_4 <= select_ln97_fu_284_p3;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state3)) begin
        outputCount_4 <= ap_phi_mux_empty_phi_fu_114_p4;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln86_fu_164_p1 == 2'd0) & (1'b1 == ap_CS_fsm_state2))) begin
        outputRow_12_0 <= p_read;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln86_fu_164_p1 == 2'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        outputRow_12_1 <= p_read;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln86_fu_164_p1 == 2'd2) & (1'b1 == ap_CS_fsm_state2))) begin
        outputRow_12_2 <= p_read;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln86_fu_164_p1 == 2'd3) & (1'b1 == ap_CS_fsm_state2))) begin
        outputRow_12_3 <= p_read;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state3)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln88_reg_317 == 1'd1) & (1'b1 == ap_CS_fsm_state3))) begin
        ap_phi_mux_empty_phi_fu_114_p4 = 16'd0;
    end else begin
        ap_phi_mux_empty_phi_fu_114_p4 = empty_reg_111;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state3)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((trunc_ln86_fu_164_p1 == 2'd0) & (1'b1 == ap_CS_fsm_state2))) begin
        ap_sig_allocacmp_outputRow_12_0_load = p_read;
    end else begin
        ap_sig_allocacmp_outputRow_12_0_load = outputRow_12_0;
    end
end

always @ (*) begin
    if (((trunc_ln86_fu_164_p1 == 2'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        ap_sig_allocacmp_outputRow_12_1_load = p_read;
    end else begin
        ap_sig_allocacmp_outputRow_12_1_load = outputRow_12_1;
    end
end

always @ (*) begin
    if (((trunc_ln86_fu_164_p1 == 2'd2) & (1'b1 == ap_CS_fsm_state2))) begin
        ap_sig_allocacmp_outputRow_12_2_load = p_read;
    end else begin
        ap_sig_allocacmp_outputRow_12_2_load = outputRow_12_2;
    end
end

always @ (*) begin
    if (((trunc_ln86_fu_164_p1 == 2'd3) & (1'b1 == ap_CS_fsm_state2))) begin
        ap_sig_allocacmp_outputRow_12_3_load = p_read;
    end else begin
        ap_sig_allocacmp_outputRow_12_3_load = outputRow_12_3;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_01_blk_n = indices_01_empty_n;
    end else begin
        indices_01_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_01_read = 1'b1;
    end else begin
        indices_01_read = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_12_blk_n = indices_12_empty_n;
    end else begin
        indices_12_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_12_read = 1'b1;
    end else begin
        indices_12_read = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state2))) begin
        out_data_ce1 = 1'b1;
    end else begin
        out_data_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln88_fu_198_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        out_data_we1 = 1'b1;
    end else begin
        out_data_we1 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_start == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_state2 : begin
            ap_NS_fsm = ap_ST_fsm_state3;
        end
        ap_ST_fsm_state3 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln87_fu_192_p2 = (outputCount_4 + 16'd1);

assign add_ln94_3_fu_220_p2 = (tmp_53_cast_fu_153_p3 + zext_ln94_5_fu_216_p1);

assign add_ln94_fu_147_p2 = (sub_ln94_fu_141_p2 + indices_12_dout);

assign add_ln96_fu_272_p2 = (outputChanIdx_4 + 16'd1);

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1));
end

assign bitcast_ln94_7_fu_239_p1 = ap_sig_allocacmp_outputRow_12_1_load;

assign bitcast_ln94_8_fu_247_p1 = ap_sig_allocacmp_outputRow_12_2_load;

assign bitcast_ln94_9_fu_255_p1 = ap_sig_allocacmp_outputRow_12_3_load;

assign bitcast_ln94_fu_231_p1 = ap_sig_allocacmp_outputRow_12_0_load;

assign icmp_ln88_fu_198_p2 = ((add_ln87_fu_192_p2 == 16'd4) ? 1'b1 : 1'b0);

assign icmp_ln97_fu_278_p2 = ((add_ln96_fu_272_p2 == 16'd8) ? 1'b1 : 1'b0);

assign out_data_address1 = zext_ln94_6_fu_226_p1;

assign out_data_d1 = {{{{bitcast_ln94_9_fu_255_p1}, {bitcast_ln94_8_fu_247_p1}}, {bitcast_ln94_7_fu_239_p1}}, {bitcast_ln94_fu_231_p1}};

assign select_ln97_fu_284_p3 = ((icmp_ln97_fu_278_p2[0:0] == 1'b1) ? 16'd0 : add_ln96_fu_272_p2);

assign sub_ln94_fu_141_p2 = (tmp_fu_121_p3 - zext_ln94_fu_137_p1);

assign tmp_53_cast_fu_153_p3 = {{add_ln94_reg_304}, {3'd0}};

assign tmp_fu_121_p3 = {{indices_01_dout}, {5'd0}};

assign tmp_s_fu_129_p3 = {{indices_01_dout}, {2'd0}};

assign trunc_ln86_fu_164_p1 = outputCount_4[1:0];

assign trunc_ln94_fu_212_p1 = outputChanIdx_4[4:0];

assign zext_ln94_5_fu_216_p1 = trunc_ln94_fu_212_p1;

assign zext_ln94_6_fu_226_p1 = add_ln94_3_fu_220_p2;

assign zext_ln94_fu_137_p1 = tmp_s_fu_129_p3;

endmodule //td_fused_top_tdf6_writeOutputs_unaligned
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf7_18 (
        in_data_address0,
        in_data_ce0,
        in_data_d0,
        in_data_q0,
        in_data_we0,
        in_data_address1,
        in_data_ce1,
        in_data_d1,
        in_data_q1,
        in_data_we1,
        out_data_address0,
        out_data_ce0,
        out_data_d0,
        out_data_q0,
        out_data_we0,
        out_data_address1,
        out_data_ce1,
        out_data_d1,
        out_data_q1,
        out_data_we1,
        l1_filter_data_address0,
        l1_filter_data_ce0,
        l1_filter_data_d0,
        l1_filter_data_q0,
        l1_filter_data_we0,
        l1_filter_data_address1,
        l1_filter_data_ce1,
        l1_filter_data_d1,
        l1_filter_data_q1,
        l1_filter_data_we1,
        l2_filter_data_address0,
        l2_filter_data_ce0,
        l2_filter_data_d0,
        l2_filter_data_q0,
        l2_filter_data_we0,
        l2_filter_data_address1,
        l2_filter_data_ce1,
        l2_filter_data_d1,
        l2_filter_data_q1,
        l2_filter_data_we1,
        l1_adjustments_address0,
        l1_adjustments_ce0,
        l1_adjustments_d0,
        l1_adjustments_q0,
        l1_adjustments_we0,
        l1_adjustments_address1,
        l1_adjustments_ce1,
        l1_adjustments_d1,
        l1_adjustments_q1,
        l1_adjustments_we1,
        l2_adjustments_address0,
        l2_adjustments_ce0,
        l2_adjustments_d0,
        l2_adjustments_q0,
        l2_adjustments_we0,
        l2_adjustments_address1,
        l2_adjustments_ce1,
        l2_adjustments_d1,
        l2_adjustments_q1,
        l2_adjustments_we1,
        ap_clk,
        ap_rst,
        in_data_empty_n,
        in_data_read,
        out_data_full_n,
        out_data_write,
        ap_start,
        ap_done,
        ap_ready,
        ap_idle,
        ap_continue
);


output  [12:0] in_data_address0;
output   in_data_ce0;
output  [63:0] in_data_d0;
input  [63:0] in_data_q0;
output   in_data_we0;
output  [12:0] in_data_address1;
output   in_data_ce1;
output  [63:0] in_data_d1;
input  [63:0] in_data_q1;
output   in_data_we1;
output  [12:0] out_data_address0;
output   out_data_ce0;
output  [63:0] out_data_d0;
input  [63:0] out_data_q0;
output   out_data_we0;
output  [12:0] out_data_address1;
output   out_data_ce1;
output  [63:0] out_data_d1;
input  [63:0] out_data_q1;
output   out_data_we1;
output  [16:0] l1_filter_data_address0;
output   l1_filter_data_ce0;
output  [15:0] l1_filter_data_d0;
input  [15:0] l1_filter_data_q0;
output   l1_filter_data_we0;
output  [16:0] l1_filter_data_address1;
output   l1_filter_data_ce1;
output  [15:0] l1_filter_data_d1;
input  [15:0] l1_filter_data_q1;
output   l1_filter_data_we1;
output  [12:0] l2_filter_data_address0;
output   l2_filter_data_ce0;
output  [15:0] l2_filter_data_d0;
input  [15:0] l2_filter_data_q0;
output   l2_filter_data_we0;
output  [12:0] l2_filter_data_address1;
output   l2_filter_data_ce1;
output  [15:0] l2_filter_data_d1;
input  [15:0] l2_filter_data_q1;
output   l2_filter_data_we1;
output  [7:0] l1_adjustments_address0;
output   l1_adjustments_ce0;
output  [47:0] l1_adjustments_d0;
input  [47:0] l1_adjustments_q0;
output   l1_adjustments_we0;
output  [7:0] l1_adjustments_address1;
output   l1_adjustments_ce1;
output  [47:0] l1_adjustments_d1;
input  [47:0] l1_adjustments_q1;
output   l1_adjustments_we1;
output  [4:0] l2_adjustments_address0;
output   l2_adjustments_ce0;
output  [47:0] l2_adjustments_d0;
input  [47:0] l2_adjustments_q0;
output   l2_adjustments_we0;
output  [4:0] l2_adjustments_address1;
output   l2_adjustments_ce1;
output  [47:0] l2_adjustments_d1;
input  [47:0] l2_adjustments_q1;
output   l2_adjustments_we1;
input   ap_clk;
input   ap_rst;
input   in_data_empty_n;
output   in_data_read;
input   out_data_full_n;
output   out_data_write;
input   ap_start;
output   ap_done;
output   ap_ready;
output   ap_idle;
input   ap_continue;

reg ap_done;
reg ap_ready;
reg ap_idle;

wire   [12:0] dataflow_in_loop_TOP_LOOP37548_U0_in_data_address0;
wire    dataflow_in_loop_TOP_LOOP37548_U0_in_data_ce0;
wire   [63:0] dataflow_in_loop_TOP_LOOP37548_U0_in_data_d0;
wire    dataflow_in_loop_TOP_LOOP37548_U0_in_data_we0;
wire   [12:0] dataflow_in_loop_TOP_LOOP37548_U0_in_data_address1;
wire    dataflow_in_loop_TOP_LOOP37548_U0_in_data_ce1;
wire   [63:0] dataflow_in_loop_TOP_LOOP37548_U0_in_data_d1;
wire    dataflow_in_loop_TOP_LOOP37548_U0_in_data_we1;
wire   [16:0] dataflow_in_loop_TOP_LOOP37548_U0_l1_filter_data_address0;
wire    dataflow_in_loop_TOP_LOOP37548_U0_l1_filter_data_ce0;
wire   [15:0] dataflow_in_loop_TOP_LOOP37548_U0_l1_filter_data_d0;
wire    dataflow_in_loop_TOP_LOOP37548_U0_l1_filter_data_we0;
wire   [16:0] dataflow_in_loop_TOP_LOOP37548_U0_l1_filter_data_address1;
wire    dataflow_in_loop_TOP_LOOP37548_U0_l1_filter_data_ce1;
wire   [15:0] dataflow_in_loop_TOP_LOOP37548_U0_l1_filter_data_d1;
wire    dataflow_in_loop_TOP_LOOP37548_U0_l1_filter_data_we1;
wire   [7:0] dataflow_in_loop_TOP_LOOP37548_U0_l1_adjustments_address0;
wire    dataflow_in_loop_TOP_LOOP37548_U0_l1_adjustments_ce0;
wire   [47:0] dataflow_in_loop_TOP_LOOP37548_U0_l1_adjustments_d0;
wire    dataflow_in_loop_TOP_LOOP37548_U0_l1_adjustments_we0;
wire   [7:0] dataflow_in_loop_TOP_LOOP37548_U0_l1_adjustments_address1;
wire    dataflow_in_loop_TOP_LOOP37548_U0_l1_adjustments_ce1;
wire   [47:0] dataflow_in_loop_TOP_LOOP37548_U0_l1_adjustments_d1;
wire    dataflow_in_loop_TOP_LOOP37548_U0_l1_adjustments_we1;
wire   [12:0] dataflow_in_loop_TOP_LOOP37548_U0_l2_filter_data_address0;
wire    dataflow_in_loop_TOP_LOOP37548_U0_l2_filter_data_ce0;
wire   [15:0] dataflow_in_loop_TOP_LOOP37548_U0_l2_filter_data_d0;
wire    dataflow_in_loop_TOP_LOOP37548_U0_l2_filter_data_we0;
wire   [12:0] dataflow_in_loop_TOP_LOOP37548_U0_l2_filter_data_address1;
wire    dataflow_in_loop_TOP_LOOP37548_U0_l2_filter_data_ce1;
wire   [15:0] dataflow_in_loop_TOP_LOOP37548_U0_l2_filter_data_d1;
wire    dataflow_in_loop_TOP_LOOP37548_U0_l2_filter_data_we1;
wire   [12:0] dataflow_in_loop_TOP_LOOP37548_U0_out_data_address0;
wire    dataflow_in_loop_TOP_LOOP37548_U0_out_data_ce0;
wire   [63:0] dataflow_in_loop_TOP_LOOP37548_U0_out_data_d0;
wire    dataflow_in_loop_TOP_LOOP37548_U0_out_data_we0;
wire   [12:0] dataflow_in_loop_TOP_LOOP37548_U0_out_data_address1;
wire    dataflow_in_loop_TOP_LOOP37548_U0_out_data_ce1;
wire   [63:0] dataflow_in_loop_TOP_LOOP37548_U0_out_data_d1;
wire    dataflow_in_loop_TOP_LOOP37548_U0_out_data_we1;
wire   [4:0] dataflow_in_loop_TOP_LOOP37548_U0_l2_adjustments_address0;
wire    dataflow_in_loop_TOP_LOOP37548_U0_l2_adjustments_ce0;
wire   [47:0] dataflow_in_loop_TOP_LOOP37548_U0_l2_adjustments_d0;
wire    dataflow_in_loop_TOP_LOOP37548_U0_l2_adjustments_we0;
wire   [4:0] dataflow_in_loop_TOP_LOOP37548_U0_l2_adjustments_address1;
wire    dataflow_in_loop_TOP_LOOP37548_U0_l2_adjustments_ce1;
wire   [47:0] dataflow_in_loop_TOP_LOOP37548_U0_l2_adjustments_d1;
wire    dataflow_in_loop_TOP_LOOP37548_U0_l2_adjustments_we1;
wire    dataflow_in_loop_TOP_LOOP37548_U0_ap_start;
wire    dataflow_in_loop_TOP_LOOP37548_U0_in_data_read;
wire    dataflow_in_loop_TOP_LOOP37548_U0_out_data_write;
wire    dataflow_in_loop_TOP_LOOP37548_U0_ap_done;
wire    dataflow_in_loop_TOP_LOOP37548_U0_ap_ready;
wire    dataflow_in_loop_TOP_LOOP37548_U0_ap_idle;
reg    dataflow_in_loop_TOP_LOOP37548_U0_ap_continue;
wire    dataflow_in_loop_TOP_LOOP37548_U0_in_data_full_n;
wire    dataflow_in_loop_TOP_LOOP37548_U0_in_data_write;
wire    ap_sync_continue;
wire    ap_sync_done;
wire    ap_sync_ready;
reg   [17:0] loop_dataflow_input_count;
reg   [17:0] loop_dataflow_output_count;
wire   [17:0] bound_minus_1;
wire    dataflow_in_loop_TOP_LOOP37548_U0_start_full_n;
wire    dataflow_in_loop_TOP_LOOP37548_U0_start_write;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 loop_dataflow_input_count = 18'd0;
#0 loop_dataflow_output_count = 18'd0;
end

td_fused_top_dataflow_in_loop_TOP_LOOP37548 dataflow_in_loop_TOP_LOOP37548_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .in_data_address0(dataflow_in_loop_TOP_LOOP37548_U0_in_data_address0),
    .in_data_ce0(dataflow_in_loop_TOP_LOOP37548_U0_in_data_ce0),
    .in_data_d0(dataflow_in_loop_TOP_LOOP37548_U0_in_data_d0),
    .in_data_q0(in_data_q0),
    .in_data_we0(dataflow_in_loop_TOP_LOOP37548_U0_in_data_we0),
    .in_data_address1(dataflow_in_loop_TOP_LOOP37548_U0_in_data_address1),
    .in_data_ce1(dataflow_in_loop_TOP_LOOP37548_U0_in_data_ce1),
    .in_data_d1(dataflow_in_loop_TOP_LOOP37548_U0_in_data_d1),
    .in_data_q1(64'd0),
    .in_data_we1(dataflow_in_loop_TOP_LOOP37548_U0_in_data_we1),
    .l1_filter_data_address0(dataflow_in_loop_TOP_LOOP37548_U0_l1_filter_data_address0),
    .l1_filter_data_ce0(dataflow_in_loop_TOP_LOOP37548_U0_l1_filter_data_ce0),
    .l1_filter_data_d0(dataflow_in_loop_TOP_LOOP37548_U0_l1_filter_data_d0),
    .l1_filter_data_q0(l1_filter_data_q0),
    .l1_filter_data_we0(dataflow_in_loop_TOP_LOOP37548_U0_l1_filter_data_we0),
    .l1_filter_data_address1(dataflow_in_loop_TOP_LOOP37548_U0_l1_filter_data_address1),
    .l1_filter_data_ce1(dataflow_in_loop_TOP_LOOP37548_U0_l1_filter_data_ce1),
    .l1_filter_data_d1(dataflow_in_loop_TOP_LOOP37548_U0_l1_filter_data_d1),
    .l1_filter_data_q1(16'd0),
    .l1_filter_data_we1(dataflow_in_loop_TOP_LOOP37548_U0_l1_filter_data_we1),
    .l1_adjustments_address0(dataflow_in_loop_TOP_LOOP37548_U0_l1_adjustments_address0),
    .l1_adjustments_ce0(dataflow_in_loop_TOP_LOOP37548_U0_l1_adjustments_ce0),
    .l1_adjustments_d0(dataflow_in_loop_TOP_LOOP37548_U0_l1_adjustments_d0),
    .l1_adjustments_q0(l1_adjustments_q0),
    .l1_adjustments_we0(dataflow_in_loop_TOP_LOOP37548_U0_l1_adjustments_we0),
    .l1_adjustments_address1(dataflow_in_loop_TOP_LOOP37548_U0_l1_adjustments_address1),
    .l1_adjustments_ce1(dataflow_in_loop_TOP_LOOP37548_U0_l1_adjustments_ce1),
    .l1_adjustments_d1(dataflow_in_loop_TOP_LOOP37548_U0_l1_adjustments_d1),
    .l1_adjustments_q1(48'd0),
    .l1_adjustments_we1(dataflow_in_loop_TOP_LOOP37548_U0_l1_adjustments_we1),
    .l2_filter_data_address0(dataflow_in_loop_TOP_LOOP37548_U0_l2_filter_data_address0),
    .l2_filter_data_ce0(dataflow_in_loop_TOP_LOOP37548_U0_l2_filter_data_ce0),
    .l2_filter_data_d0(dataflow_in_loop_TOP_LOOP37548_U0_l2_filter_data_d0),
    .l2_filter_data_q0(l2_filter_data_q0),
    .l2_filter_data_we0(dataflow_in_loop_TOP_LOOP37548_U0_l2_filter_data_we0),
    .l2_filter_data_address1(dataflow_in_loop_TOP_LOOP37548_U0_l2_filter_data_address1),
    .l2_filter_data_ce1(dataflow_in_loop_TOP_LOOP37548_U0_l2_filter_data_ce1),
    .l2_filter_data_d1(dataflow_in_loop_TOP_LOOP37548_U0_l2_filter_data_d1),
    .l2_filter_data_q1(16'd0),
    .l2_filter_data_we1(dataflow_in_loop_TOP_LOOP37548_U0_l2_filter_data_we1),
    .out_data_address0(dataflow_in_loop_TOP_LOOP37548_U0_out_data_address0),
    .out_data_ce0(dataflow_in_loop_TOP_LOOP37548_U0_out_data_ce0),
    .out_data_d0(dataflow_in_loop_TOP_LOOP37548_U0_out_data_d0),
    .out_data_q0(64'd0),
    .out_data_we0(dataflow_in_loop_TOP_LOOP37548_U0_out_data_we0),
    .out_data_address1(dataflow_in_loop_TOP_LOOP37548_U0_out_data_address1),
    .out_data_ce1(dataflow_in_loop_TOP_LOOP37548_U0_out_data_ce1),
    .out_data_d1(dataflow_in_loop_TOP_LOOP37548_U0_out_data_d1),
    .out_data_q1(64'd0),
    .out_data_we1(dataflow_in_loop_TOP_LOOP37548_U0_out_data_we1),
    .l2_adjustments_address0(dataflow_in_loop_TOP_LOOP37548_U0_l2_adjustments_address0),
    .l2_adjustments_ce0(dataflow_in_loop_TOP_LOOP37548_U0_l2_adjustments_ce0),
    .l2_adjustments_d0(dataflow_in_loop_TOP_LOOP37548_U0_l2_adjustments_d0),
    .l2_adjustments_q0(l2_adjustments_q0),
    .l2_adjustments_we0(dataflow_in_loop_TOP_LOOP37548_U0_l2_adjustments_we0),
    .l2_adjustments_address1(dataflow_in_loop_TOP_LOOP37548_U0_l2_adjustments_address1),
    .l2_adjustments_ce1(dataflow_in_loop_TOP_LOOP37548_U0_l2_adjustments_ce1),
    .l2_adjustments_d1(dataflow_in_loop_TOP_LOOP37548_U0_l2_adjustments_d1),
    .l2_adjustments_q1(48'd0),
    .l2_adjustments_we1(dataflow_in_loop_TOP_LOOP37548_U0_l2_adjustments_we1),
    .ap_start(dataflow_in_loop_TOP_LOOP37548_U0_ap_start),
    .in_data_empty_n(1'b0),
    .in_data_read(dataflow_in_loop_TOP_LOOP37548_U0_in_data_read),
    .out_data_full_n(out_data_full_n),
    .out_data_write(dataflow_in_loop_TOP_LOOP37548_U0_out_data_write),
    .ap_done(dataflow_in_loop_TOP_LOOP37548_U0_ap_done),
    .ap_ready(dataflow_in_loop_TOP_LOOP37548_U0_ap_ready),
    .ap_idle(dataflow_in_loop_TOP_LOOP37548_U0_ap_idle),
    .ap_continue(dataflow_in_loop_TOP_LOOP37548_U0_ap_continue)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        loop_dataflow_input_count <= 18'd0;
    end else begin
        if ((~(loop_dataflow_input_count == bound_minus_1) & (ap_start == 1'b1) & (dataflow_in_loop_TOP_LOOP37548_U0_ap_ready == 1'b1))) begin
            loop_dataflow_input_count <= (loop_dataflow_input_count + 18'd1);
        end else if (((loop_dataflow_input_count == bound_minus_1) & (ap_start == 1'b1) & (dataflow_in_loop_TOP_LOOP37548_U0_ap_ready == 1'b1))) begin
            loop_dataflow_input_count <= 18'd0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        loop_dataflow_output_count <= 18'd0;
    end else begin
        if ((~(loop_dataflow_output_count == bound_minus_1) & (dataflow_in_loop_TOP_LOOP37548_U0_ap_continue == 1'b1) & (dataflow_in_loop_TOP_LOOP37548_U0_ap_done == 1'b1))) begin
            loop_dataflow_output_count <= (loop_dataflow_output_count + 18'd1);
        end else if (((loop_dataflow_output_count == bound_minus_1) & (dataflow_in_loop_TOP_LOOP37548_U0_ap_continue == 1'b1) & (dataflow_in_loop_TOP_LOOP37548_U0_ap_done == 1'b1))) begin
            loop_dataflow_output_count <= 18'd0;
        end
    end
end

always @ (*) begin
    if (((loop_dataflow_output_count == bound_minus_1) & (dataflow_in_loop_TOP_LOOP37548_U0_ap_done == 1'b1))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = 1'b0;
    end
end

always @ (*) begin
    if (((loop_dataflow_output_count == 18'd0) & (ap_start == 1'b0) & (dataflow_in_loop_TOP_LOOP37548_U0_ap_idle == 1'b1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((loop_dataflow_input_count == bound_minus_1) & (ap_start == 1'b1) & (dataflow_in_loop_TOP_LOOP37548_U0_ap_ready == 1'b1))) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((~(loop_dataflow_output_count == bound_minus_1) | (ap_continue == 1'b1))) begin
        dataflow_in_loop_TOP_LOOP37548_U0_ap_continue = 1'b1;
    end else begin
        dataflow_in_loop_TOP_LOOP37548_U0_ap_continue = 1'b0;
    end
end

assign ap_sync_continue = ap_continue;

assign ap_sync_done = dataflow_in_loop_TOP_LOOP37548_U0_ap_done;

assign ap_sync_ready = dataflow_in_loop_TOP_LOOP37548_U0_ap_ready;

assign bound_minus_1 = (18'd200704 - 18'd1);

assign dataflow_in_loop_TOP_LOOP37548_U0_ap_start = ap_start;

assign dataflow_in_loop_TOP_LOOP37548_U0_in_data_full_n = in_data_empty_n;

assign dataflow_in_loop_TOP_LOOP37548_U0_in_data_write = 1'b0;

assign dataflow_in_loop_TOP_LOOP37548_U0_start_full_n = 1'b1;

assign dataflow_in_loop_TOP_LOOP37548_U0_start_write = 1'b0;

assign in_data_address0 = dataflow_in_loop_TOP_LOOP37548_U0_in_data_address0;

assign in_data_address1 = 13'd0;

assign in_data_ce0 = dataflow_in_loop_TOP_LOOP37548_U0_in_data_ce0;

assign in_data_ce1 = 1'b0;

assign in_data_d0 = 64'd0;

assign in_data_d1 = 64'd0;

assign in_data_read = dataflow_in_loop_TOP_LOOP37548_U0_in_data_write;

assign in_data_we0 = 1'b0;

assign in_data_we1 = 1'b0;

assign l1_adjustments_address0 = dataflow_in_loop_TOP_LOOP37548_U0_l1_adjustments_address0;

assign l1_adjustments_address1 = 8'd0;

assign l1_adjustments_ce0 = dataflow_in_loop_TOP_LOOP37548_U0_l1_adjustments_ce0;

assign l1_adjustments_ce1 = 1'b0;

assign l1_adjustments_d0 = 48'd0;

assign l1_adjustments_d1 = 48'd0;

assign l1_adjustments_we0 = 1'b0;

assign l1_adjustments_we1 = 1'b0;

assign l1_filter_data_address0 = dataflow_in_loop_TOP_LOOP37548_U0_l1_filter_data_address0;

assign l1_filter_data_address1 = 17'd0;

assign l1_filter_data_ce0 = dataflow_in_loop_TOP_LOOP37548_U0_l1_filter_data_ce0;

assign l1_filter_data_ce1 = 1'b0;

assign l1_filter_data_d0 = 16'd0;

assign l1_filter_data_d1 = 16'd0;

assign l1_filter_data_we0 = 1'b0;

assign l1_filter_data_we1 = 1'b0;

assign l2_adjustments_address0 = dataflow_in_loop_TOP_LOOP37548_U0_l2_adjustments_address0;

assign l2_adjustments_address1 = 5'd0;

assign l2_adjustments_ce0 = dataflow_in_loop_TOP_LOOP37548_U0_l2_adjustments_ce0;

assign l2_adjustments_ce1 = 1'b0;

assign l2_adjustments_d0 = 48'd0;

assign l2_adjustments_d1 = 48'd0;

assign l2_adjustments_we0 = 1'b0;

assign l2_adjustments_we1 = 1'b0;

assign l2_filter_data_address0 = dataflow_in_loop_TOP_LOOP37548_U0_l2_filter_data_address0;

assign l2_filter_data_address1 = 13'd0;

assign l2_filter_data_ce0 = dataflow_in_loop_TOP_LOOP37548_U0_l2_filter_data_ce0;

assign l2_filter_data_ce1 = 1'b0;

assign l2_filter_data_d0 = 16'd0;

assign l2_filter_data_d1 = 16'd0;

assign l2_filter_data_we0 = 1'b0;

assign l2_filter_data_we1 = 1'b0;

assign out_data_address0 = 13'd0;

assign out_data_address1 = dataflow_in_loop_TOP_LOOP37548_U0_out_data_address1;

assign out_data_ce0 = 1'b0;

assign out_data_ce1 = dataflow_in_loop_TOP_LOOP37548_U0_out_data_ce1;

assign out_data_d0 = 64'd0;

assign out_data_d1 = dataflow_in_loop_TOP_LOOP37548_U0_out_data_d1;

assign out_data_we0 = 1'b0;

assign out_data_we1 = dataflow_in_loop_TOP_LOOP37548_U0_out_data_we1;

assign out_data_write = dataflow_in_loop_TOP_LOOP37548_U0_out_data_write;

endmodule //td_fused_top_tdf7_18
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf7_accum_1 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        accum_in_0_address0,
        accum_in_0_ce0,
        accum_in_0_q0,
        accum_in_0_address1,
        accum_in_0_ce1,
        accum_in_0_q1,
        accum_out_address0,
        accum_out_ce0,
        accum_out_we0,
        accum_out_d0,
        accum_out_address1,
        accum_out_ce1,
        accum_out_we1,
        accum_out_d1
);

parameter    ap_ST_fsm_state1 = 8'd1;
parameter    ap_ST_fsm_pp0_stage0 = 8'd2;
parameter    ap_ST_fsm_pp0_stage1 = 8'd4;
parameter    ap_ST_fsm_pp0_stage2 = 8'd8;
parameter    ap_ST_fsm_pp0_stage3 = 8'd16;
parameter    ap_ST_fsm_state12 = 8'd32;
parameter    ap_ST_fsm_state13 = 8'd64;
parameter    ap_ST_fsm_state14 = 8'd128;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [8:0] accum_in_0_address0;
output   accum_in_0_ce0;
input  [15:0] accum_in_0_q0;
output  [8:0] accum_in_0_address1;
output   accum_in_0_ce1;
input  [15:0] accum_in_0_q1;
output  [2:0] accum_out_address0;
output   accum_out_ce0;
output   accum_out_we0;
output  [15:0] accum_out_d0;
output  [2:0] accum_out_address1;
output   accum_out_ce1;
output   accum_out_we1;
output  [15:0] accum_out_d1;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg[8:0] accum_in_0_address0;
reg accum_in_0_ce0;
reg[8:0] accum_in_0_address1;
reg accum_in_0_ce1;
reg accum_out_ce0;
reg accum_out_we0;
reg accum_out_ce1;
reg accum_out_we1;

reg    ap_done_reg;
  reg   [7:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg   [8:0] x_reg_168;
reg   [15:0] psum_7_08_reg_180;
reg   [15:0] psum_6_07_reg_192;
reg   [15:0] psum_5_06_reg_204;
reg   [15:0] psum_4_05_reg_216;
reg   [15:0] psum_3_04_reg_228;
reg   [15:0] psum_2_03_reg_240;
reg   [15:0] psum_1_02_reg_252;
reg   [15:0] psum_0_01_reg_264;
wire   [0:0] icmp_ln132_fu_321_p2;
reg   [0:0] icmp_ln132_reg_492;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state6_pp0_stage0_iter1;
wire    ap_block_state10_pp0_stage0_iter2;
wire    ap_block_pp0_stage0_11001;
reg   [0:0] icmp_ln132_reg_492_pp0_iter1_reg;
reg   [0:0] icmp_ln132_reg_492_pp0_iter2_reg;
reg   [15:0] accum_in_0_load_reg_506;
wire    ap_CS_fsm_pp0_stage1;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_state3_pp0_stage1_iter0;
wire    ap_block_state7_pp0_stage1_iter1;
wire    ap_block_state11_pp0_stage1_iter2;
wire    ap_block_pp0_stage1_11001;
reg   [15:0] accum_in_0_load_15_reg_511;
reg   [15:0] accum_in_0_load_16_reg_526;
wire    ap_CS_fsm_pp0_stage2;
wire    ap_block_state4_pp0_stage2_iter0;
wire    ap_block_state8_pp0_stage2_iter1;
wire    ap_block_pp0_stage2_11001;
reg   [15:0] accum_in_0_load_17_reg_531;
wire   [8:0] add_ln132_fu_387_p2;
reg   [8:0] add_ln132_reg_546;
wire    ap_CS_fsm_pp0_stage3;
wire    ap_block_state5_pp0_stage3_iter0;
wire    ap_block_state9_pp0_stage3_iter1;
wire    ap_block_pp0_stage3_11001;
reg   [15:0] accum_in_0_load_18_reg_551;
reg   [15:0] accum_in_0_load_19_reg_556;
reg   [15:0] accum_in_0_load_20_reg_571;
reg    ap_enable_reg_pp0_iter1;
reg   [15:0] accum_in_0_load_21_reg_576;
wire   [15:0] grp_fu_305_p2;
wire   [15:0] grp_fu_310_p2;
reg    ap_enable_reg_pp0_iter2;
wire   [3:0] add_ln140_fu_432_p2;
wire    ap_CS_fsm_state13;
wire   [0:0] tmp_fu_415_p3;
reg    ap_block_state1;
wire    ap_block_pp0_stage2_subdone;
reg    ap_condition_pp0_exit_iter0_state4;
wire    ap_block_pp0_stage3_subdone;
wire    ap_block_pp0_stage1_subdone;
reg   [8:0] ap_phi_mux_x_phi_fu_172_p4;
wire    ap_block_pp0_stage0;
wire   [15:0] ap_phi_mux_psum_7_08_phi_fu_184_p4;
wire    ap_block_pp0_stage1;
wire   [15:0] ap_phi_mux_psum_6_07_phi_fu_196_p4;
wire   [15:0] ap_phi_mux_psum_5_06_phi_fu_208_p4;
wire   [15:0] ap_phi_mux_psum_4_05_phi_fu_220_p4;
wire   [15:0] ap_phi_mux_psum_3_04_phi_fu_232_p4;
wire    ap_block_pp0_stage3;
wire   [15:0] ap_phi_mux_psum_2_03_phi_fu_244_p4;
wire    ap_block_pp0_stage2;
reg   [3:0] q_reg_276;
wire    ap_CS_fsm_state12;
reg   [15:0] ap_phi_mux_phi_ln152_phi_fu_290_p8;
wire   [2:0] trunc_ln140_fu_428_p1;
wire   [63:0] zext_ln132_fu_327_p1;
wire   [63:0] zext_ln136_fu_338_p1;
wire   [63:0] zext_ln136_1_fu_349_p1;
wire   [63:0] zext_ln136_2_fu_360_p1;
wire   [63:0] zext_ln136_3_fu_371_p1;
wire   [63:0] zext_ln136_4_fu_382_p1;
wire   [63:0] zext_ln136_5_fu_399_p1;
wire   [63:0] zext_ln136_6_fu_410_p1;
wire   [63:0] zext_ln140_fu_423_p1;
wire   [63:0] zext_ln140_1_fu_444_p1;
reg   [15:0] grp_fu_305_p0;
reg   [15:0] grp_fu_305_p1;
reg   [15:0] grp_fu_310_p0;
reg   [15:0] grp_fu_310_p1;
wire   [8:0] or_ln136_fu_332_p2;
wire   [8:0] or_ln136_1_fu_343_p2;
wire   [8:0] or_ln136_2_fu_354_p2;
wire   [8:0] or_ln136_3_fu_365_p2;
wire   [8:0] or_ln136_4_fu_376_p2;
wire   [8:0] or_ln136_5_fu_393_p2;
wire   [8:0] or_ln136_6_fu_404_p2;
wire   [2:0] or_ln140_fu_438_p2;
wire   [0:0] icmp_ln152_fu_449_p2;
wire   [0:0] icmp_ln152_1_fu_463_p2;
wire   [15:0] select_ln152_fu_455_p3;
wire   [0:0] icmp_ln152_2_fu_477_p2;
wire   [15:0] select_ln152_1_fu_469_p3;
wire    ap_CS_fsm_state14;
reg   [7:0] ap_NS_fsm;
wire    ap_block_pp0_stage0_subdone;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
reg    ap_condition_514;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 8'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
end

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U421(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(grp_fu_305_p0),
    .din1(grp_fu_305_p1),
    .dout(grp_fu_305_p2)
);

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U422(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(grp_fu_310_p0),
    .din1(grp_fu_310_p1),
    .dout(grp_fu_310_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state14)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage2_subdone) & (1'b1 == ap_condition_pp0_exit_iter0_state4) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage3_subdone) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b0)) | ((1'b0 == ap_block_pp0_stage3_subdone) & (1'b1 == ap_CS_fsm_pp0_stage3)))) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end else if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter2 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state12)) begin
        q_reg_276 <= 4'd0;
    end else if (((tmp_fu_415_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state13))) begin
        q_reg_276 <= add_ln140_fu_432_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln132_reg_492 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        x_reg_168 <= add_ln132_reg_546;
    end else if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        x_reg_168 <= 9'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage1_11001) & (icmp_ln132_reg_492 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
        accum_in_0_load_15_reg_511 <= accum_in_0_q0;
        accum_in_0_load_reg_506 <= accum_in_0_q1;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2_11001) & (icmp_ln132_reg_492 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
        accum_in_0_load_16_reg_526 <= accum_in_0_q1;
        accum_in_0_load_17_reg_531 <= accum_in_0_q0;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage3_11001) & (icmp_ln132_reg_492 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
        accum_in_0_load_18_reg_551 <= accum_in_0_q1;
        accum_in_0_load_19_reg_556 <= accum_in_0_q0;
        add_ln132_reg_546 <= add_ln132_fu_387_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln132_reg_492 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        accum_in_0_load_20_reg_571 <= accum_in_0_q1;
        accum_in_0_load_21_reg_576 <= accum_in_0_q0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln132_reg_492 <= icmp_ln132_fu_321_p2;
        icmp_ln132_reg_492_pp0_iter1_reg <= icmp_ln132_reg_492;
        icmp_ln132_reg_492_pp0_iter2_reg <= icmp_ln132_reg_492_pp0_iter1_reg;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln132_reg_492_pp0_iter1_reg == 1'd1) & (1'b0 == ap_block_pp0_stage2_11001) & (1'b1 == ap_CS_fsm_pp0_stage2) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        psum_0_01_reg_264 <= grp_fu_305_p2;
        psum_1_02_reg_252 <= grp_fu_310_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln132_reg_492_pp0_iter1_reg == 1'd1) & (1'b0 == ap_block_pp0_stage3_11001) & (1'b1 == ap_CS_fsm_pp0_stage3) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        psum_2_03_reg_240 <= grp_fu_305_p2;
        psum_3_04_reg_228 <= grp_fu_310_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln132_reg_492_pp0_iter1_reg == 1'd1) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        psum_4_05_reg_216 <= grp_fu_305_p2;
        psum_5_06_reg_204 <= grp_fu_310_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln132_reg_492_pp0_iter2_reg == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        psum_6_07_reg_192 <= grp_fu_305_p2;
        psum_7_08_reg_180 <= grp_fu_310_p2;
    end
end

always @ (*) begin
    if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
        if (((1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            accum_in_0_address0 = zext_ln136_6_fu_410_p1;
        end else if (((1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            accum_in_0_address0 = zext_ln136_4_fu_382_p1;
        end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            accum_in_0_address0 = zext_ln136_2_fu_360_p1;
        end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            accum_in_0_address0 = zext_ln136_fu_338_p1;
        end else begin
            accum_in_0_address0 = 'bx;
        end
    end else begin
        accum_in_0_address0 = 'bx;
    end
end

always @ (*) begin
    if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
        if (((1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            accum_in_0_address1 = zext_ln136_5_fu_399_p1;
        end else if (((1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            accum_in_0_address1 = zext_ln136_3_fu_371_p1;
        end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            accum_in_0_address1 = zext_ln136_1_fu_349_p1;
        end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            accum_in_0_address1 = zext_ln132_fu_327_p1;
        end else begin
            accum_in_0_address1 = 'bx;
        end
    end else begin
        accum_in_0_address1 = 'bx;
    end
end

always @ (*) begin
    if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage3_11001) & (1'b1 == ap_CS_fsm_pp0_stage3)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2_11001) & (1'b1 == ap_CS_fsm_pp0_stage2)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1)))) begin
        accum_in_0_ce0 = 1'b1;
    end else begin
        accum_in_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage3_11001) & (1'b1 == ap_CS_fsm_pp0_stage3)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2_11001) & (1'b1 == ap_CS_fsm_pp0_stage2)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1)))) begin
        accum_in_0_ce1 = 1'b1;
    end else begin
        accum_in_0_ce1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state13)) begin
        accum_out_ce0 = 1'b1;
    end else begin
        accum_out_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state13)) begin
        accum_out_ce1 = 1'b1;
    end else begin
        accum_out_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((tmp_fu_415_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state13))) begin
        accum_out_we0 = 1'b1;
    end else begin
        accum_out_we0 = 1'b0;
    end
end

always @ (*) begin
    if (((tmp_fu_415_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state13))) begin
        accum_out_we1 = 1'b1;
    end else begin
        accum_out_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((icmp_ln132_reg_492 == 1'd0)) begin
        ap_condition_pp0_exit_iter0_state4 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state4 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state14)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((tmp_fu_415_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state13))) begin
        if ((trunc_ln140_fu_428_p1 == 3'd0)) begin
            ap_phi_mux_phi_ln152_phi_fu_290_p8 = psum_0_01_reg_264;
        end else if ((1'b1 == ap_condition_514)) begin
            ap_phi_mux_phi_ln152_phi_fu_290_p8 = psum_6_07_reg_192;
        end else if ((trunc_ln140_fu_428_p1 == 3'd4)) begin
            ap_phi_mux_phi_ln152_phi_fu_290_p8 = psum_4_05_reg_216;
        end else if ((trunc_ln140_fu_428_p1 == 3'd2)) begin
            ap_phi_mux_phi_ln152_phi_fu_290_p8 = psum_2_03_reg_240;
        end else begin
            ap_phi_mux_phi_ln152_phi_fu_290_p8 = 'bx;
        end
    end else begin
        ap_phi_mux_phi_ln152_phi_fu_290_p8 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0) & (icmp_ln132_reg_492 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_x_phi_fu_172_p4 = add_ln132_reg_546;
    end else begin
        ap_phi_mux_x_phi_fu_172_p4 = x_reg_168;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state14)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_305_p0 = ap_phi_mux_psum_6_07_phi_fu_196_p4;
    end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_305_p0 = ap_phi_mux_psum_4_05_phi_fu_220_p4;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
        grp_fu_305_p0 = ap_phi_mux_psum_2_03_phi_fu_244_p4;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
        grp_fu_305_p0 = grp_fu_305_p2;
    end else begin
        grp_fu_305_p0 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_305_p1 = accum_in_0_load_20_reg_571;
    end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_305_p1 = accum_in_0_load_18_reg_551;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
        grp_fu_305_p1 = accum_in_0_load_16_reg_526;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
        grp_fu_305_p1 = accum_in_0_load_reg_506;
    end else begin
        grp_fu_305_p1 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_310_p0 = ap_phi_mux_psum_7_08_phi_fu_184_p4;
    end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_310_p0 = ap_phi_mux_psum_5_06_phi_fu_208_p4;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
        grp_fu_310_p0 = ap_phi_mux_psum_3_04_phi_fu_232_p4;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
        grp_fu_310_p0 = grp_fu_310_p2;
    end else begin
        grp_fu_310_p0 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_310_p1 = accum_in_0_load_21_reg_576;
    end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_310_p1 = accum_in_0_load_19_reg_556;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
        grp_fu_310_p1 = accum_in_0_load_17_reg_531;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
        grp_fu_310_p1 = accum_in_0_load_15_reg_511;
    end else begin
        grp_fu_310_p1 = 'bx;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_pp0_stage1 : begin
            if ((~((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter2 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0)) & (1'b0 == ap_block_pp0_stage1_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage2;
            end else if (((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter2 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
                ap_NS_fsm = ap_ST_fsm_state12;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end
        end
        ap_ST_fsm_pp0_stage2 : begin
            if ((~((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2_subdone) & (icmp_ln132_reg_492 == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b0)) & (1'b0 == ap_block_pp0_stage2_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage3;
            end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2_subdone) & (icmp_ln132_reg_492 == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
                ap_NS_fsm = ap_ST_fsm_state12;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage2;
            end
        end
        ap_ST_fsm_pp0_stage3 : begin
            if ((1'b0 == ap_block_pp0_stage3_subdone)) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage3;
            end
        end
        ap_ST_fsm_state12 : begin
            ap_NS_fsm = ap_ST_fsm_state13;
        end
        ap_ST_fsm_state13 : begin
            if (((tmp_fu_415_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state13))) begin
                ap_NS_fsm = ap_ST_fsm_state13;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state14;
            end
        end
        ap_ST_fsm_state14 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign accum_out_address0 = zext_ln140_1_fu_444_p1;

assign accum_out_address1 = zext_ln140_fu_423_p1;

assign accum_out_d0 = ((icmp_ln152_2_fu_477_p2[0:0] == 1'b1) ? psum_5_06_reg_204 : select_ln152_1_fu_469_p3);

assign accum_out_d1 = ap_phi_mux_phi_ln152_phi_fu_290_p8;

assign add_ln132_fu_387_p2 = (x_reg_168 + 9'd8);

assign add_ln140_fu_432_p2 = (q_reg_276 + 4'd2);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_pp0_stage1 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_pp0_stage2 = ap_CS_fsm[32'd3];

assign ap_CS_fsm_pp0_stage3 = ap_CS_fsm[32'd4];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state12 = ap_CS_fsm[32'd5];

assign ap_CS_fsm_state13 = ap_CS_fsm[32'd6];

assign ap_CS_fsm_state14 = ap_CS_fsm[32'd7];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1_subdone = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage2 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage2_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage2_subdone = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage3 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage3_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage3_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((ap_done_reg == 1'b1) | (ap_start == 1'b0));
end

assign ap_block_state10_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state11_pp0_stage1_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage1_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage2_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage3_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage1_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage2_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state9_pp0_stage3_iter1 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_condition_514 = (~(trunc_ln140_fu_428_p1 == 3'd0) & ~(trunc_ln140_fu_428_p1 == 3'd4) & ~(trunc_ln140_fu_428_p1 == 3'd2));
end

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign ap_phi_mux_psum_2_03_phi_fu_244_p4 = grp_fu_305_p2;

assign ap_phi_mux_psum_3_04_phi_fu_232_p4 = grp_fu_310_p2;

assign ap_phi_mux_psum_4_05_phi_fu_220_p4 = grp_fu_305_p2;

assign ap_phi_mux_psum_5_06_phi_fu_208_p4 = grp_fu_310_p2;

assign ap_phi_mux_psum_6_07_phi_fu_196_p4 = grp_fu_305_p2;

assign ap_phi_mux_psum_7_08_phi_fu_184_p4 = grp_fu_310_p2;

assign icmp_ln132_fu_321_p2 = ((ap_phi_mux_x_phi_fu_172_p4 < 9'd288) ? 1'b1 : 1'b0);

assign icmp_ln152_1_fu_463_p2 = ((or_ln140_fu_438_p2 == 3'd3) ? 1'b1 : 1'b0);

assign icmp_ln152_2_fu_477_p2 = ((or_ln140_fu_438_p2 == 3'd5) ? 1'b1 : 1'b0);

assign icmp_ln152_fu_449_p2 = ((or_ln140_fu_438_p2 == 3'd1) ? 1'b1 : 1'b0);

assign or_ln136_1_fu_343_p2 = (x_reg_168 | 9'd2);

assign or_ln136_2_fu_354_p2 = (x_reg_168 | 9'd3);

assign or_ln136_3_fu_365_p2 = (x_reg_168 | 9'd4);

assign or_ln136_4_fu_376_p2 = (x_reg_168 | 9'd5);

assign or_ln136_5_fu_393_p2 = (x_reg_168 | 9'd6);

assign or_ln136_6_fu_404_p2 = (x_reg_168 | 9'd7);

assign or_ln136_fu_332_p2 = (ap_phi_mux_x_phi_fu_172_p4 | 9'd1);

assign or_ln140_fu_438_p2 = (trunc_ln140_fu_428_p1 | 3'd1);

assign select_ln152_1_fu_469_p3 = ((icmp_ln152_1_fu_463_p2[0:0] == 1'b1) ? psum_3_04_reg_228 : select_ln152_fu_455_p3);

assign select_ln152_fu_455_p3 = ((icmp_ln152_fu_449_p2[0:0] == 1'b1) ? psum_1_02_reg_252 : psum_7_08_reg_180);

assign tmp_fu_415_p3 = q_reg_276[32'd3];

assign trunc_ln140_fu_428_p1 = q_reg_276[2:0];

assign zext_ln132_fu_327_p1 = ap_phi_mux_x_phi_fu_172_p4;

assign zext_ln136_1_fu_349_p1 = or_ln136_1_fu_343_p2;

assign zext_ln136_2_fu_360_p1 = or_ln136_2_fu_354_p2;

assign zext_ln136_3_fu_371_p1 = or_ln136_3_fu_365_p2;

assign zext_ln136_4_fu_382_p1 = or_ln136_4_fu_376_p2;

assign zext_ln136_5_fu_399_p1 = or_ln136_5_fu_393_p2;

assign zext_ln136_6_fu_410_p1 = or_ln136_6_fu_404_p2;

assign zext_ln136_fu_338_p1 = or_ln136_fu_332_p2;

assign zext_ln140_1_fu_444_p1 = or_ln140_fu_438_p2;

assign zext_ln140_fu_423_p1 = q_reg_276;

endmodule //td_fused_top_tdf7_accum_1
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf7_accum_2 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        accum_in_6,
        accum_in_6_ap_vld,
        accum_in_address0,
        accum_in_ce0,
        accum_in_q0
);

parameter    ap_ST_fsm_state1 = 7'd1;
parameter    ap_ST_fsm_state2 = 7'd2;
parameter    ap_ST_fsm_state3 = 7'd4;
parameter    ap_ST_fsm_state4 = 7'd8;
parameter    ap_ST_fsm_state5 = 7'd16;
parameter    ap_ST_fsm_state6 = 7'd32;
parameter    ap_ST_fsm_state7 = 7'd64;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [15:0] accum_in_6;
output   accum_in_6_ap_vld;
output  [2:0] accum_in_address0;
output   accum_in_ce0;
input  [15:0] accum_in_q0;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg[15:0] accum_in_6;
reg accum_in_6_ap_vld;
reg accum_in_ce0;

reg    ap_done_reg;
  reg   [6:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
wire   [3:0] add_ln164_fu_74_p2;
reg   [3:0] add_ln164_reg_91;
wire    ap_CS_fsm_state2;
wire   [0:0] icmp_ln164_fu_85_p2;
wire    ap_CS_fsm_state3;
wire   [15:0] grp_fu_68_p2;
wire    ap_CS_fsm_state7;
reg   [3:0] i_1_1_reg_44;
reg    ap_block_state1;
reg   [15:0] sum_01_reg_55;
wire   [63:0] zext_ln164_fu_80_p1;
reg   [15:0] accum_in_6_preg;
reg   [6:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 7'd1;
#0 accum_in_6_preg = 16'd0;
end

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U425(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(sum_01_reg_55),
    .din1(accum_in_q0),
    .dout(grp_fu_68_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        accum_in_6_preg <= 16'd0;
    end else begin
        if (((icmp_ln164_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
            accum_in_6_preg <= sum_01_reg_55;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if (((icmp_ln164_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        i_1_1_reg_44 <= 4'd0;
    end else if ((1'b1 == ap_CS_fsm_state7)) begin
        i_1_1_reg_44 <= add_ln164_reg_91;
    end
end

always @ (posedge ap_clk) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        sum_01_reg_55 <= 16'd0;
    end else if ((1'b1 == ap_CS_fsm_state7)) begin
        sum_01_reg_55 <= grp_fu_68_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        add_ln164_reg_91 <= add_ln164_fu_74_p2;
    end
end

always @ (*) begin
    if (((icmp_ln164_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        accum_in_6 = sum_01_reg_55;
    end else begin
        accum_in_6 = accum_in_6_preg;
    end
end

always @ (*) begin
    if (((icmp_ln164_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        accum_in_6_ap_vld = 1'b1;
    end else begin
        accum_in_6_ap_vld = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        accum_in_ce0 = 1'b1;
    end else begin
        accum_in_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln164_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln164_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_state2 : begin
            if (((icmp_ln164_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end
        end
        ap_ST_fsm_state3 : begin
            ap_NS_fsm = ap_ST_fsm_state4;
        end
        ap_ST_fsm_state4 : begin
            ap_NS_fsm = ap_ST_fsm_state5;
        end
        ap_ST_fsm_state5 : begin
            ap_NS_fsm = ap_ST_fsm_state6;
        end
        ap_ST_fsm_state6 : begin
            ap_NS_fsm = ap_ST_fsm_state7;
        end
        ap_ST_fsm_state7 : begin
            ap_NS_fsm = ap_ST_fsm_state2;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign accum_in_address0 = zext_ln164_fu_80_p1;

assign add_ln164_fu_74_p2 = (i_1_1_reg_44 + 4'd1);

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state7 = ap_CS_fsm[32'd6];

always @ (*) begin
    ap_block_state1 = ((ap_done_reg == 1'b1) | (ap_start == 1'b0));
end

assign icmp_ln164_fu_85_p2 = ((i_1_1_reg_44 == 4'd8) ? 1'b1 : 1'b0);

assign zext_ln164_fu_80_p1 = i_1_1_reg_44;

endmodule //td_fused_top_tdf7_accum_2
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_tdf7_adjustments_ram (addr0, ce0, q0, addr1, ce1, d1, we1,  clk);

parameter DWIDTH = 48;
parameter AWIDTH = 8;
parameter MEM_SIZE = 256;

input[AWIDTH-1:0] addr0;
input ce0;
output wire[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
input clk;

 reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];
wire [AWIDTH-1:0] addr0_t0; 
reg [AWIDTH-1:0] addr0_t1; 
reg [DWIDTH-1:0] q0_t0;
reg [DWIDTH-1:0] q0_t1;
wire [AWIDTH-1:0] addr1_t0; 
reg [AWIDTH-1:0] addr1_t1; 
wire [DWIDTH-1:0] d1_t0; 
wire we1_t0; 
reg [DWIDTH-1:0] d1_t1; 
reg we1_t1; 


assign addr0_t0 = addr0;
assign q0 = q0_t1;
assign addr1_t0 = addr1;
assign d1_t0 = d1;
assign we1_t0 = we1;

always @(posedge clk)  
begin
    if (ce0) 
    begin
        addr0_t1 <= addr0_t0; 
        q0_t1 <= q0_t0;
    end
    if (ce1) 
    begin
        addr1_t1 <= addr1_t0; 
        d1_t1 <= d1_t0;
        we1_t1 <= we1_t0;
    end
end


always @(posedge clk)  
begin 
    if (ce0) begin
        q0_t0 <= ram[addr0_t1];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1_t1) 
            ram[addr1_t1] <= d1_t1; 
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_tdf7_adjustments(
    reset,
    clk,
    address0,
    ce0,
    q0,
    address1,
    ce1,
    we1,
    d1);

parameter DataWidth = 32'd48;
parameter AddressRange = 32'd256;
parameter AddressWidth = 32'd8;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;



td_fused_top_tdf7_adjustments_ram td_fused_top_tdf7_adjustments_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 )
);

endmodule

// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf7_adjust (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        sums_read,
        adjustments_address0,
        adjustments_ce0,
        adjustments_q0,
        indices_23_dout,
        indices_23_empty_n,
        indices_23_read,
        indices_23_out_din,
        indices_23_out_full_n,
        indices_23_out_write,
        ap_return
);

parameter    ap_ST_fsm_state1 = 17'd1;
parameter    ap_ST_fsm_state2 = 17'd2;
parameter    ap_ST_fsm_state3 = 17'd4;
parameter    ap_ST_fsm_state4 = 17'd8;
parameter    ap_ST_fsm_state5 = 17'd16;
parameter    ap_ST_fsm_state6 = 17'd32;
parameter    ap_ST_fsm_state7 = 17'd64;
parameter    ap_ST_fsm_state8 = 17'd128;
parameter    ap_ST_fsm_state9 = 17'd256;
parameter    ap_ST_fsm_state10 = 17'd512;
parameter    ap_ST_fsm_state11 = 17'd1024;
parameter    ap_ST_fsm_state12 = 17'd2048;
parameter    ap_ST_fsm_state13 = 17'd4096;
parameter    ap_ST_fsm_state14 = 17'd8192;
parameter    ap_ST_fsm_state15 = 17'd16384;
parameter    ap_ST_fsm_state16 = 17'd32768;
parameter    ap_ST_fsm_state17 = 17'd65536;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
input  [15:0] sums_read;
output  [7:0] adjustments_address0;
output   adjustments_ce0;
input  [47:0] adjustments_q0;
input  [12:0] indices_23_dout;
input   indices_23_empty_n;
output   indices_23_read;
output  [12:0] indices_23_out_din;
input   indices_23_out_full_n;
output   indices_23_out_write;
output  [15:0] ap_return;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg adjustments_ce0;
reg indices_23_read;
reg indices_23_out_write;

reg    ap_done_reg;
  reg   [16:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    indices_23_blk_n;
reg    indices_23_out_blk_n;
wire    ap_CS_fsm_state4;
reg   [15:0] tmp_26_i_i_reg_183;
reg   [15:0] tmp_27_i_i_reg_188;
wire   [15:0] grp_fu_93_p2;
reg   [15:0] sub_i_i_i_reg_193;
wire    ap_CS_fsm_state8;
wire    ap_CS_fsm_state9;
wire   [15:0] grp_fu_98_p2;
reg   [15:0] mul_i_i_i_reg_203;
wire    ap_CS_fsm_state12;
wire    ap_CS_fsm_state13;
wire   [63:0] zext_ln220_fu_106_p1;
reg    ap_block_state1;
wire    ap_CS_fsm_state2;
wire    ap_CS_fsm_state3;
wire   [15:0] grp_fu_89_p1;
wire   [15:0] grp_fu_93_p1;
wire   [15:0] grp_fu_98_p1;
wire   [7:0] trunc_ln251_fu_102_p1;
wire   [15:0] trunc_ln220_fu_111_p1;
wire   [15:0] grp_fu_89_p2;
wire    ap_CS_fsm_state17;
wire   [15:0] bitcast_ln648_fu_148_p1;
wire   [0:0] tmp_fu_152_p3;
reg   [16:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 17'd1;
end

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U429(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(mul_i_i_i_reg_203),
    .din1(grp_fu_89_p1),
    .dout(grp_fu_89_p2)
);

td_fused_top_hsub_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hsub_16ns_16ns_16_5_full_dsp_1_U430(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(sums_read),
    .din1(grp_fu_93_p1),
    .dout(grp_fu_93_p2)
);

td_fused_top_hmul_16ns_16ns_16_4_max_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hmul_16ns_16ns_16_4_max_dsp_1_U431(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(sub_i_i_i_reg_193),
    .din1(grp_fu_98_p1),
    .dout(grp_fu_98_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state17)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state12)) begin
        mul_i_i_i_reg_203 <= grp_fu_98_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state8)) begin
        sub_i_i_i_reg_193 <= grp_fu_93_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        tmp_26_i_i_reg_183 <= {{adjustments_q0[31:16]}};
        tmp_27_i_i_reg_188 <= {{adjustments_q0[47:32]}};
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state2) | (~((indices_23_out_full_n == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1)))) begin
        adjustments_ce0 = 1'b1;
    end else begin
        adjustments_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state17)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state17)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_23_blk_n = indices_23_empty_n;
    end else begin
        indices_23_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_23_out_blk_n = indices_23_out_full_n;
    end else begin
        indices_23_out_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((indices_23_out_full_n == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_23_out_write = 1'b1;
    end else begin
        indices_23_out_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((indices_23_out_full_n == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_23_read = 1'b1;
    end else begin
        indices_23_read = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((indices_23_out_full_n == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_state2 : begin
            ap_NS_fsm = ap_ST_fsm_state3;
        end
        ap_ST_fsm_state3 : begin
            ap_NS_fsm = ap_ST_fsm_state4;
        end
        ap_ST_fsm_state4 : begin
            ap_NS_fsm = ap_ST_fsm_state5;
        end
        ap_ST_fsm_state5 : begin
            ap_NS_fsm = ap_ST_fsm_state6;
        end
        ap_ST_fsm_state6 : begin
            ap_NS_fsm = ap_ST_fsm_state7;
        end
        ap_ST_fsm_state7 : begin
            ap_NS_fsm = ap_ST_fsm_state8;
        end
        ap_ST_fsm_state8 : begin
            ap_NS_fsm = ap_ST_fsm_state9;
        end
        ap_ST_fsm_state9 : begin
            ap_NS_fsm = ap_ST_fsm_state10;
        end
        ap_ST_fsm_state10 : begin
            ap_NS_fsm = ap_ST_fsm_state11;
        end
        ap_ST_fsm_state11 : begin
            ap_NS_fsm = ap_ST_fsm_state12;
        end
        ap_ST_fsm_state12 : begin
            ap_NS_fsm = ap_ST_fsm_state13;
        end
        ap_ST_fsm_state13 : begin
            ap_NS_fsm = ap_ST_fsm_state14;
        end
        ap_ST_fsm_state14 : begin
            ap_NS_fsm = ap_ST_fsm_state15;
        end
        ap_ST_fsm_state15 : begin
            ap_NS_fsm = ap_ST_fsm_state16;
        end
        ap_ST_fsm_state16 : begin
            ap_NS_fsm = ap_ST_fsm_state17;
        end
        ap_ST_fsm_state17 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign adjustments_address0 = zext_ln220_fu_106_p1;

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state12 = ap_CS_fsm[32'd11];

assign ap_CS_fsm_state13 = ap_CS_fsm[32'd12];

assign ap_CS_fsm_state17 = ap_CS_fsm[32'd16];

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

assign ap_CS_fsm_state8 = ap_CS_fsm[32'd7];

assign ap_CS_fsm_state9 = ap_CS_fsm[32'd8];

always @ (*) begin
    ap_block_state1 = ((indices_23_out_full_n == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0));
end

assign ap_return = ((tmp_fu_152_p3[0:0] == 1'b1) ? 16'd0 : grp_fu_89_p2);

assign bitcast_ln648_fu_148_p1 = grp_fu_89_p2;

assign grp_fu_89_p1 = tmp_27_i_i_reg_188;

assign grp_fu_93_p1 = trunc_ln220_fu_111_p1;

assign grp_fu_98_p1 = tmp_26_i_i_reg_183;

assign indices_23_out_din = indices_23_dout;

assign tmp_fu_152_p3 = bitcast_ln648_fu_148_p1[32'd15];

assign trunc_ln220_fu_111_p1 = adjustments_q0[15:0];

assign trunc_ln251_fu_102_p1 = indices_23_dout[7:0];

assign zext_ln220_fu_106_p1 = trunc_ln251_fu_102_p1;

endmodule //td_fused_top_tdf7_adjust
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf7_dot_product (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        ifmap_vec_address0,
        ifmap_vec_ce0,
        ifmap_vec_q0,
        weight_vecs_0_address0,
        weight_vecs_0_ce0,
        weight_vecs_0_q0,
        products_0_address0,
        products_0_ce0,
        products_0_we0,
        products_0_d0
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state10 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [8:0] ifmap_vec_address0;
output   ifmap_vec_ce0;
input  [15:0] ifmap_vec_q0;
output  [8:0] weight_vecs_0_address0;
output   weight_vecs_0_ce0;
input  [15:0] weight_vecs_0_q0;
output  [8:0] products_0_address0;
output   products_0_ce0;
output   products_0_we0;
output  [15:0] products_0_d0;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg ifmap_vec_ce0;
reg weight_vecs_0_ce0;
reg products_0_ce0;
reg products_0_we0;

reg    ap_done_reg;
  reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg   [8:0] indvar_flatten17_reg_97;
reg   [7:0] indvar_flatten_reg_108;
reg   [1:0] jj_reg_119;
reg   [5:0] ic_reg_131;
reg   [1:0] ii_reg_142;
wire   [8:0] add_ln147_2_fu_157_p2;
wire    ap_CS_fsm_pp0_stage0;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
wire    ap_block_state4_pp0_stage0_iter2;
wire    ap_block_state5_pp0_stage0_iter3;
wire    ap_block_state6_pp0_stage0_iter4;
wire    ap_block_state7_pp0_stage0_iter5;
wire    ap_block_state8_pp0_stage0_iter6;
wire    ap_block_state9_pp0_stage0_iter7;
wire    ap_block_pp0_stage0_11001;
wire   [0:0] icmp_ln147_fu_163_p2;
reg   [0:0] icmp_ln147_reg_408;
reg   [0:0] icmp_ln147_reg_408_pp0_iter1_reg;
reg   [0:0] icmp_ln147_reg_408_pp0_iter2_reg;
reg   [0:0] icmp_ln147_reg_408_pp0_iter3_reg;
reg   [0:0] icmp_ln147_reg_408_pp0_iter4_reg;
reg   [0:0] icmp_ln147_reg_408_pp0_iter5_reg;
reg   [0:0] icmp_ln147_reg_408_pp0_iter6_reg;
wire   [0:0] icmp_ln148_fu_169_p2;
reg   [0:0] icmp_ln148_reg_412;
wire   [0:0] and_ln147_fu_195_p2;
reg   [0:0] and_ln147_reg_419;
wire   [1:0] add_ln148_fu_201_p2;
reg   [1:0] add_ln148_reg_424;
wire   [5:0] select_ln148_fu_213_p3;
reg   [5:0] select_ln148_reg_429;
wire   [1:0] select_ln148_4_fu_221_p3;
reg   [1:0] select_ln148_4_reg_434;
wire   [4:0] trunc_ln150_fu_229_p1;
reg   [4:0] trunc_ln150_reg_440;
reg   [4:0] trunc_ln150_reg_440_pp0_iter1_reg;
reg   [4:0] trunc_ln150_reg_440_pp0_iter2_reg;
reg   [4:0] trunc_ln150_reg_440_pp0_iter3_reg;
reg   [4:0] trunc_ln150_reg_440_pp0_iter4_reg;
reg   [4:0] trunc_ln150_reg_440_pp0_iter5_reg;
reg   [4:0] trunc_ln150_reg_440_pp0_iter6_reg;
wire   [5:0] add_ln149_fu_233_p2;
wire   [7:0] select_ln148_6_fu_245_p3;
wire   [1:0] select_ln147_5_fu_287_p3;
reg   [1:0] select_ln147_5_reg_455;
reg    ap_enable_reg_pp0_iter1;
wire   [3:0] select_ln148_5_fu_370_p3;
reg   [3:0] select_ln148_5_reg_460;
reg   [3:0] select_ln148_5_reg_460_pp0_iter2_reg;
reg   [3:0] select_ln148_5_reg_460_pp0_iter3_reg;
reg   [3:0] select_ln148_5_reg_460_pp0_iter4_reg;
reg   [3:0] select_ln148_5_reg_460_pp0_iter5_reg;
reg   [3:0] select_ln148_5_reg_460_pp0_iter6_reg;
reg   [15:0] ifmap_vec_load_reg_475;
reg   [15:0] weight_vecs_0_load_reg_480;
wire   [15:0] grp_fu_153_p2;
reg   [15:0] mul_reg_485;
reg    ap_block_state1;
wire    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_flush_enable;
reg    ap_enable_reg_pp0_iter2;
reg    ap_condition_pp0_exit_iter1_state3;
reg    ap_enable_reg_pp0_iter3;
reg    ap_enable_reg_pp0_iter4;
reg    ap_enable_reg_pp0_iter5;
reg    ap_enable_reg_pp0_iter6;
reg    ap_enable_reg_pp0_iter7;
reg   [1:0] ap_phi_mux_jj_phi_fu_123_p4;
wire    ap_block_pp0_stage0;
reg   [1:0] ap_phi_mux_ii_phi_fu_146_p4;
wire   [63:0] p_cast25_fu_386_p1;
wire   [63:0] idxprom30_fu_398_p1;
wire   [0:0] icmp_ln149_fu_189_p2;
wire   [0:0] xor_ln147_fu_183_p2;
wire   [1:0] select_ln147_fu_175_p3;
wire   [0:0] or_ln148_fu_207_p2;
wire   [7:0] add_ln148_2_fu_239_p2;
wire   [3:0] shl_ln_fu_257_p3;
wire   [3:0] zext_ln150_fu_253_p1;
wire   [3:0] sub_ln150_fu_265_p2;
wire   [3:0] zext_ln150_2_fu_271_p1;
wire   [1:0] add_ln147_fu_281_p2;
wire   [3:0] tmp_fu_298_p3;
wire   [3:0] select_ln147_6_cast_fu_294_p1;
wire   [3:0] shl_ln150_mid1_fu_316_p3;
wire   [3:0] zext_ln150_4_fu_312_p1;
wire   [3:0] sub_ln150_2_fu_324_p2;
wire   [3:0] add_ln150_fu_275_p2;
wire   [3:0] empty_74_fu_306_p2;
wire   [3:0] select_ln148_5_cast_fu_344_p1;
wire   [3:0] empty_75_fu_347_p2;
wire   [3:0] select_ln147_6_fu_330_p3;
wire   [3:0] zext_ln150_5_fu_361_p1;
wire   [3:0] add_ln150_2_fu_364_p2;
wire   [3:0] select_ln147_7_fu_337_p3;
wire   [8:0] tmp_50_cast_fu_353_p3;
wire   [8:0] select_ln148_cast_fu_377_p1;
wire   [8:0] empty_76_fu_380_p2;
wire   [8:0] p_fu_392_p3;
wire    ap_CS_fsm_state10;
reg   [2:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
#0 ap_enable_reg_pp0_iter4 = 1'b0;
#0 ap_enable_reg_pp0_iter5 = 1'b0;
#0 ap_enable_reg_pp0_iter6 = 1'b0;
#0 ap_enable_reg_pp0_iter7 = 1'b0;
end

td_fused_top_hmul_16ns_16ns_16_4_max_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hmul_16ns_16ns_16_4_max_dsp_1_U417(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(ifmap_vec_load_reg_475),
    .din1(weight_vecs_0_load_reg_480),
    .dout(grp_fu_153_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state10)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if ((1'b1 == ap_condition_pp0_flush_enable)) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            if ((1'b1 == ap_condition_pp0_exit_iter1_state3)) begin
                ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter0;
            end else if ((1'b1 == 1'b1)) begin
                ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
            end
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter4 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter5 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter5 <= ap_enable_reg_pp0_iter4;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter6 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter6 <= ap_enable_reg_pp0_iter5;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter7 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter7 <= ap_enable_reg_pp0_iter6;
        end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter7 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_fu_163_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ic_reg_131 <= add_ln149_fu_233_p2;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ic_reg_131 <= 6'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_reg_408_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        ii_reg_142 <= select_ln147_5_reg_455;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ii_reg_142 <= 2'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_fu_163_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        indvar_flatten17_reg_97 <= add_ln147_2_fu_157_p2;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indvar_flatten17_reg_97 <= 9'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_fu_163_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        indvar_flatten_reg_108 <= select_ln148_6_fu_245_p3;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indvar_flatten_reg_108 <= 8'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_reg_408 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        jj_reg_119 <= select_ln148_4_reg_434;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        jj_reg_119 <= 2'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_fu_163_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        add_ln148_reg_424 <= add_ln148_fu_201_p2;
        and_ln147_reg_419 <= and_ln147_fu_195_p2;
        icmp_ln148_reg_412 <= icmp_ln148_fu_169_p2;
        select_ln148_reg_429 <= select_ln148_fu_213_p3;
        trunc_ln150_reg_440 <= trunc_ln150_fu_229_p1;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln147_reg_408 <= icmp_ln147_fu_163_p2;
        icmp_ln147_reg_408_pp0_iter1_reg <= icmp_ln147_reg_408;
        trunc_ln150_reg_440_pp0_iter1_reg <= trunc_ln150_reg_440;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        icmp_ln147_reg_408_pp0_iter2_reg <= icmp_ln147_reg_408_pp0_iter1_reg;
        icmp_ln147_reg_408_pp0_iter3_reg <= icmp_ln147_reg_408_pp0_iter2_reg;
        icmp_ln147_reg_408_pp0_iter4_reg <= icmp_ln147_reg_408_pp0_iter3_reg;
        icmp_ln147_reg_408_pp0_iter5_reg <= icmp_ln147_reg_408_pp0_iter4_reg;
        icmp_ln147_reg_408_pp0_iter6_reg <= icmp_ln147_reg_408_pp0_iter5_reg;
        select_ln148_5_reg_460_pp0_iter2_reg <= select_ln148_5_reg_460;
        select_ln148_5_reg_460_pp0_iter3_reg <= select_ln148_5_reg_460_pp0_iter2_reg;
        select_ln148_5_reg_460_pp0_iter4_reg <= select_ln148_5_reg_460_pp0_iter3_reg;
        select_ln148_5_reg_460_pp0_iter5_reg <= select_ln148_5_reg_460_pp0_iter4_reg;
        select_ln148_5_reg_460_pp0_iter6_reg <= select_ln148_5_reg_460_pp0_iter5_reg;
        trunc_ln150_reg_440_pp0_iter2_reg <= trunc_ln150_reg_440_pp0_iter1_reg;
        trunc_ln150_reg_440_pp0_iter3_reg <= trunc_ln150_reg_440_pp0_iter2_reg;
        trunc_ln150_reg_440_pp0_iter4_reg <= trunc_ln150_reg_440_pp0_iter3_reg;
        trunc_ln150_reg_440_pp0_iter5_reg <= trunc_ln150_reg_440_pp0_iter4_reg;
        trunc_ln150_reg_440_pp0_iter6_reg <= trunc_ln150_reg_440_pp0_iter5_reg;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_reg_408_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        ifmap_vec_load_reg_475 <= ifmap_vec_q0;
        weight_vecs_0_load_reg_480 <= weight_vecs_0_q0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_reg_408_pp0_iter5_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        mul_reg_485 <= grp_fu_153_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_reg_408 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        select_ln147_5_reg_455 <= select_ln147_5_fu_287_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_fu_163_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        select_ln148_4_reg_434 <= select_ln148_4_fu_221_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_reg_408 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        select_ln148_5_reg_460 <= select_ln148_5_fu_370_p3;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_condition_pp0_exit_iter1_state3 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter1_state3 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln147_fu_163_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_condition_pp0_flush_enable = 1'b1;
    end else begin
        ap_condition_pp0_flush_enable = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state10)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter7 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln147_reg_408_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        ap_phi_mux_ii_phi_fu_146_p4 = select_ln147_5_reg_455;
    end else begin
        ap_phi_mux_ii_phi_fu_146_p4 = ii_reg_142;
    end
end

always @ (*) begin
    if (((icmp_ln147_reg_408 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_jj_phi_fu_123_p4 = select_ln148_4_reg_434;
    end else begin
        ap_phi_mux_jj_phi_fu_123_p4 = jj_reg_119;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state10)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ifmap_vec_ce0 = 1'b1;
    end else begin
        ifmap_vec_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter7 == 1'b1))) begin
        products_0_ce0 = 1'b1;
    end else begin
        products_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln147_reg_408_pp0_iter6_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter7 == 1'b1))) begin
        products_0_we0 = 1'b1;
    end else begin
        products_0_we0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        weight_vecs_0_ce0 = 1'b1;
    end else begin
        weight_vecs_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((~((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b1)) & ~((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter7 == 1'b1) & (ap_enable_reg_pp0_iter6 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if ((((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter7 == 1'b1) & (ap_enable_reg_pp0_iter6 == 1'b0)) | ((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b1)))) begin
                ap_NS_fsm = ap_ST_fsm_state10;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state10 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln147_2_fu_157_p2 = (indvar_flatten17_reg_97 + 9'd1);

assign add_ln147_fu_281_p2 = (ap_phi_mux_ii_phi_fu_146_p4 + 2'd1);

assign add_ln148_2_fu_239_p2 = (indvar_flatten_reg_108 + 8'd1);

assign add_ln148_fu_201_p2 = (select_ln147_fu_175_p3 + 2'd1);

assign add_ln149_fu_233_p2 = (select_ln148_fu_213_p3 + 6'd1);

assign add_ln150_2_fu_364_p2 = (select_ln147_6_fu_330_p3 + zext_ln150_5_fu_361_p1);

assign add_ln150_fu_275_p2 = (sub_ln150_fu_265_p2 + zext_ln150_2_fu_271_p1);

assign and_ln147_fu_195_p2 = (xor_ln147_fu_183_p2 & icmp_ln149_fu_189_p2);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state10 = ap_CS_fsm[32'd2];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (ap_done_reg == 1'b1));
end

assign ap_block_state2_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter4 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage0_iter5 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage0_iter6 = ~(1'b1 == 1'b1);

assign ap_block_state9_pp0_stage0_iter7 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign empty_74_fu_306_p2 = (tmp_fu_298_p3 - select_ln147_6_cast_fu_294_p1);

assign empty_75_fu_347_p2 = (empty_74_fu_306_p2 + select_ln148_5_cast_fu_344_p1);

assign empty_76_fu_380_p2 = (tmp_50_cast_fu_353_p3 + select_ln148_cast_fu_377_p1);

assign icmp_ln147_fu_163_p2 = ((indvar_flatten17_reg_97 == 9'd288) ? 1'b1 : 1'b0);

assign icmp_ln148_fu_169_p2 = ((indvar_flatten_reg_108 == 8'd96) ? 1'b1 : 1'b0);

assign icmp_ln149_fu_189_p2 = ((ic_reg_131 == 6'd32) ? 1'b1 : 1'b0);

assign idxprom30_fu_398_p1 = p_fu_392_p3;

assign ifmap_vec_address0 = p_cast25_fu_386_p1;

assign or_ln148_fu_207_p2 = (icmp_ln148_fu_169_p2 | and_ln147_fu_195_p2);

assign p_cast25_fu_386_p1 = empty_76_fu_380_p2;

assign p_fu_392_p3 = {{select_ln148_5_reg_460_pp0_iter6_reg}, {trunc_ln150_reg_440_pp0_iter6_reg}};

assign products_0_address0 = idxprom30_fu_398_p1;

assign products_0_d0 = mul_reg_485;

assign select_ln147_5_fu_287_p3 = ((icmp_ln148_reg_412[0:0] == 1'b1) ? add_ln147_fu_281_p2 : ap_phi_mux_ii_phi_fu_146_p4);

assign select_ln147_6_cast_fu_294_p1 = select_ln147_5_fu_287_p3;

assign select_ln147_6_fu_330_p3 = ((icmp_ln148_reg_412[0:0] == 1'b1) ? sub_ln150_2_fu_324_p2 : sub_ln150_fu_265_p2);

assign select_ln147_7_fu_337_p3 = ((icmp_ln148_reg_412[0:0] == 1'b1) ? sub_ln150_2_fu_324_p2 : add_ln150_fu_275_p2);

assign select_ln147_fu_175_p3 = ((icmp_ln148_fu_169_p2[0:0] == 1'b1) ? 2'd0 : ap_phi_mux_jj_phi_fu_123_p4);

assign select_ln148_4_fu_221_p3 = ((and_ln147_fu_195_p2[0:0] == 1'b1) ? add_ln148_fu_201_p2 : select_ln147_fu_175_p3);

assign select_ln148_5_cast_fu_344_p1 = select_ln148_4_reg_434;

assign select_ln148_5_fu_370_p3 = ((and_ln147_reg_419[0:0] == 1'b1) ? add_ln150_2_fu_364_p2 : select_ln147_7_fu_337_p3);

assign select_ln148_6_fu_245_p3 = ((icmp_ln148_fu_169_p2[0:0] == 1'b1) ? 8'd1 : add_ln148_2_fu_239_p2);

assign select_ln148_cast_fu_377_p1 = select_ln148_reg_429;

assign select_ln148_fu_213_p3 = ((or_ln148_fu_207_p2[0:0] == 1'b1) ? 6'd0 : ic_reg_131);

assign shl_ln150_mid1_fu_316_p3 = {{add_ln147_fu_281_p2}, {2'd0}};

assign shl_ln_fu_257_p3 = {{ap_phi_mux_ii_phi_fu_146_p4}, {2'd0}};

assign sub_ln150_2_fu_324_p2 = (shl_ln150_mid1_fu_316_p3 - zext_ln150_4_fu_312_p1);

assign sub_ln150_fu_265_p2 = (shl_ln_fu_257_p3 - zext_ln150_fu_253_p1);

assign tmp_50_cast_fu_353_p3 = {{empty_75_fu_347_p2}, {5'd0}};

assign tmp_fu_298_p3 = {{select_ln147_5_fu_287_p3}, {2'd0}};

assign trunc_ln150_fu_229_p1 = select_ln148_fu_213_p3[4:0];

assign weight_vecs_0_address0 = p_cast25_fu_386_p1;

assign xor_ln147_fu_183_p2 = (icmp_ln148_fu_169_p2 ^ 1'd1);

assign zext_ln150_2_fu_271_p1 = jj_reg_119;

assign zext_ln150_4_fu_312_p1 = add_ln147_fu_281_p2;

assign zext_ln150_5_fu_361_p1 = add_ln148_reg_424;

assign zext_ln150_fu_253_p1 = ap_phi_mux_ii_phi_fu_146_p4;

endmodule //td_fused_top_tdf7_dot_product
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_tdf7_filters_ram (addr0, ce0, q0, addr1, ce1, d1, we1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 17;
parameter MEM_SIZE = 73728;

input[AWIDTH-1:0] addr0;
input ce0;
output wire[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
input clk;

 reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];
wire [AWIDTH-1:0] addr0_t0; 
reg [AWIDTH-1:0] addr0_t1; 
reg [DWIDTH-1:0] q0_t0;
reg [DWIDTH-1:0] q0_t1;
wire [AWIDTH-1:0] addr1_t0; 
reg [AWIDTH-1:0] addr1_t1; 
wire [DWIDTH-1:0] d1_t0; 
wire we1_t0; 
reg [DWIDTH-1:0] d1_t1; 
reg we1_t1; 


assign addr0_t0 = addr0;
assign q0 = q0_t1;
assign addr1_t0 = addr1;
assign d1_t0 = d1;
assign we1_t0 = we1;

always @(posedge clk)  
begin
    if (ce0) 
    begin
        addr0_t1 <= addr0_t0; 
        q0_t1 <= q0_t0;
    end
    if (ce1) 
    begin
        addr1_t1 <= addr1_t0; 
        d1_t1 <= d1_t0;
        we1_t1 <= we1_t0;
    end
end


always @(posedge clk)  
begin 
    if (ce0) begin
        q0_t0 <= ram[addr0_t1];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1_t1) 
            ram[addr1_t1] <= d1_t1; 
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_tdf7_filters(
    reset,
    clk,
    address0,
    ce0,
    q0,
    address1,
    ce1,
    we1,
    d1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd73728;
parameter AddressWidth = 32'd17;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;



td_fused_top_tdf7_filters_ram td_fused_top_tdf7_filters_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 )
);

endmodule

// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf7_get_next_ijk (
        ap_clk,
        ap_rst,
        ap_start,
        start_full_n,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        start_out,
        start_write,
        indices_0_din,
        indices_0_full_n,
        indices_0_write,
        indices_1_din,
        indices_1_full_n,
        indices_1_write,
        indices_2_out_din,
        indices_2_out_full_n,
        indices_2_out_write,
        indices_2_out1_din,
        indices_2_out1_full_n,
        indices_2_out1_write,
        write_r_din,
        write_r_full_n,
        write_r_write
);

parameter    ap_ST_fsm_state1 = 1'd1;

input   ap_clk;
input   ap_rst;
input   ap_start;
input   start_full_n;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output   start_out;
output   start_write;
output  [15:0] indices_0_din;
input   indices_0_full_n;
output   indices_0_write;
output  [15:0] indices_1_din;
input   indices_1_full_n;
output   indices_1_write;
output  [7:0] indices_2_out_din;
input   indices_2_out_full_n;
output   indices_2_out_write;
output  [12:0] indices_2_out1_din;
input   indices_2_out1_full_n;
output   indices_2_out1_write;
output   write_r_din;
input   write_r_full_n;
output   write_r_write;

reg ap_done;
reg ap_idle;
reg start_write;
reg indices_0_write;
reg indices_1_write;
reg indices_2_out_write;
reg indices_2_out1_write;
reg write_r_write;

reg    real_start;
reg    start_once_reg;
reg    ap_done_reg;
  reg   [0:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    internal_ap_ready;
reg   [15:0] i_11;
reg   [15:0] j_11;
reg   [15:0] k_11;
reg    indices_0_blk_n;
reg    indices_1_blk_n;
reg    indices_2_out_blk_n;
reg    indices_2_out1_blk_n;
reg    write_r_blk_n;
reg   [0:0] ap_phi_mux_j_18_flag_0_i_phi_fu_92_p6;
reg    ap_block_state1;
wire   [0:0] icmp_ln188_fu_167_p2;
wire   [0:0] icmp_ln191_fu_180_p2;
reg   [15:0] ap_phi_mux_j_18_new_0_i_phi_fu_106_p6;
wire   [15:0] add_ln190_fu_173_p2;
reg   [15:0] ap_phi_mux_k_18_new_0_i_phi_fu_119_p6;
wire   [15:0] add_ln187_fu_160_p2;
wire   [15:0] select_ln194_fu_198_p3;
wire   [15:0] add_ln193_fu_186_p2;
wire   [0:0] icmp_ln194_fu_192_p2;
reg   [0:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 start_once_reg = 1'b0;
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 1'd1;
#0 i_11 = 16'd0;
#0 j_11 = 16'd0;
#0 k_11 = 16'd0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((~((real_start == 1'b0) | (write_r_full_n == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        start_once_reg <= 1'b0;
    end else begin
        if (((real_start == 1'b1) & (internal_ap_ready == 1'b0))) begin
            start_once_reg <= 1'b1;
        end else if ((internal_ap_ready == 1'b1)) begin
            start_once_reg <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((~((real_start == 1'b0) | (write_r_full_n == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (icmp_ln191_fu_180_p2 == 1'd1) & (icmp_ln188_fu_167_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1))) begin
        i_11 <= select_ln194_fu_198_p3;
    end
end

always @ (posedge ap_clk) begin
    if ((~((real_start == 1'b0) | (write_r_full_n == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (ap_phi_mux_j_18_flag_0_i_phi_fu_92_p6 == 1'd1) & (1'b1 == ap_CS_fsm_state1))) begin
        j_11 <= ap_phi_mux_j_18_new_0_i_phi_fu_106_p6;
    end
end

always @ (posedge ap_clk) begin
    if ((~((real_start == 1'b0) | (write_r_full_n == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        k_11 <= ap_phi_mux_k_18_new_0_i_phi_fu_119_p6;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (write_r_full_n == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((real_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln188_fu_167_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_phi_mux_j_18_flag_0_i_phi_fu_92_p6 = 1'd0;
    end else if ((((icmp_ln191_fu_180_p2 == 1'd0) & (icmp_ln188_fu_167_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1)) | ((icmp_ln191_fu_180_p2 == 1'd1) & (icmp_ln188_fu_167_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1)))) begin
        ap_phi_mux_j_18_flag_0_i_phi_fu_92_p6 = 1'd1;
    end else begin
        ap_phi_mux_j_18_flag_0_i_phi_fu_92_p6 = 'bx;
    end
end

always @ (*) begin
    if (((icmp_ln188_fu_167_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1))) begin
        if ((icmp_ln191_fu_180_p2 == 1'd0)) begin
            ap_phi_mux_j_18_new_0_i_phi_fu_106_p6 = add_ln190_fu_173_p2;
        end else if ((icmp_ln191_fu_180_p2 == 1'd1)) begin
            ap_phi_mux_j_18_new_0_i_phi_fu_106_p6 = 16'd0;
        end else begin
            ap_phi_mux_j_18_new_0_i_phi_fu_106_p6 = 'bx;
        end
    end else begin
        ap_phi_mux_j_18_new_0_i_phi_fu_106_p6 = 'bx;
    end
end

always @ (*) begin
    if (((icmp_ln188_fu_167_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_phi_mux_k_18_new_0_i_phi_fu_119_p6 = add_ln187_fu_160_p2;
    end else if ((((icmp_ln191_fu_180_p2 == 1'd0) & (icmp_ln188_fu_167_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1)) | ((icmp_ln191_fu_180_p2 == 1'd1) & (icmp_ln188_fu_167_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1)))) begin
        ap_phi_mux_k_18_new_0_i_phi_fu_119_p6 = 16'd0;
    end else begin
        ap_phi_mux_k_18_new_0_i_phi_fu_119_p6 = 'bx;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_0_blk_n = indices_0_full_n;
    end else begin
        indices_0_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (write_r_full_n == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_0_write = 1'b1;
    end else begin
        indices_0_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_1_blk_n = indices_1_full_n;
    end else begin
        indices_1_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (write_r_full_n == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_1_write = 1'b1;
    end else begin
        indices_1_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_2_out1_blk_n = indices_2_out1_full_n;
    end else begin
        indices_2_out1_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (write_r_full_n == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_2_out1_write = 1'b1;
    end else begin
        indices_2_out1_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_2_out_blk_n = indices_2_out_full_n;
    end else begin
        indices_2_out_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (write_r_full_n == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_2_out_write = 1'b1;
    end else begin
        indices_2_out_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (write_r_full_n == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        internal_ap_ready = 1'b1;
    end else begin
        internal_ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((start_full_n == 1'b0) & (start_once_reg == 1'b0))) begin
        real_start = 1'b0;
    end else begin
        real_start = ap_start;
    end
end

always @ (*) begin
    if (((real_start == 1'b1) & (start_once_reg == 1'b0))) begin
        start_write = 1'b1;
    end else begin
        start_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        write_r_blk_n = write_r_full_n;
    end else begin
        write_r_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (write_r_full_n == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        write_r_write = 1'b1;
    end else begin
        write_r_write = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln187_fu_160_p2 = (k_11 + 16'd1);

assign add_ln190_fu_173_p2 = (j_11 + 16'd1);

assign add_ln193_fu_186_p2 = (i_11 + 16'd1);

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

always @ (*) begin
    ap_block_state1 = ((real_start == 1'b0) | (write_r_full_n == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1));
end

assign ap_ready = internal_ap_ready;

assign icmp_ln188_fu_167_p2 = ((add_ln187_fu_160_p2 == 16'd256) ? 1'b1 : 1'b0);

assign icmp_ln191_fu_180_p2 = ((add_ln190_fu_173_p2 == 16'd28) ? 1'b1 : 1'b0);

assign icmp_ln194_fu_192_p2 = ((add_ln193_fu_186_p2 == 16'd28) ? 1'b1 : 1'b0);

assign indices_0_din = i_11;

assign indices_1_din = j_11;

assign indices_2_out1_din = k_11[12:0];

assign indices_2_out_din = k_11[7:0];

assign select_ln194_fu_198_p3 = ((icmp_ln194_fu_192_p2[0:0] == 1'b1) ? 16'd0 : add_ln193_fu_186_p2);

assign start_out = real_start;

assign write_r_din = ((k_11 == 16'd255) ? 1'b1 : 1'b0);

endmodule //td_fused_top_tdf7_get_next_ijk
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_tdf7_l2_filters_ram (addr0, ce0, q0, addr1, ce1, d1, we1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 13;
parameter MEM_SIZE = 8192;

input[AWIDTH-1:0] addr0;
input ce0;
output wire[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
input clk;

 reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];
wire [AWIDTH-1:0] addr0_t0; 
reg [AWIDTH-1:0] addr0_t1; 
reg [DWIDTH-1:0] q0_t0;
reg [DWIDTH-1:0] q0_t1;
wire [AWIDTH-1:0] addr1_t0; 
reg [AWIDTH-1:0] addr1_t1; 
wire [DWIDTH-1:0] d1_t0; 
wire we1_t0; 
reg [DWIDTH-1:0] d1_t1; 
reg we1_t1; 


assign addr0_t0 = addr0;
assign q0 = q0_t1;
assign addr1_t0 = addr1;
assign d1_t0 = d1;
assign we1_t0 = we1;

always @(posedge clk)  
begin
    if (ce0) 
    begin
        addr0_t1 <= addr0_t0; 
        q0_t1 <= q0_t0;
    end
    if (ce1) 
    begin
        addr1_t1 <= addr1_t0; 
        d1_t1 <= d1_t0;
        we1_t1 <= we1_t0;
    end
end


always @(posedge clk)  
begin 
    if (ce0) begin
        q0_t0 <= ram[addr0_t1];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1_t1) 
            ram[addr1_t1] <= d1_t1; 
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_tdf7_l2_filters(
    reset,
    clk,
    address0,
    ce0,
    q0,
    address1,
    ce1,
    we1,
    d1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd8192;
parameter AddressWidth = 32'd13;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;



td_fused_top_tdf7_l2_filters_ram td_fused_top_tdf7_l2_filters_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 )
);

endmodule

// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf7_l2_multiply50 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        intermediate_fmaps_read,
        l2_filter_data_address0,
        l2_filter_data_ce0,
        l2_filter_data_q0,
        l2_products_address0,
        l2_products_ce0,
        l2_products_we0,
        l2_products_d0,
        indices_23_dout,
        indices_23_empty_n,
        indices_23_read
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state10 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
input  [15:0] intermediate_fmaps_read;
output  [12:0] l2_filter_data_address0;
output   l2_filter_data_ce0;
input  [15:0] l2_filter_data_q0;
output  [4:0] l2_products_address0;
output   l2_products_ce0;
output   l2_products_we0;
output  [15:0] l2_products_d0;
input  [12:0] indices_23_dout;
input   indices_23_empty_n;
output   indices_23_read;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg l2_filter_data_ce0;
reg l2_products_ce0;
reg l2_products_we0;
reg indices_23_read;

reg    ap_done_reg;
  reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    indices_23_blk_n;
reg   [5:0] i_1_1_reg_106;
reg   [12:0] l2_ichan_reg_165;
wire   [5:0] add_ln20_fu_122_p2;
wire    ap_CS_fsm_pp0_stage0;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
wire    ap_block_state4_pp0_stage0_iter2;
wire    ap_block_state5_pp0_stage0_iter3;
wire    ap_block_state6_pp0_stage0_iter4;
wire    ap_block_state7_pp0_stage0_iter5;
wire    ap_block_state8_pp0_stage0_iter6;
wire    ap_block_state9_pp0_stage0_iter7;
wire    ap_block_pp0_stage0_11001;
wire   [0:0] icmp_ln20_fu_128_p2;
reg   [0:0] icmp_ln20_reg_175;
reg   [0:0] icmp_ln20_reg_175_pp0_iter1_reg;
reg   [0:0] icmp_ln20_reg_175_pp0_iter2_reg;
reg   [0:0] icmp_ln20_reg_175_pp0_iter3_reg;
reg   [0:0] icmp_ln20_reg_175_pp0_iter4_reg;
reg   [0:0] icmp_ln20_reg_175_pp0_iter5_reg;
reg   [0:0] icmp_ln20_reg_175_pp0_iter6_reg;
wire   [4:0] l2_o_fu_134_p1;
reg   [4:0] l2_o_reg_179;
reg   [4:0] l2_o_reg_179_pp0_iter1_reg;
reg   [4:0] l2_o_reg_179_pp0_iter2_reg;
reg   [4:0] l2_o_reg_179_pp0_iter3_reg;
reg   [4:0] l2_o_reg_179_pp0_iter4_reg;
reg   [4:0] l2_o_reg_179_pp0_iter5_reg;
reg   [4:0] l2_o_reg_179_pp0_iter6_reg;
wire   [15:0] grp_fu_117_p2;
reg   [15:0] mul_i_i_reg_194;
reg    ap_block_state1;
wire    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_exit_iter0_state2;
reg    ap_enable_reg_pp0_iter1;
reg    ap_enable_reg_pp0_iter2;
reg    ap_enable_reg_pp0_iter3;
reg    ap_enable_reg_pp0_iter4;
reg    ap_enable_reg_pp0_iter5;
reg    ap_enable_reg_pp0_iter6;
reg    ap_enable_reg_pp0_iter7;
wire   [63:0] zext_ln29_7_fu_151_p1;
wire    ap_block_pp0_stage0;
wire   [63:0] zext_ln29_fu_156_p1;
wire   [12:0] tmp_s_fu_138_p3;
wire   [12:0] add_ln29_fu_146_p2;
wire    ap_CS_fsm_state10;
reg   [2:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
#0 ap_enable_reg_pp0_iter4 = 1'b0;
#0 ap_enable_reg_pp0_iter5 = 1'b0;
#0 ap_enable_reg_pp0_iter6 = 1'b0;
#0 ap_enable_reg_pp0_iter7 = 1'b0;
end

td_fused_top_hmul_16ns_16ns_16_4_max_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hmul_16ns_16ns_16_4_max_dsp_1_U436(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(l2_filter_data_q0),
    .din1(intermediate_fmaps_read),
    .dout(grp_fu_117_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state10)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b1 == ap_condition_pp0_exit_iter0_state2))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            if ((1'b1 == ap_condition_pp0_exit_iter0_state2)) begin
                ap_enable_reg_pp0_iter1 <= (1'b1 ^ ap_condition_pp0_exit_iter0_state2);
            end else if ((1'b1 == 1'b1)) begin
                ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
            end
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter4 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter5 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter5 <= ap_enable_reg_pp0_iter4;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter6 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter6 <= ap_enable_reg_pp0_iter5;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter7 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter7 <= ap_enable_reg_pp0_iter6;
        end else if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter7 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        i_1_1_reg_106 <= 6'd0;
    end else if (((icmp_ln20_fu_128_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        i_1_1_reg_106 <= add_ln20_fu_122_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln20_reg_175 <= icmp_ln20_fu_128_p2;
        icmp_ln20_reg_175_pp0_iter1_reg <= icmp_ln20_reg_175;
        l2_o_reg_179_pp0_iter1_reg <= l2_o_reg_179;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        icmp_ln20_reg_175_pp0_iter2_reg <= icmp_ln20_reg_175_pp0_iter1_reg;
        icmp_ln20_reg_175_pp0_iter3_reg <= icmp_ln20_reg_175_pp0_iter2_reg;
        icmp_ln20_reg_175_pp0_iter4_reg <= icmp_ln20_reg_175_pp0_iter3_reg;
        icmp_ln20_reg_175_pp0_iter5_reg <= icmp_ln20_reg_175_pp0_iter4_reg;
        icmp_ln20_reg_175_pp0_iter6_reg <= icmp_ln20_reg_175_pp0_iter5_reg;
        l2_o_reg_179_pp0_iter2_reg <= l2_o_reg_179_pp0_iter1_reg;
        l2_o_reg_179_pp0_iter3_reg <= l2_o_reg_179_pp0_iter2_reg;
        l2_o_reg_179_pp0_iter4_reg <= l2_o_reg_179_pp0_iter3_reg;
        l2_o_reg_179_pp0_iter5_reg <= l2_o_reg_179_pp0_iter4_reg;
        l2_o_reg_179_pp0_iter6_reg <= l2_o_reg_179_pp0_iter5_reg;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state1)) begin
        l2_ichan_reg_165 <= indices_23_dout;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln20_fu_128_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        l2_o_reg_179 <= l2_o_fu_134_p1;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln20_reg_175_pp0_iter5_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        mul_i_i_reg_194 <= grp_fu_117_p2;
    end
end

always @ (*) begin
    if ((icmp_ln20_fu_128_p2 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state2 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state2 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state10)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter7 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state10)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_23_blk_n = indices_23_empty_n;
    end else begin
        indices_23_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_23_read = 1'b1;
    end else begin
        indices_23_read = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter3 == 1'b1)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1)))) begin
        l2_filter_data_ce0 = 1'b1;
    end else begin
        l2_filter_data_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter7 == 1'b1))) begin
        l2_products_ce0 = 1'b1;
    end else begin
        l2_products_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln20_reg_175_pp0_iter6_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter7 == 1'b1))) begin
        l2_products_we0 = 1'b1;
    end else begin
        l2_products_we0 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((~((icmp_ln20_fu_128_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0)) & ~((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter7 == 1'b1) & (ap_enable_reg_pp0_iter6 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if ((((icmp_ln20_fu_128_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0)) | ((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter7 == 1'b1) & (ap_enable_reg_pp0_iter6 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_state10;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state10 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln20_fu_122_p2 = (i_1_1_reg_106 + 6'd1);

assign add_ln29_fu_146_p2 = (tmp_s_fu_138_p3 + l2_ichan_reg_165);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state10 = ap_CS_fsm[32'd2];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1));
end

assign ap_block_state2_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter4 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage0_iter5 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage0_iter6 = ~(1'b1 == 1'b1);

assign ap_block_state9_pp0_stage0_iter7 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign icmp_ln20_fu_128_p2 = ((i_1_1_reg_106 == 6'd32) ? 1'b1 : 1'b0);

assign l2_filter_data_address0 = zext_ln29_7_fu_151_p1;

assign l2_o_fu_134_p1 = i_1_1_reg_106[4:0];

assign l2_products_address0 = zext_ln29_fu_156_p1;

assign l2_products_d0 = mul_i_i_reg_194;

assign tmp_s_fu_138_p3 = {{l2_o_fu_134_p1}, {8'd0}};

assign zext_ln29_7_fu_151_p1 = add_ln29_fu_146_p2;

assign zext_ln29_fu_156_p1 = l2_o_reg_179_pp0_iter6_reg;

endmodule //td_fused_top_tdf7_l2_multiply50
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_tdf7_l2_writeOutputs_149_running_sums_ram (addr0, ce0, d0, we0, addr1, ce1, q1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 5;
parameter MEM_SIZE = 32;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
input[AWIDTH-1:0] addr1;
input ce1;
output reg[DWIDTH-1:0] q1;
input clk;

 reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];

//initial begin
//    $readmemh("./td_fused_top_tdf7_l2_writeOutputs_149_running_sums_ram.dat", ram);
//end



always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[addr0] <= d0; 
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        q1 <= ram[addr1];
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_tdf7_l2_writeOutputs_149_running_sums(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    address1,
    ce1,
    q1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd32;
parameter AddressWidth = 32'd5;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
input[AddressWidth - 1:0] address1;
input ce1;
output[DataWidth - 1:0] q1;



td_fused_top_tdf7_l2_writeOutputs_149_running_sums_ram td_fused_top_tdf7_l2_writeOutputs_149_running_sums_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .q1( q1 )
);

endmodule

// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf7_l2_writeOutputs_149 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        indices_01_dout,
        indices_01_empty_n,
        indices_01_read,
        indices_12_dout,
        indices_12_empty_n,
        indices_12_read,
        write4_dout,
        write4_empty_n,
        write4_read,
        l2_partial_sums_address0,
        l2_partial_sums_ce0,
        l2_partial_sums_q0,
        out_data_address1,
        out_data_ce1,
        out_data_we1,
        out_data_d1,
        l2_adjustments_address0,
        l2_adjustments_ce0,
        l2_adjustments_q0
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state25 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
input  [4:0] indices_01_dout;
input   indices_01_empty_n;
output   indices_01_read;
input  [9:0] indices_12_dout;
input   indices_12_empty_n;
output   indices_12_read;
input  [0:0] write4_dout;
input   write4_empty_n;
output   write4_read;
output  [4:0] l2_partial_sums_address0;
output   l2_partial_sums_ce0;
input  [15:0] l2_partial_sums_q0;
output  [12:0] out_data_address1;
output   out_data_ce1;
output   out_data_we1;
output  [63:0] out_data_d1;
output  [4:0] l2_adjustments_address0;
output   l2_adjustments_ce0;
input  [47:0] l2_adjustments_q0;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg indices_01_read;
reg indices_12_read;
reg write4_read;
reg l2_partial_sums_ce0;
reg out_data_ce1;
reg out_data_we1;
reg l2_adjustments_ce0;

reg    ap_done_reg;
  reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    running_sums_ce0;
reg    running_sums_we0;
wire   [15:0] running_sums_d0;
wire   [4:0] running_sums_address1;
reg    running_sums_ce1;
wire   [15:0] running_sums_q1;
reg    indices_01_blk_n;
reg    indices_12_blk_n;
reg    write4_blk_n;
reg   [5:0] ochan_reg_206;
reg   [0:0] write4_read_reg_565;
wire   [11:0] add_ln109_fu_271_p2;
reg   [11:0] add_ln109_reg_571;
wire   [5:0] add_ln86_fu_277_p2;
wire    ap_CS_fsm_pp0_stage0;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
wire    ap_block_state4_pp0_stage0_iter2;
wire    ap_block_state5_pp0_stage0_iter3;
wire    ap_block_state6_pp0_stage0_iter4;
wire    ap_block_state7_pp0_stage0_iter5;
wire    ap_block_state8_pp0_stage0_iter6;
wire    ap_block_state9_pp0_stage0_iter7;
wire    ap_block_state10_pp0_stage0_iter8;
wire    ap_block_state11_pp0_stage0_iter9;
wire    ap_block_state12_pp0_stage0_iter10;
wire    ap_block_state13_pp0_stage0_iter11;
wire    ap_block_state14_pp0_stage0_iter12;
wire    ap_block_state15_pp0_stage0_iter13;
wire    ap_block_state16_pp0_stage0_iter14;
wire    ap_block_state17_pp0_stage0_iter15;
wire    ap_block_state18_pp0_stage0_iter16;
wire    ap_block_state19_pp0_stage0_iter17;
wire    ap_block_state20_pp0_stage0_iter18;
wire    ap_block_state21_pp0_stage0_iter19;
wire    ap_block_state22_pp0_stage0_iter20;
wire    ap_block_state23_pp0_stage0_iter21;
wire    ap_block_state24_pp0_stage0_iter22;
wire    ap_block_pp0_stage0_11001;
wire   [0:0] icmp_ln86_fu_283_p2;
wire   [63:0] zext_ln86_fu_289_p1;
reg   [63:0] zext_ln86_reg_585;
reg   [63:0] zext_ln86_reg_585_pp0_iter1_reg;
reg   [63:0] zext_ln86_reg_585_pp0_iter2_reg;
reg   [63:0] zext_ln86_reg_585_pp0_iter3_reg;
reg   [4:0] running_sums_addr_reg_595;
reg   [4:0] running_sums_addr_reg_595_pp0_iter1_reg;
reg   [4:0] running_sums_addr_reg_595_pp0_iter2_reg;
reg   [4:0] running_sums_addr_reg_595_pp0_iter3_reg;
reg   [4:0] running_sums_addr_reg_595_pp0_iter4_reg;
reg   [4:0] running_sums_addr_reg_595_pp0_iter5_reg;
reg   [4:0] running_sums_addr_reg_595_pp0_iter6_reg;
wire   [1:0] trunc_ln99_fu_295_p1;
reg   [1:0] trunc_ln99_reg_601;
reg   [1:0] trunc_ln99_reg_601_pp0_iter1_reg;
reg   [1:0] trunc_ln99_reg_601_pp0_iter2_reg;
reg   [1:0] trunc_ln99_reg_601_pp0_iter3_reg;
reg   [1:0] trunc_ln99_reg_601_pp0_iter4_reg;
reg   [1:0] trunc_ln99_reg_601_pp0_iter5_reg;
reg   [1:0] trunc_ln99_reg_601_pp0_iter6_reg;
reg   [1:0] trunc_ln99_reg_601_pp0_iter7_reg;
reg   [1:0] trunc_ln99_reg_601_pp0_iter8_reg;
reg   [1:0] trunc_ln99_reg_601_pp0_iter9_reg;
reg   [1:0] trunc_ln99_reg_601_pp0_iter10_reg;
reg   [1:0] trunc_ln99_reg_601_pp0_iter11_reg;
reg   [1:0] trunc_ln99_reg_601_pp0_iter12_reg;
reg   [1:0] trunc_ln99_reg_601_pp0_iter13_reg;
reg   [1:0] trunc_ln99_reg_601_pp0_iter14_reg;
reg   [1:0] trunc_ln99_reg_601_pp0_iter15_reg;
reg   [1:0] trunc_ln99_reg_601_pp0_iter16_reg;
reg   [1:0] trunc_ln99_reg_601_pp0_iter17_reg;
reg   [1:0] trunc_ln99_reg_601_pp0_iter18_reg;
reg   [1:0] trunc_ln99_reg_601_pp0_iter19_reg;
reg   [1:0] trunc_ln99_reg_601_pp0_iter20_reg;
wire   [0:0] and_ln103_fu_305_p2;
reg   [0:0] and_ln103_reg_608;
reg   [0:0] and_ln103_reg_608_pp0_iter1_reg;
reg   [0:0] and_ln103_reg_608_pp0_iter2_reg;
reg   [0:0] and_ln103_reg_608_pp0_iter3_reg;
reg   [0:0] and_ln103_reg_608_pp0_iter4_reg;
reg   [0:0] and_ln103_reg_608_pp0_iter5_reg;
reg   [0:0] and_ln103_reg_608_pp0_iter6_reg;
reg   [0:0] and_ln103_reg_608_pp0_iter7_reg;
reg   [0:0] and_ln103_reg_608_pp0_iter8_reg;
reg   [0:0] and_ln103_reg_608_pp0_iter9_reg;
reg   [0:0] and_ln103_reg_608_pp0_iter10_reg;
reg   [0:0] and_ln103_reg_608_pp0_iter11_reg;
reg   [0:0] and_ln103_reg_608_pp0_iter12_reg;
reg   [0:0] and_ln103_reg_608_pp0_iter13_reg;
reg   [0:0] and_ln103_reg_608_pp0_iter14_reg;
reg   [0:0] and_ln103_reg_608_pp0_iter15_reg;
reg   [0:0] and_ln103_reg_608_pp0_iter16_reg;
reg   [0:0] and_ln103_reg_608_pp0_iter17_reg;
reg   [0:0] and_ln103_reg_608_pp0_iter18_reg;
reg   [0:0] and_ln103_reg_608_pp0_iter19_reg;
reg   [0:0] and_ln103_reg_608_pp0_iter20_reg;
reg   [2:0] lshr_ln_reg_612;
reg   [2:0] lshr_ln_reg_612_pp0_iter1_reg;
reg   [2:0] lshr_ln_reg_612_pp0_iter2_reg;
reg   [2:0] lshr_ln_reg_612_pp0_iter3_reg;
reg   [2:0] lshr_ln_reg_612_pp0_iter4_reg;
reg   [2:0] lshr_ln_reg_612_pp0_iter5_reg;
reg   [2:0] lshr_ln_reg_612_pp0_iter6_reg;
reg   [2:0] lshr_ln_reg_612_pp0_iter7_reg;
reg   [2:0] lshr_ln_reg_612_pp0_iter8_reg;
reg   [2:0] lshr_ln_reg_612_pp0_iter9_reg;
reg   [2:0] lshr_ln_reg_612_pp0_iter10_reg;
reg   [2:0] lshr_ln_reg_612_pp0_iter11_reg;
reg   [2:0] lshr_ln_reg_612_pp0_iter12_reg;
reg   [2:0] lshr_ln_reg_612_pp0_iter13_reg;
reg   [2:0] lshr_ln_reg_612_pp0_iter14_reg;
reg   [2:0] lshr_ln_reg_612_pp0_iter15_reg;
reg   [2:0] lshr_ln_reg_612_pp0_iter16_reg;
reg   [2:0] lshr_ln_reg_612_pp0_iter17_reg;
reg   [2:0] lshr_ln_reg_612_pp0_iter18_reg;
reg   [2:0] lshr_ln_reg_612_pp0_iter19_reg;
reg   [2:0] lshr_ln_reg_612_pp0_iter20_reg;
reg   [15:0] val_reg_617;
reg   [15:0] running_sums_load_reg_622;
reg    ap_enable_reg_pp0_iter1;
wire   [15:0] grp_fu_217_p2;
reg   [15:0] sum_reg_632;
reg   [15:0] tmp_20_i_i_reg_643;
reg   [15:0] tmp_20_i_i_reg_643_pp0_iter8_reg;
reg   [15:0] tmp_20_i_i_reg_643_pp0_iter9_reg;
reg   [15:0] tmp_20_i_i_reg_643_pp0_iter10_reg;
reg   [15:0] tmp_20_i_i_reg_643_pp0_iter11_reg;
reg   [15:0] tmp_21_i_i_reg_648;
reg   [15:0] tmp_21_i_i_reg_648_pp0_iter8_reg;
reg   [15:0] tmp_21_i_i_reg_648_pp0_iter9_reg;
reg   [15:0] tmp_21_i_i_reg_648_pp0_iter10_reg;
reg   [15:0] tmp_21_i_i_reg_648_pp0_iter11_reg;
reg   [15:0] tmp_21_i_i_reg_648_pp0_iter12_reg;
reg   [15:0] tmp_21_i_i_reg_648_pp0_iter13_reg;
reg   [15:0] tmp_21_i_i_reg_648_pp0_iter14_reg;
reg   [15:0] tmp_21_i_i_reg_648_pp0_iter15_reg;
wire   [15:0] grp_fu_225_p2;
reg   [15:0] sub_i_i_i_reg_653;
wire   [15:0] grp_fu_229_p2;
reg   [15:0] normalized_reg_663;
wire   [15:0] grp_fu_221_p2;
reg   [15:0] biased_reg_673;
reg    ap_block_state1;
wire    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_exit_iter0_state2;
reg    ap_enable_reg_pp0_iter2;
reg    ap_enable_reg_pp0_iter3;
reg    ap_enable_reg_pp0_iter4;
reg    ap_enable_reg_pp0_iter5;
reg    ap_enable_reg_pp0_iter6;
reg    ap_enable_reg_pp0_iter7;
reg    ap_enable_reg_pp0_iter8;
reg    ap_enable_reg_pp0_iter9;
reg    ap_enable_reg_pp0_iter10;
reg    ap_enable_reg_pp0_iter11;
reg    ap_enable_reg_pp0_iter12;
reg    ap_enable_reg_pp0_iter13;
reg    ap_enable_reg_pp0_iter14;
reg    ap_enable_reg_pp0_iter15;
reg    ap_enable_reg_pp0_iter16;
reg    ap_enable_reg_pp0_iter17;
reg    ap_enable_reg_pp0_iter18;
reg    ap_enable_reg_pp0_iter19;
reg    ap_enable_reg_pp0_iter20;
reg    ap_enable_reg_pp0_iter21;
reg    ap_enable_reg_pp0_iter22;
wire    ap_block_pp0_stage0;
wire   [63:0] sext_ln109_fu_507_p1;
reg   [15:0] quad_3_1_fu_112;
wire   [15:0] quad_3_13_fu_473_p3;
reg   [15:0] quad_3_2_fu_116;
wire   [15:0] quad_3_12_fu_465_p3;
reg   [15:0] quad_3_3_fu_120;
wire   [15:0] quad_3_10_fu_449_p3;
reg   [15:0] quad_3_4_fu_124;
wire   [15:0] quad_3_7_fu_425_p3;
wire   [15:0] grp_fu_221_p1;
wire   [15:0] grp_fu_225_p1;
wire   [15:0] grp_fu_229_p1;
wire   [9:0] tmp_fu_233_p3;
wire   [6:0] tmp_s_fu_245_p3;
wire   [10:0] zext_ln109_fu_241_p1;
wire   [10:0] zext_ln109_1_fu_253_p1;
wire   [10:0] sub_ln109_fu_257_p2;
wire   [11:0] sub_ln109_cast_fu_263_p1;
wire   [11:0] zext_ln109_2_fu_267_p1;
wire   [0:0] icmp_ln103_fu_299_p2;
wire   [15:0] trunc_ln95_fu_327_p1;
wire   [15:0] data_V_fu_376_p1;
wire   [0:0] p_Result_s_fu_379_p3;
wire   [0:0] icmp_ln99_fu_394_p2;
wire   [15:0] quad_0_fu_387_p3;
wire   [0:0] icmp_ln99_1_fu_407_p2;
wire   [15:0] quad_3_fu_399_p3;
wire   [0:0] icmp_ln99_2_fu_420_p2;
wire   [15:0] quad_3_6_fu_412_p3;
wire   [15:0] quad_3_8_fu_433_p3;
wire   [15:0] quad_3_9_fu_441_p3;
wire   [15:0] quad_3_11_fu_457_p3;
wire   [14:0] tmp_17_fu_501_p3;
wire   [15:0] bitcast_ln109_3_fu_524_p1;
wire   [15:0] bitcast_ln109_2_fu_520_p1;
wire   [15:0] bitcast_ln109_1_fu_516_p1;
wire   [15:0] bitcast_ln109_fu_512_p1;
wire    ap_CS_fsm_state25;
reg   [2:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
#0 ap_enable_reg_pp0_iter4 = 1'b0;
#0 ap_enable_reg_pp0_iter5 = 1'b0;
#0 ap_enable_reg_pp0_iter6 = 1'b0;
#0 ap_enable_reg_pp0_iter7 = 1'b0;
#0 ap_enable_reg_pp0_iter8 = 1'b0;
#0 ap_enable_reg_pp0_iter9 = 1'b0;
#0 ap_enable_reg_pp0_iter10 = 1'b0;
#0 ap_enable_reg_pp0_iter11 = 1'b0;
#0 ap_enable_reg_pp0_iter12 = 1'b0;
#0 ap_enable_reg_pp0_iter13 = 1'b0;
#0 ap_enable_reg_pp0_iter14 = 1'b0;
#0 ap_enable_reg_pp0_iter15 = 1'b0;
#0 ap_enable_reg_pp0_iter16 = 1'b0;
#0 ap_enable_reg_pp0_iter17 = 1'b0;
#0 ap_enable_reg_pp0_iter18 = 1'b0;
#0 ap_enable_reg_pp0_iter19 = 1'b0;
#0 ap_enable_reg_pp0_iter20 = 1'b0;
#0 ap_enable_reg_pp0_iter21 = 1'b0;
#0 ap_enable_reg_pp0_iter22 = 1'b0;
end

td_fused_top_tdf7_l2_writeOutputs_149_running_sums #(
    .DataWidth( 16 ),
    .AddressRange( 32 ),
    .AddressWidth( 5 ))
running_sums_U(
    .reset(ap_rst),
    .clk(ap_clk),
    .address0(running_sums_addr_reg_595_pp0_iter6_reg),
    .ce0(running_sums_ce0),
    .we0(running_sums_we0),
    .d0(running_sums_d0),
    .address1(running_sums_address1),
    .ce1(running_sums_ce1),
    .q1(running_sums_q1)
);

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U441(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(running_sums_load_reg_622),
    .din1(val_reg_617),
    .dout(grp_fu_217_p2)
);

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U442(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(normalized_reg_663),
    .din1(grp_fu_221_p1),
    .dout(grp_fu_221_p2)
);

td_fused_top_hsub_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hsub_16ns_16ns_16_5_full_dsp_1_U443(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(sum_reg_632),
    .din1(grp_fu_225_p1),
    .dout(grp_fu_225_p2)
);

td_fused_top_hmul_16ns_16ns_16_4_max_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hmul_16ns_16ns_16_4_max_dsp_1_U444(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(sub_i_i_i_reg_653),
    .din1(grp_fu_229_p1),
    .dout(grp_fu_229_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state25)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b1 == ap_condition_pp0_exit_iter0_state2) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((~((ap_start == 1'b0) | (write4_empty_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            if ((1'b1 == ap_condition_pp0_exit_iter0_state2)) begin
                ap_enable_reg_pp0_iter1 <= (1'b1 ^ ap_condition_pp0_exit_iter0_state2);
            end else if ((1'b1 == 1'b1)) begin
                ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
            end
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter10 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter10 <= ap_enable_reg_pp0_iter9;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter11 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter11 <= ap_enable_reg_pp0_iter10;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter12 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter12 <= ap_enable_reg_pp0_iter11;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter13 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter13 <= ap_enable_reg_pp0_iter12;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter14 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter14 <= ap_enable_reg_pp0_iter13;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter15 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter15 <= ap_enable_reg_pp0_iter14;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter16 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter16 <= ap_enable_reg_pp0_iter15;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter17 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter17 <= ap_enable_reg_pp0_iter16;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter18 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter18 <= ap_enable_reg_pp0_iter17;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter19 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter19 <= ap_enable_reg_pp0_iter18;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter20 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter20 <= ap_enable_reg_pp0_iter19;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter21 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter21 <= ap_enable_reg_pp0_iter20;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter22 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter22 <= ap_enable_reg_pp0_iter21;
        end else if ((~((ap_start == 1'b0) | (write4_empty_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter22 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter4 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter5 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter5 <= ap_enable_reg_pp0_iter4;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter6 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter6 <= ap_enable_reg_pp0_iter5;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter7 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter7 <= ap_enable_reg_pp0_iter6;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter8 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter8 <= ap_enable_reg_pp0_iter7;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter9 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter9 <= ap_enable_reg_pp0_iter8;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (icmp_ln86_fu_283_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        ochan_reg_206 <= add_ln86_fu_277_p2;
    end else if ((~((ap_start == 1'b0) | (write4_empty_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ochan_reg_206 <= 6'd0;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state1)) begin
        add_ln109_reg_571 <= add_ln109_fu_271_p2;
        write4_read_reg_565 <= write4_dout;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (icmp_ln86_fu_283_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        and_ln103_reg_608 <= and_ln103_fu_305_p2;
        running_sums_addr_reg_595 <= zext_ln86_fu_289_p1;
        trunc_ln99_reg_601 <= trunc_ln99_fu_295_p1;
        zext_ln86_reg_585[5 : 0] <= zext_ln86_fu_289_p1[5 : 0];
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        and_ln103_reg_608_pp0_iter10_reg <= and_ln103_reg_608_pp0_iter9_reg;
        and_ln103_reg_608_pp0_iter11_reg <= and_ln103_reg_608_pp0_iter10_reg;
        and_ln103_reg_608_pp0_iter12_reg <= and_ln103_reg_608_pp0_iter11_reg;
        and_ln103_reg_608_pp0_iter13_reg <= and_ln103_reg_608_pp0_iter12_reg;
        and_ln103_reg_608_pp0_iter14_reg <= and_ln103_reg_608_pp0_iter13_reg;
        and_ln103_reg_608_pp0_iter15_reg <= and_ln103_reg_608_pp0_iter14_reg;
        and_ln103_reg_608_pp0_iter16_reg <= and_ln103_reg_608_pp0_iter15_reg;
        and_ln103_reg_608_pp0_iter17_reg <= and_ln103_reg_608_pp0_iter16_reg;
        and_ln103_reg_608_pp0_iter18_reg <= and_ln103_reg_608_pp0_iter17_reg;
        and_ln103_reg_608_pp0_iter19_reg <= and_ln103_reg_608_pp0_iter18_reg;
        and_ln103_reg_608_pp0_iter20_reg <= and_ln103_reg_608_pp0_iter19_reg;
        and_ln103_reg_608_pp0_iter2_reg <= and_ln103_reg_608_pp0_iter1_reg;
        and_ln103_reg_608_pp0_iter3_reg <= and_ln103_reg_608_pp0_iter2_reg;
        and_ln103_reg_608_pp0_iter4_reg <= and_ln103_reg_608_pp0_iter3_reg;
        and_ln103_reg_608_pp0_iter5_reg <= and_ln103_reg_608_pp0_iter4_reg;
        and_ln103_reg_608_pp0_iter6_reg <= and_ln103_reg_608_pp0_iter5_reg;
        and_ln103_reg_608_pp0_iter7_reg <= and_ln103_reg_608_pp0_iter6_reg;
        and_ln103_reg_608_pp0_iter8_reg <= and_ln103_reg_608_pp0_iter7_reg;
        and_ln103_reg_608_pp0_iter9_reg <= and_ln103_reg_608_pp0_iter8_reg;
        biased_reg_673 <= grp_fu_221_p2;
        lshr_ln_reg_612_pp0_iter10_reg <= lshr_ln_reg_612_pp0_iter9_reg;
        lshr_ln_reg_612_pp0_iter11_reg <= lshr_ln_reg_612_pp0_iter10_reg;
        lshr_ln_reg_612_pp0_iter12_reg <= lshr_ln_reg_612_pp0_iter11_reg;
        lshr_ln_reg_612_pp0_iter13_reg <= lshr_ln_reg_612_pp0_iter12_reg;
        lshr_ln_reg_612_pp0_iter14_reg <= lshr_ln_reg_612_pp0_iter13_reg;
        lshr_ln_reg_612_pp0_iter15_reg <= lshr_ln_reg_612_pp0_iter14_reg;
        lshr_ln_reg_612_pp0_iter16_reg <= lshr_ln_reg_612_pp0_iter15_reg;
        lshr_ln_reg_612_pp0_iter17_reg <= lshr_ln_reg_612_pp0_iter16_reg;
        lshr_ln_reg_612_pp0_iter18_reg <= lshr_ln_reg_612_pp0_iter17_reg;
        lshr_ln_reg_612_pp0_iter19_reg <= lshr_ln_reg_612_pp0_iter18_reg;
        lshr_ln_reg_612_pp0_iter20_reg <= lshr_ln_reg_612_pp0_iter19_reg;
        lshr_ln_reg_612_pp0_iter2_reg <= lshr_ln_reg_612_pp0_iter1_reg;
        lshr_ln_reg_612_pp0_iter3_reg <= lshr_ln_reg_612_pp0_iter2_reg;
        lshr_ln_reg_612_pp0_iter4_reg <= lshr_ln_reg_612_pp0_iter3_reg;
        lshr_ln_reg_612_pp0_iter5_reg <= lshr_ln_reg_612_pp0_iter4_reg;
        lshr_ln_reg_612_pp0_iter6_reg <= lshr_ln_reg_612_pp0_iter5_reg;
        lshr_ln_reg_612_pp0_iter7_reg <= lshr_ln_reg_612_pp0_iter6_reg;
        lshr_ln_reg_612_pp0_iter8_reg <= lshr_ln_reg_612_pp0_iter7_reg;
        lshr_ln_reg_612_pp0_iter9_reg <= lshr_ln_reg_612_pp0_iter8_reg;
        normalized_reg_663 <= grp_fu_229_p2;
        running_sums_addr_reg_595_pp0_iter2_reg <= running_sums_addr_reg_595_pp0_iter1_reg;
        running_sums_addr_reg_595_pp0_iter3_reg <= running_sums_addr_reg_595_pp0_iter2_reg;
        running_sums_addr_reg_595_pp0_iter4_reg <= running_sums_addr_reg_595_pp0_iter3_reg;
        running_sums_addr_reg_595_pp0_iter5_reg <= running_sums_addr_reg_595_pp0_iter4_reg;
        running_sums_addr_reg_595_pp0_iter6_reg <= running_sums_addr_reg_595_pp0_iter5_reg;
        sub_i_i_i_reg_653 <= grp_fu_225_p2;
        sum_reg_632 <= grp_fu_217_p2;
        tmp_20_i_i_reg_643 <= {{l2_adjustments_q0[31:16]}};
        tmp_20_i_i_reg_643_pp0_iter10_reg <= tmp_20_i_i_reg_643_pp0_iter9_reg;
        tmp_20_i_i_reg_643_pp0_iter11_reg <= tmp_20_i_i_reg_643_pp0_iter10_reg;
        tmp_20_i_i_reg_643_pp0_iter8_reg <= tmp_20_i_i_reg_643;
        tmp_20_i_i_reg_643_pp0_iter9_reg <= tmp_20_i_i_reg_643_pp0_iter8_reg;
        tmp_21_i_i_reg_648 <= {{l2_adjustments_q0[47:32]}};
        tmp_21_i_i_reg_648_pp0_iter10_reg <= tmp_21_i_i_reg_648_pp0_iter9_reg;
        tmp_21_i_i_reg_648_pp0_iter11_reg <= tmp_21_i_i_reg_648_pp0_iter10_reg;
        tmp_21_i_i_reg_648_pp0_iter12_reg <= tmp_21_i_i_reg_648_pp0_iter11_reg;
        tmp_21_i_i_reg_648_pp0_iter13_reg <= tmp_21_i_i_reg_648_pp0_iter12_reg;
        tmp_21_i_i_reg_648_pp0_iter14_reg <= tmp_21_i_i_reg_648_pp0_iter13_reg;
        tmp_21_i_i_reg_648_pp0_iter15_reg <= tmp_21_i_i_reg_648_pp0_iter14_reg;
        tmp_21_i_i_reg_648_pp0_iter8_reg <= tmp_21_i_i_reg_648;
        tmp_21_i_i_reg_648_pp0_iter9_reg <= tmp_21_i_i_reg_648_pp0_iter8_reg;
        trunc_ln99_reg_601_pp0_iter10_reg <= trunc_ln99_reg_601_pp0_iter9_reg;
        trunc_ln99_reg_601_pp0_iter11_reg <= trunc_ln99_reg_601_pp0_iter10_reg;
        trunc_ln99_reg_601_pp0_iter12_reg <= trunc_ln99_reg_601_pp0_iter11_reg;
        trunc_ln99_reg_601_pp0_iter13_reg <= trunc_ln99_reg_601_pp0_iter12_reg;
        trunc_ln99_reg_601_pp0_iter14_reg <= trunc_ln99_reg_601_pp0_iter13_reg;
        trunc_ln99_reg_601_pp0_iter15_reg <= trunc_ln99_reg_601_pp0_iter14_reg;
        trunc_ln99_reg_601_pp0_iter16_reg <= trunc_ln99_reg_601_pp0_iter15_reg;
        trunc_ln99_reg_601_pp0_iter17_reg <= trunc_ln99_reg_601_pp0_iter16_reg;
        trunc_ln99_reg_601_pp0_iter18_reg <= trunc_ln99_reg_601_pp0_iter17_reg;
        trunc_ln99_reg_601_pp0_iter19_reg <= trunc_ln99_reg_601_pp0_iter18_reg;
        trunc_ln99_reg_601_pp0_iter20_reg <= trunc_ln99_reg_601_pp0_iter19_reg;
        trunc_ln99_reg_601_pp0_iter2_reg <= trunc_ln99_reg_601_pp0_iter1_reg;
        trunc_ln99_reg_601_pp0_iter3_reg <= trunc_ln99_reg_601_pp0_iter2_reg;
        trunc_ln99_reg_601_pp0_iter4_reg <= trunc_ln99_reg_601_pp0_iter3_reg;
        trunc_ln99_reg_601_pp0_iter5_reg <= trunc_ln99_reg_601_pp0_iter4_reg;
        trunc_ln99_reg_601_pp0_iter6_reg <= trunc_ln99_reg_601_pp0_iter5_reg;
        trunc_ln99_reg_601_pp0_iter7_reg <= trunc_ln99_reg_601_pp0_iter6_reg;
        trunc_ln99_reg_601_pp0_iter8_reg <= trunc_ln99_reg_601_pp0_iter7_reg;
        trunc_ln99_reg_601_pp0_iter9_reg <= trunc_ln99_reg_601_pp0_iter8_reg;
        zext_ln86_reg_585_pp0_iter2_reg[5 : 0] <= zext_ln86_reg_585_pp0_iter1_reg[5 : 0];
        zext_ln86_reg_585_pp0_iter3_reg[5 : 0] <= zext_ln86_reg_585_pp0_iter2_reg[5 : 0];
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        and_ln103_reg_608_pp0_iter1_reg <= and_ln103_reg_608;
        lshr_ln_reg_612_pp0_iter1_reg <= lshr_ln_reg_612;
        running_sums_addr_reg_595_pp0_iter1_reg <= running_sums_addr_reg_595;
        trunc_ln99_reg_601_pp0_iter1_reg <= trunc_ln99_reg_601;
        val_reg_617 <= l2_partial_sums_q0;
        zext_ln86_reg_585_pp0_iter1_reg[5 : 0] <= zext_ln86_reg_585[5 : 0];
    end
end

always @ (posedge ap_clk) begin
    if (((1'd1 == and_ln103_fu_305_p2) & (1'b1 == ap_CS_fsm_pp0_stage0) & (icmp_ln86_fu_283_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        lshr_ln_reg_612 <= {{ochan_reg_206[4:2]}};
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        quad_3_1_fu_112 <= quad_3_13_fu_473_p3;
        quad_3_2_fu_116 <= quad_3_12_fu_465_p3;
        quad_3_3_fu_120 <= quad_3_10_fu_449_p3;
        quad_3_4_fu_124 <= quad_3_7_fu_425_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        running_sums_load_reg_622 <= running_sums_q1;
    end
end

always @ (*) begin
    if ((icmp_ln86_fu_283_p2 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state2 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state2 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state25)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter22 == 1'b0) & (ap_enable_reg_pp0_iter21 == 1'b0) & (ap_enable_reg_pp0_iter20 == 1'b0) & (ap_enable_reg_pp0_iter19 == 1'b0) & (ap_enable_reg_pp0_iter18 == 1'b0) & (ap_enable_reg_pp0_iter17 == 1'b0) & (ap_enable_reg_pp0_iter16 == 1'b0) & (ap_enable_reg_pp0_iter15 == 1'b0) & (ap_enable_reg_pp0_iter14 == 1'b0) & (ap_enable_reg_pp0_iter13 == 1'b0) & (ap_enable_reg_pp0_iter12 == 1'b0) & (ap_enable_reg_pp0_iter11 == 1'b0) & (ap_enable_reg_pp0_iter10 == 1'b0) & (ap_enable_reg_pp0_iter9 == 1'b0) & (ap_enable_reg_pp0_iter8 == 1'b0) & (ap_enable_reg_pp0_iter7 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state25)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_01_blk_n = indices_01_empty_n;
    end else begin
        indices_01_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (write4_empty_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_01_read = 1'b1;
    end else begin
        indices_01_read = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_12_blk_n = indices_12_empty_n;
    end else begin
        indices_12_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (write4_empty_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_12_read = 1'b1;
    end else begin
        indices_12_read = 1'b0;
    end
end

always @ (*) begin
    if ((((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001)) | ((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001)) | ((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001)) | ((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
        l2_adjustments_ce0 = 1'b1;
    end else begin
        l2_adjustments_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        l2_partial_sums_ce0 = 1'b1;
    end else begin
        l2_partial_sums_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((((ap_enable_reg_pp0_iter22 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001)) | ((ap_enable_reg_pp0_iter21 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
        out_data_ce1 = 1'b1;
    end else begin
        out_data_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter21 == 1'b1) & (1'd1 == and_ln103_reg_608_pp0_iter20_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        out_data_we1 = 1'b1;
    end else begin
        out_data_we1 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        running_sums_ce0 = 1'b1;
    end else begin
        running_sums_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        running_sums_ce1 = 1'b1;
    end else begin
        running_sums_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        running_sums_we0 = 1'b1;
    end else begin
        running_sums_we0 = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        write4_blk_n = write4_empty_n;
    end else begin
        write4_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (write4_empty_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        write4_read = 1'b1;
    end else begin
        write4_read = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_start == 1'b0) | (write4_empty_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((~((ap_enable_reg_pp0_iter0 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0) & (icmp_ln86_fu_283_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone)) & ~((ap_enable_reg_pp0_iter22 == 1'b1) & (ap_enable_reg_pp0_iter21 == 1'b0) & (1'b0 == ap_block_pp0_stage0_subdone)))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0) & (icmp_ln86_fu_283_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone)) | ((ap_enable_reg_pp0_iter22 == 1'b1) & (ap_enable_reg_pp0_iter21 == 1'b0) & (1'b0 == ap_block_pp0_stage0_subdone)))) begin
                ap_NS_fsm = ap_ST_fsm_state25;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state25 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln109_fu_271_p2 = ((sub_ln109_cast_fu_263_p1) + (zext_ln109_2_fu_267_p1));

assign add_ln86_fu_277_p2 = (ochan_reg_206 + 6'd1);

assign and_ln103_fu_305_p2 = (write4_read_reg_565 & icmp_ln103_fu_299_p2);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state25 = ap_CS_fsm[32'd2];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (write4_empty_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1));
end

assign ap_block_state10_pp0_stage0_iter8 = ~(1'b1 == 1'b1);

assign ap_block_state11_pp0_stage0_iter9 = ~(1'b1 == 1'b1);

assign ap_block_state12_pp0_stage0_iter10 = ~(1'b1 == 1'b1);

assign ap_block_state13_pp0_stage0_iter11 = ~(1'b1 == 1'b1);

assign ap_block_state14_pp0_stage0_iter12 = ~(1'b1 == 1'b1);

assign ap_block_state15_pp0_stage0_iter13 = ~(1'b1 == 1'b1);

assign ap_block_state16_pp0_stage0_iter14 = ~(1'b1 == 1'b1);

assign ap_block_state17_pp0_stage0_iter15 = ~(1'b1 == 1'b1);

assign ap_block_state18_pp0_stage0_iter16 = ~(1'b1 == 1'b1);

assign ap_block_state19_pp0_stage0_iter17 = ~(1'b1 == 1'b1);

assign ap_block_state20_pp0_stage0_iter18 = ~(1'b1 == 1'b1);

assign ap_block_state21_pp0_stage0_iter19 = ~(1'b1 == 1'b1);

assign ap_block_state22_pp0_stage0_iter20 = ~(1'b1 == 1'b1);

assign ap_block_state23_pp0_stage0_iter21 = ~(1'b1 == 1'b1);

assign ap_block_state24_pp0_stage0_iter22 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter4 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage0_iter5 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage0_iter6 = ~(1'b1 == 1'b1);

assign ap_block_state9_pp0_stage0_iter7 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign bitcast_ln109_1_fu_516_p1 = quad_3_12_fu_465_p3;

assign bitcast_ln109_2_fu_520_p1 = quad_3_10_fu_449_p3;

assign bitcast_ln109_3_fu_524_p1 = quad_3_7_fu_425_p3;

assign bitcast_ln109_fu_512_p1 = quad_3_13_fu_473_p3;

assign data_V_fu_376_p1 = biased_reg_673;

assign grp_fu_221_p1 = tmp_21_i_i_reg_648_pp0_iter15_reg;

assign grp_fu_225_p1 = trunc_ln95_fu_327_p1;

assign grp_fu_229_p1 = tmp_20_i_i_reg_643_pp0_iter11_reg;

assign icmp_ln103_fu_299_p2 = ((trunc_ln99_fu_295_p1 == 2'd3) ? 1'b1 : 1'b0);

assign icmp_ln86_fu_283_p2 = ((ochan_reg_206 == 6'd32) ? 1'b1 : 1'b0);

assign icmp_ln99_1_fu_407_p2 = ((trunc_ln99_reg_601_pp0_iter20_reg == 2'd1) ? 1'b1 : 1'b0);

assign icmp_ln99_2_fu_420_p2 = ((trunc_ln99_reg_601_pp0_iter20_reg == 2'd0) ? 1'b1 : 1'b0);

assign icmp_ln99_fu_394_p2 = ((trunc_ln99_reg_601_pp0_iter20_reg == 2'd2) ? 1'b1 : 1'b0);

assign l2_adjustments_address0 = zext_ln86_reg_585_pp0_iter3_reg;

assign l2_partial_sums_address0 = zext_ln86_fu_289_p1;

assign out_data_address1 = sext_ln109_fu_507_p1;

assign out_data_d1 = {{{{bitcast_ln109_3_fu_524_p1}, {bitcast_ln109_2_fu_520_p1}}, {bitcast_ln109_1_fu_516_p1}}, {bitcast_ln109_fu_512_p1}};

assign p_Result_s_fu_379_p3 = data_V_fu_376_p1[32'd15];

assign quad_0_fu_387_p3 = ((p_Result_s_fu_379_p3[0:0] == 1'b1) ? 16'd0 : biased_reg_673);

assign quad_3_10_fu_449_p3 = ((icmp_ln99_2_fu_420_p2[0:0] == 1'b1) ? quad_3_3_fu_120 : quad_3_9_fu_441_p3);

assign quad_3_11_fu_457_p3 = ((icmp_ln99_1_fu_407_p2[0:0] == 1'b1) ? quad_0_fu_387_p3 : quad_3_2_fu_116);

assign quad_3_12_fu_465_p3 = ((icmp_ln99_2_fu_420_p2[0:0] == 1'b1) ? quad_3_2_fu_116 : quad_3_11_fu_457_p3);

assign quad_3_13_fu_473_p3 = ((icmp_ln99_2_fu_420_p2[0:0] == 1'b1) ? quad_0_fu_387_p3 : quad_3_1_fu_112);

assign quad_3_6_fu_412_p3 = ((icmp_ln99_1_fu_407_p2[0:0] == 1'b1) ? quad_3_4_fu_124 : quad_3_fu_399_p3);

assign quad_3_7_fu_425_p3 = ((icmp_ln99_2_fu_420_p2[0:0] == 1'b1) ? quad_3_4_fu_124 : quad_3_6_fu_412_p3);

assign quad_3_8_fu_433_p3 = ((icmp_ln99_fu_394_p2[0:0] == 1'b1) ? quad_0_fu_387_p3 : quad_3_3_fu_120);

assign quad_3_9_fu_441_p3 = ((icmp_ln99_1_fu_407_p2[0:0] == 1'b1) ? quad_3_3_fu_120 : quad_3_8_fu_433_p3);

assign quad_3_fu_399_p3 = ((icmp_ln99_fu_394_p2[0:0] == 1'b1) ? quad_3_4_fu_124 : quad_0_fu_387_p3);

assign running_sums_address1 = zext_ln86_fu_289_p1;

assign running_sums_d0 = ((write4_read_reg_565[0:0] == 1'b1) ? 16'd0 : sum_reg_632);

assign sext_ln109_fu_507_p1 = (tmp_17_fu_501_p3);

assign sub_ln109_cast_fu_263_p1 = (sub_ln109_fu_257_p2);

assign sub_ln109_fu_257_p2 = (zext_ln109_fu_241_p1 - zext_ln109_1_fu_253_p1);

assign tmp_17_fu_501_p3 = {{add_ln109_reg_571}, {lshr_ln_reg_612_pp0_iter20_reg}};

assign tmp_fu_233_p3 = {{indices_01_dout}, {5'd0}};

assign tmp_s_fu_245_p3 = {{indices_01_dout}, {2'd0}};

assign trunc_ln95_fu_327_p1 = l2_adjustments_q0[15:0];

assign trunc_ln99_fu_295_p1 = ochan_reg_206[1:0];

assign zext_ln109_1_fu_253_p1 = tmp_s_fu_245_p3;

assign zext_ln109_2_fu_267_p1 = indices_12_dout;

assign zext_ln109_fu_241_p1 = tmp_fu_233_p3;

assign zext_ln86_fu_289_p1 = ochan_reg_206;

always @ (posedge ap_clk) begin
    zext_ln86_reg_585[63:6] <= 58'b0000000000000000000000000000000000000000000000000000000000;
    zext_ln86_reg_585_pp0_iter1_reg[63:6] <= 58'b0000000000000000000000000000000000000000000000000000000000;
    zext_ln86_reg_585_pp0_iter2_reg[63:6] <= 58'b0000000000000000000000000000000000000000000000000000000000;
    zext_ln86_reg_585_pp0_iter3_reg[63:6] <= 58'b0000000000000000000000000000000000000000000000000000000000;
end

endmodule //td_fused_top_tdf7_l2_writeOutputs_149
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf7_readFilters52 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        filter_data_address0,
        filter_data_ce0,
        filter_data_q0,
        indices_23_dout,
        indices_23_empty_n,
        indices_23_read,
        weight_vecs_0_address0,
        weight_vecs_0_ce0,
        weight_vecs_0_we0,
        weight_vecs_0_d0
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state7 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [16:0] filter_data_address0;
output   filter_data_ce0;
input  [15:0] filter_data_q0;
input  [7:0] indices_23_dout;
input   indices_23_empty_n;
output   indices_23_read;
output  [8:0] weight_vecs_0_address0;
output   weight_vecs_0_ce0;
output   weight_vecs_0_we0;
output  [15:0] weight_vecs_0_d0;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg filter_data_ce0;
reg indices_23_read;
reg weight_vecs_0_ce0;
reg weight_vecs_0_we0;

reg    ap_done_reg;
  reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    indices_23_blk_n;
reg   [8:0] indvar_flatten13_reg_123;
reg   [1:0] ii_reg_134;
reg   [7:0] indvar_flatten_reg_145;
reg   [1:0] jj_reg_156;
reg   [5:0] kk_reg_167;
wire   [11:0] sext_ln47_fu_200_p1;
reg   [11:0] sext_ln47_reg_408;
wire   [8:0] add_ln47_2_fu_204_p2;
wire    ap_CS_fsm_pp0_stage0;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
wire    ap_block_state4_pp0_stage0_iter2;
wire    ap_block_state5_pp0_stage0_iter3;
wire    ap_block_state6_pp0_stage0_iter4;
wire    ap_block_pp0_stage0_11001;
wire   [0:0] icmp_ln47_fu_210_p2;
reg   [0:0] icmp_ln47_reg_418;
reg   [0:0] icmp_ln47_reg_418_pp0_iter1_reg;
reg   [0:0] icmp_ln47_reg_418_pp0_iter2_reg;
reg   [0:0] icmp_ln47_reg_418_pp0_iter3_reg;
wire   [0:0] icmp_ln48_fu_222_p2;
reg   [0:0] icmp_ln48_reg_422;
wire   [1:0] select_ln47_2_fu_228_p3;
reg   [1:0] select_ln47_2_reg_429;
wire   [7:0] select_ln48_4_fu_242_p3;
wire   [1:0] select_ln48_3_fu_329_p3;
reg   [1:0] select_ln48_3_reg_442;
reg    ap_enable_reg_pp0_iter1;
wire   [8:0] add_ln55_8_fu_392_p2;
reg   [8:0] add_ln55_8_reg_452;
reg   [8:0] add_ln55_8_reg_452_pp0_iter2_reg;
reg   [8:0] add_ln55_8_reg_452_pp0_iter3_reg;
wire   [5:0] add_ln49_fu_398_p2;
reg    ap_block_state1;
wire    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_flush_enable;
reg    ap_enable_reg_pp0_iter2;
reg    ap_condition_pp0_exit_iter1_state3;
reg    ap_enable_reg_pp0_iter3;
reg    ap_enable_reg_pp0_iter4;
reg   [1:0] ap_phi_mux_ii_phi_fu_138_p4;
wire    ap_block_pp0_stage0;
reg   [1:0] ap_phi_mux_jj_phi_fu_160_p4;
wire   [63:0] zext_ln55_18_fu_387_p1;
wire   [63:0] zext_ln55_19_fu_404_p1;
wire   [9:0] tmp_fu_182_p3;
wire   [10:0] zext_ln55_11_fu_190_p1;
wire   [10:0] zext_ln55_fu_178_p1;
wire   [10:0] sub_ln55_fu_194_p2;
wire   [1:0] add_ln47_fu_216_p2;
wire   [7:0] add_ln48_2_fu_236_p2;
wire   [11:0] zext_ln55_13_fu_260_p1;
wire   [11:0] add_ln55_fu_263_p2;
wire   [11:0] shl_ln55_fu_268_p2;
wire   [3:0] tmp_s_fu_280_p3;
wire   [3:0] zext_ln55_12_fu_257_p1;
wire   [0:0] icmp_ln49_fu_298_p2;
wire   [0:0] xor_ln47_fu_293_p2;
wire   [1:0] select_ln47_fu_250_p3;
wire   [0:0] and_ln47_fu_304_p2;
wire   [0:0] or_ln48_fu_316_p2;
wire   [1:0] add_ln48_fu_310_p2;
wire   [11:0] sub_ln55_3_fu_274_p2;
wire   [11:0] zext_ln55_15_fu_341_p1;
wire   [11:0] add_ln55_5_fu_345_p2;
wire   [3:0] sub_ln55_4_fu_287_p2;
wire   [3:0] zext_ln55_14_fu_337_p1;
wire   [3:0] add_ln55_6_fu_359_p2;
wire   [5:0] select_ln48_fu_321_p3;
wire   [16:0] tmp_41_cast_fu_351_p3;
wire   [16:0] zext_ln55_17_fu_377_p1;
wire   [16:0] add_ln55_7_fu_381_p2;
wire   [8:0] tmp_43_cast_fu_365_p3;
wire   [8:0] zext_ln55_16_fu_373_p1;
wire    ap_CS_fsm_state7;
reg   [2:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
#0 ap_enable_reg_pp0_iter4 = 1'b0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state7)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if ((1'b1 == ap_condition_pp0_flush_enable)) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            if ((1'b1 == ap_condition_pp0_exit_iter1_state3)) begin
                ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter0;
            end else if ((1'b1 == 1'b1)) begin
                ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
            end
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter4 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
        end else if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter4 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln47_reg_418 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ii_reg_134 <= select_ln47_2_reg_429;
    end else if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ii_reg_134 <= 2'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_fu_210_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        indvar_flatten13_reg_123 <= add_ln47_2_fu_204_p2;
    end else if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indvar_flatten13_reg_123 <= 9'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_fu_210_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        indvar_flatten_reg_145 <= select_ln48_4_fu_242_p3;
    end else if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indvar_flatten_reg_145 <= 8'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_reg_418_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        jj_reg_156 <= select_ln48_3_reg_442;
    end else if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        jj_reg_156 <= 2'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln47_reg_418 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        kk_reg_167 <= add_ln49_fu_398_p2;
    end else if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        kk_reg_167 <= 6'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_reg_418 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        add_ln55_8_reg_452 <= add_ln55_8_fu_392_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        add_ln55_8_reg_452_pp0_iter2_reg <= add_ln55_8_reg_452;
        add_ln55_8_reg_452_pp0_iter3_reg <= add_ln55_8_reg_452_pp0_iter2_reg;
        icmp_ln47_reg_418_pp0_iter2_reg <= icmp_ln47_reg_418_pp0_iter1_reg;
        icmp_ln47_reg_418_pp0_iter3_reg <= icmp_ln47_reg_418_pp0_iter2_reg;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln47_reg_418 <= icmp_ln47_fu_210_p2;
        icmp_ln47_reg_418_pp0_iter1_reg <= icmp_ln47_reg_418;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_fu_210_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln48_reg_422 <= icmp_ln48_fu_222_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_fu_210_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        select_ln47_2_reg_429 <= select_ln47_2_fu_228_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln47_reg_418 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        select_ln48_3_reg_442 <= select_ln48_3_fu_329_p3;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state1)) begin
        sext_ln47_reg_408 <= sext_ln47_fu_200_p1;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_condition_pp0_exit_iter1_state3 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter1_state3 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln47_fu_210_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_condition_pp0_flush_enable = 1'b1;
    end else begin
        ap_condition_pp0_flush_enable = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state7)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln47_reg_418 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_phi_mux_ii_phi_fu_138_p4 = select_ln47_2_reg_429;
    end else begin
        ap_phi_mux_ii_phi_fu_138_p4 = ii_reg_134;
    end
end

always @ (*) begin
    if (((icmp_ln47_reg_418_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        ap_phi_mux_jj_phi_fu_160_p4 = select_ln48_3_reg_442;
    end else begin
        ap_phi_mux_jj_phi_fu_160_p4 = jj_reg_156;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state7)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter3 == 1'b1)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter4 == 1'b1)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1)))) begin
        filter_data_ce0 = 1'b1;
    end else begin
        filter_data_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_23_blk_n = indices_23_empty_n;
    end else begin
        indices_23_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_23_read = 1'b1;
    end else begin
        indices_23_read = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter4 == 1'b1))) begin
        weight_vecs_0_ce0 = 1'b1;
    end else begin
        weight_vecs_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln47_reg_418_pp0_iter3_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter4 == 1'b1))) begin
        weight_vecs_0_we0 = 1'b1;
    end else begin
        weight_vecs_0_we0 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((~((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b0)) & ~((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter4 == 1'b1) & (ap_enable_reg_pp0_iter3 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if ((((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b0)) | ((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter4 == 1'b1) & (ap_enable_reg_pp0_iter3 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_state7;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state7 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln47_2_fu_204_p2 = (indvar_flatten13_reg_123 + 9'd1);

assign add_ln47_fu_216_p2 = (ap_phi_mux_ii_phi_fu_138_p4 + 2'd1);

assign add_ln48_2_fu_236_p2 = (indvar_flatten_reg_145 + 8'd1);

assign add_ln48_fu_310_p2 = (select_ln47_fu_250_p3 + 2'd1);

assign add_ln49_fu_398_p2 = (select_ln48_fu_321_p3 + 6'd1);

assign add_ln55_5_fu_345_p2 = (sub_ln55_3_fu_274_p2 + zext_ln55_15_fu_341_p1);

assign add_ln55_6_fu_359_p2 = (sub_ln55_4_fu_287_p2 + zext_ln55_14_fu_337_p1);

assign add_ln55_7_fu_381_p2 = (tmp_41_cast_fu_351_p3 + zext_ln55_17_fu_377_p1);

assign add_ln55_8_fu_392_p2 = (tmp_43_cast_fu_365_p3 + zext_ln55_16_fu_373_p1);

assign add_ln55_fu_263_p2 = ((sext_ln47_reg_408) + (zext_ln55_13_fu_260_p1));

assign and_ln47_fu_304_p2 = (xor_ln47_fu_293_p2 & icmp_ln49_fu_298_p2);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state7 = ap_CS_fsm[32'd2];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1));
end

assign ap_block_state2_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter4 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign filter_data_address0 = zext_ln55_18_fu_387_p1;

assign icmp_ln47_fu_210_p2 = ((indvar_flatten13_reg_123 == 9'd288) ? 1'b1 : 1'b0);

assign icmp_ln48_fu_222_p2 = ((indvar_flatten_reg_145 == 8'd96) ? 1'b1 : 1'b0);

assign icmp_ln49_fu_298_p2 = ((kk_reg_167 == 6'd32) ? 1'b1 : 1'b0);

assign or_ln48_fu_316_p2 = (icmp_ln48_reg_422 | and_ln47_fu_304_p2);

assign select_ln47_2_fu_228_p3 = ((icmp_ln48_fu_222_p2[0:0] == 1'b1) ? add_ln47_fu_216_p2 : ap_phi_mux_ii_phi_fu_138_p4);

assign select_ln47_fu_250_p3 = ((icmp_ln48_reg_422[0:0] == 1'b1) ? 2'd0 : ap_phi_mux_jj_phi_fu_160_p4);

assign select_ln48_3_fu_329_p3 = ((and_ln47_fu_304_p2[0:0] == 1'b1) ? add_ln48_fu_310_p2 : select_ln47_fu_250_p3);

assign select_ln48_4_fu_242_p3 = ((icmp_ln48_fu_222_p2[0:0] == 1'b1) ? 8'd1 : add_ln48_2_fu_236_p2);

assign select_ln48_fu_321_p3 = ((or_ln48_fu_316_p2[0:0] == 1'b1) ? 6'd0 : kk_reg_167);

assign sext_ln47_fu_200_p1 = (sub_ln55_fu_194_p2);

assign shl_ln55_fu_268_p2 = add_ln55_fu_263_p2 << 12'd2;

assign sub_ln55_3_fu_274_p2 = (shl_ln55_fu_268_p2 - add_ln55_fu_263_p2);

assign sub_ln55_4_fu_287_p2 = (tmp_s_fu_280_p3 - zext_ln55_12_fu_257_p1);

assign sub_ln55_fu_194_p2 = (zext_ln55_11_fu_190_p1 - zext_ln55_fu_178_p1);

assign tmp_41_cast_fu_351_p3 = {{add_ln55_5_fu_345_p2}, {5'd0}};

assign tmp_43_cast_fu_365_p3 = {{add_ln55_6_fu_359_p2}, {5'd0}};

assign tmp_fu_182_p3 = {{indices_23_dout}, {2'd0}};

assign tmp_s_fu_280_p3 = {{select_ln47_2_reg_429}, {2'd0}};

assign weight_vecs_0_address0 = zext_ln55_19_fu_404_p1;

assign weight_vecs_0_d0 = filter_data_q0;

assign xor_ln47_fu_293_p2 = (icmp_ln48_reg_422 ^ 1'd1);

assign zext_ln55_11_fu_190_p1 = tmp_fu_182_p3;

assign zext_ln55_12_fu_257_p1 = select_ln47_2_reg_429;

assign zext_ln55_13_fu_260_p1 = select_ln47_2_reg_429;

assign zext_ln55_14_fu_337_p1 = select_ln48_3_fu_329_p3;

assign zext_ln55_15_fu_341_p1 = select_ln48_3_fu_329_p3;

assign zext_ln55_16_fu_373_p1 = select_ln48_fu_321_p3;

assign zext_ln55_17_fu_377_p1 = select_ln48_fu_321_p3;

assign zext_ln55_18_fu_387_p1 = add_ln55_7_fu_381_p2;

assign zext_ln55_19_fu_404_p1 = add_ln55_8_reg_452_pp0_iter3_reg;

assign zext_ln55_fu_178_p1 = indices_23_dout;

endmodule //td_fused_top_tdf7_readFilters52
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf7_readInputs53 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        in_data_address0,
        in_data_ce0,
        in_data_q0,
        indices_01_dout,
        indices_01_empty_n,
        indices_01_read,
        indices_12_dout,
        indices_12_empty_n,
        indices_12_read,
        ifmap_vec_address0,
        ifmap_vec_ce0,
        ifmap_vec_we0,
        ifmap_vec_d0,
        ifmap_vec_address1,
        ifmap_vec_ce1,
        ifmap_vec_we1,
        ifmap_vec_d1,
        indices_01_out_din,
        indices_01_out_full_n,
        indices_01_out_write,
        indices_12_out_din,
        indices_12_out_full_n,
        indices_12_out_write
);

parameter    ap_ST_fsm_state1 = 5'd1;
parameter    ap_ST_fsm_state2 = 5'd2;
parameter    ap_ST_fsm_pp0_stage0 = 5'd4;
parameter    ap_ST_fsm_pp0_stage1 = 5'd8;
parameter    ap_ST_fsm_state9 = 5'd16;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [12:0] in_data_address0;
output   in_data_ce0;
input  [63:0] in_data_q0;
input  [15:0] indices_01_dout;
input   indices_01_empty_n;
output   indices_01_read;
input  [15:0] indices_12_dout;
input   indices_12_empty_n;
output   indices_12_read;
output  [8:0] ifmap_vec_address0;
output   ifmap_vec_ce0;
output   ifmap_vec_we0;
output  [15:0] ifmap_vec_d0;
output  [8:0] ifmap_vec_address1;
output   ifmap_vec_ce1;
output   ifmap_vec_we1;
output  [15:0] ifmap_vec_d1;
output  [4:0] indices_01_out_din;
input   indices_01_out_full_n;
output   indices_01_out_write;
output  [9:0] indices_12_out_din;
input   indices_12_out_full_n;
output   indices_12_out_write;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg in_data_ce0;
reg indices_01_read;
reg indices_12_read;
reg[8:0] ifmap_vec_address0;
reg ifmap_vec_ce0;
reg ifmap_vec_we0;
reg[15:0] ifmap_vec_d0;
reg[8:0] ifmap_vec_address1;
reg ifmap_vec_ce1;
reg ifmap_vec_we1;
reg[15:0] ifmap_vec_d1;
reg indices_01_out_write;
reg indices_12_out_write;

reg    ap_done_reg;
  reg   [4:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    indices_01_blk_n;
reg    indices_12_blk_n;
reg    indices_01_out_blk_n;
reg    indices_12_out_blk_n;
reg   [6:0] indvar_flatten47_reg_222;
reg   [1:0] ii_reg_234;
reg   [5:0] indvar_flatten_reg_246;
reg   [1:0] jj_reg_257;
reg   [5:0] kk_0_i_i_reg_269;
reg   [15:0] indices_01_read_reg_957;
wire   [4:0] trunc_ln250_fu_280_p1;
reg   [4:0] trunc_ln250_reg_962;
reg   [15:0] indices_12_read_reg_967;
wire   [9:0] empty_fu_285_p1;
reg   [9:0] empty_reg_972;
wire   [17:0] p_cast_i_i_fu_302_p1;
reg   [17:0] p_cast_i_i_reg_979;
wire    ap_CS_fsm_state2;
wire   [17:0] sext_ln22_fu_312_p1;
reg   [17:0] sext_ln22_reg_985;
wire   [4:0] p_cast_fu_316_p2;
reg   [4:0] p_cast_reg_991;
wire   [0:0] or_ln23_6_fu_335_p2;
reg   [0:0] or_ln23_6_reg_997;
wire   [9:0] p_mid137_fu_341_p2;
reg   [9:0] p_mid137_reg_1002;
wire   [4:0] p_cast5_i_i_fu_359_p2;
reg   [4:0] p_cast5_i_i_reg_1007;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_block_state3_pp0_stage0_iter0;
wire    ap_block_state5_pp0_stage0_iter1;
wire    ap_block_state7_pp0_stage0_iter2;
wire    ap_block_pp0_stage0_11001;
wire   [0:0] is_padding_fu_399_p2;
reg   [0:0] is_padding_reg_1013;
wire   [0:0] icmp_ln19_fu_405_p2;
reg   [0:0] icmp_ln19_reg_1020;
reg   [0:0] icmp_ln19_reg_1020_pp0_iter1_reg;
reg   [0:0] icmp_ln19_reg_1020_pp0_iter2_reg;
wire   [1:0] add_ln19_fu_411_p2;
reg   [1:0] add_ln19_reg_1024;
wire   [0:0] icmp_ln20_fu_417_p2;
reg   [0:0] icmp_ln20_reg_1029;
wire   [1:0] select_ln19_fu_423_p3;
reg   [1:0] select_ln19_reg_1041;
wire   [4:0] p_cast5_i_i_mid1_fu_444_p2;
reg   [4:0] p_cast5_i_i_mid1_reg_1046;
wire   [0:0] or_ln23_8_fu_463_p2;
reg   [0:0] or_ln23_8_reg_1052;
wire   [1:0] add_ln20_fu_468_p2;
reg   [1:0] add_ln20_reg_1059;
wire   [0:0] or_ln23_10_fu_503_p2;
reg   [0:0] or_ln23_10_reg_1065;
wire   [5:0] add_ln20_2_fu_509_p2;
reg   [5:0] add_ln20_2_reg_1072;
wire   [6:0] add_ln19_2_fu_515_p2;
reg   [6:0] add_ln19_2_reg_1077;
wire    ap_CS_fsm_pp0_stage1;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_state4_pp0_stage1_iter0;
wire    ap_block_state6_pp0_stage1_iter1;
wire    ap_block_state8_pp0_stage1_iter2;
wire    ap_block_pp0_stage1_11001;
wire   [1:0] select_ln19_7_fu_553_p3;
reg   [1:0] select_ln19_7_reg_1082;
wire   [5:0] select_ln20_fu_617_p3;
reg   [5:0] select_ln20_reg_1089;
wire   [1:0] select_ln20_6_fu_625_p3;
reg   [1:0] select_ln20_6_reg_1095;
wire   [0:0] select_ln20_7_fu_634_p3;
reg   [0:0] select_ln20_7_reg_1101;
reg   [0:0] select_ln20_7_reg_1101_pp0_iter1_reg;
wire   [4:0] empty_73_fu_730_p1;
reg   [4:0] empty_73_reg_1109;
reg   [4:0] empty_73_reg_1109_pp0_iter1_reg;
wire   [5:0] select_ln20_10_fu_757_p3;
reg   [5:0] select_ln20_10_reg_1121;
wire   [5:0] add_ln25_fu_763_p2;
reg   [5:0] add_ln25_reg_1126;
reg    ap_enable_reg_pp0_iter1;
wire   [5:0] add_ln33_fu_795_p2;
reg   [5:0] add_ln33_reg_1131;
wire   [8:0] add_ln33_2_fu_816_p2;
reg   [8:0] add_ln33_2_reg_1138;
wire   [15:0] select_ln33_8_fu_895_p3;
reg   [15:0] select_ln33_8_reg_1143;
wire   [15:0] select_ln33_9_fu_916_p3;
reg   [15:0] select_ln33_9_reg_1148;
wire    ap_block_pp0_stage1_subdone;
reg    ap_condition_pp0_exit_iter0_state4;
reg    ap_enable_reg_pp0_iter2;
reg   [6:0] ap_phi_mux_indvar_flatten47_phi_fu_226_p4;
wire    ap_block_pp0_stage0;
reg   [1:0] ap_phi_mux_ii_phi_fu_238_p4;
reg   [5:0] ap_phi_mux_indvar_flatten_phi_fu_250_p4;
reg   [1:0] ap_phi_mux_jj_phi_fu_261_p4;
reg   [5:0] ap_phi_mux_kk_0_i_i_phi_fu_273_p4;
wire    ap_block_pp0_stage1;
wire   [63:0] sext_ln32_fu_752_p1;
wire   [63:0] zext_ln33_9_fu_822_p1;
wire   [63:0] sext_ln33_fu_854_p1;
wire   [63:0] sext_ln33_3_fu_935_p1;
wire   [63:0] sext_ln33_4_fu_952_p1;
reg    ap_block_state1;
wire   [15:0] select_ln33_fu_834_p3;
wire   [15:0] select_ln33_7_fu_873_p3;
wire   [16:0] zext_ln19_fu_293_p1;
wire   [16:0] empty_68_fu_296_p2;
wire   [16:0] j_cast_i_i_fu_290_p1;
wire   [16:0] add_ln22_fu_306_p2;
wire   [0:0] tmp_9_fu_321_p3;
wire   [0:0] icmp_ln24_fu_329_p2;
wire   [17:0] ii_cast_i_i_fu_346_p1;
wire   [4:0] ii_cast_fu_350_p1;
wire   [17:0] empty_69_fu_354_p2;
wire   [17:0] zext_ln20_fu_370_p1;
wire   [17:0] add_ln22_2_fu_374_p2;
wire   [0:0] tmp_10_fu_379_p3;
wire   [0:0] icmp_ln24_2_fu_387_p2;
wire   [0:0] or_ln23_fu_393_p2;
wire   [0:0] empty_70_fu_364_p2;
wire   [17:0] ii_cast_i_i_mid1_fu_431_p1;
wire   [4:0] ii_cast_mid1_fu_435_p1;
wire   [17:0] p_mid111_fu_439_p2;
wire   [0:0] p_mid113_fu_449_p2;
wire   [17:0] zext_ln20_2_fu_474_p1;
wire   [17:0] add_ln22_3_fu_478_p2;
wire   [0:0] tmp_11_fu_483_p3;
wire   [0:0] icmp_ln24_3_fu_491_p2;
wire   [0:0] or_ln23_9_fu_497_p2;
wire   [0:0] select_ln19_9_fu_455_p3;
wire   [2:0] zext_ln22_fu_521_p1;
wire   [2:0] tmp1_fu_531_p2;
wire   [9:0] tmp1_cast_fu_537_p1;
wire   [9:0] empty_71_fu_541_p2;
wire   [4:0] row_coord_int_mid131_fu_569_p3;
wire   [4:0] row_coord_int_fu_525_p3;
wire   [9:0] col_coord_int_mid139_fu_575_p3;
wire   [9:0] col_coord_int_fu_546_p3;
wire   [0:0] icmp_ln25_fu_600_p2;
wire   [0:0] xor_ln19_fu_595_p2;
wire   [0:0] and_ln19_fu_606_p2;
wire   [0:0] or_ln20_fu_612_p2;
wire   [0:0] select_ln19_10_fu_564_p3;
wire   [4:0] select_ln19_8_fu_559_p3;
wire   [2:0] zext_ln22_2_fu_631_p1;
wire   [2:0] tmp1_mid1_fu_648_p2;
wire   [9:0] tmp1_cast_mid1_fu_654_p1;
wire   [9:0] p_mid1_fu_658_p2;
wire   [4:0] row_coord_int_mid1_fu_641_p3;
wire   [4:0] select_ln19_11_fu_581_p3;
wire   [4:0] select_ln20_8_fu_670_p3;
wire   [9:0] tmp_s_fu_678_p3;
wire   [6:0] tmp_3_fu_690_p3;
wire   [10:0] zext_ln32_fu_686_p1;
wire   [10:0] zext_ln32_9_fu_698_p1;
wire   [10:0] sub_ln32_fu_702_p2;
wire   [9:0] col_coord_int_mid1_fu_663_p3;
wire   [9:0] select_ln19_12_fu_588_p3;
wire   [9:0] select_ln20_9_fu_712_p3;
wire   [11:0] sext_ln20_fu_708_p1;
wire   [11:0] zext_ln32_10_fu_720_p1;
wire   [11:0] add_ln32_fu_724_p2;
wire   [2:0] lshr_ln_fu_734_p4;
wire   [14:0] tmp_12_fu_744_p3;
wire   [3:0] tmp_fu_771_p3;
wire   [4:0] zext_ln33_6_fu_778_p1;
wire   [4:0] zext_ln33_fu_768_p1;
wire   [4:0] sub_ln33_fu_782_p2;
wire   [5:0] sub_ln33_cast_fu_788_p1;
wire   [5:0] zext_ln33_7_fu_792_p1;
wire   [3:0] trunc_ln33_fu_801_p1;
wire   [8:0] tmp_30_cast_fu_805_p3;
wire   [8:0] zext_ln33_8_fu_813_p1;
wire   [15:0] trunc_ln32_fu_826_p1;
wire   [15:0] bitcast_ln32_fu_830_p1;
wire   [4:0] or_ln25_fu_842_p2;
wire   [10:0] tmp_13_fu_847_p3;
wire   [15:0] tmp_17_i_i_fu_859_p4;
wire   [15:0] bitcast_ln32_7_fu_869_p1;
wire   [15:0] tmp_18_i_i_fu_881_p4;
wire   [15:0] bitcast_ln32_8_fu_891_p1;
wire   [15:0] tmp_19_i_i_fu_902_p4;
wire   [15:0] bitcast_ln32_9_fu_912_p1;
wire   [4:0] or_ln25_5_fu_923_p2;
wire   [10:0] tmp_14_fu_928_p3;
wire   [4:0] or_ln25_6_fu_940_p2;
wire   [10:0] tmp_15_fu_945_p3;
wire    ap_CS_fsm_state9;
reg   [4:0] ap_NS_fsm;
wire    ap_block_pp0_stage0_subdone;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 5'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b1 == ap_condition_pp0_exit_iter0_state4) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_subdone))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_subdone))) begin
            if ((1'b1 == ap_condition_pp0_exit_iter0_state4)) begin
                ap_enable_reg_pp0_iter1 <= (1'b1 ^ ap_condition_pp0_exit_iter0_state4);
            end else if ((1'b1 == 1'b1)) begin
                ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
            end
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_subdone))) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            ap_enable_reg_pp0_iter2 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln19_reg_1020 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        ii_reg_234 <= select_ln19_7_reg_1082;
    end else if ((1'b1 == ap_CS_fsm_state2)) begin
        ii_reg_234 <= 2'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln19_reg_1020 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        indvar_flatten47_reg_222 <= add_ln19_2_reg_1077;
    end else if ((1'b1 == ap_CS_fsm_state2)) begin
        indvar_flatten47_reg_222 <= 7'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln19_reg_1020 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        indvar_flatten_reg_246 <= select_ln20_10_reg_1121;
    end else if ((1'b1 == ap_CS_fsm_state2)) begin
        indvar_flatten_reg_246 <= 6'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln19_reg_1020 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        jj_reg_257 <= select_ln20_6_reg_1095;
    end else if ((1'b1 == ap_CS_fsm_state2)) begin
        jj_reg_257 <= 2'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln19_reg_1020_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001))) begin
        kk_0_i_i_reg_269 <= add_ln25_reg_1126;
    end else if ((1'b1 == ap_CS_fsm_state2)) begin
        kk_0_i_i_reg_269 <= 6'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
        add_ln19_2_reg_1077 <= add_ln19_2_fu_515_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (icmp_ln19_fu_405_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        add_ln19_reg_1024 <= add_ln19_fu_411_p2;
        add_ln20_2_reg_1072 <= add_ln20_2_fu_509_p2;
        add_ln20_reg_1059 <= add_ln20_fu_468_p2;
        icmp_ln20_reg_1029 <= icmp_ln20_fu_417_p2;
        or_ln23_10_reg_1065 <= or_ln23_10_fu_503_p2;
        or_ln23_8_reg_1052 <= or_ln23_8_fu_463_p2;
        p_cast5_i_i_mid1_reg_1046 <= p_cast5_i_i_mid1_fu_444_p2;
        select_ln19_reg_1041 <= select_ln19_fu_423_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln19_reg_1020 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        add_ln25_reg_1126 <= add_ln25_fu_763_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln19_reg_1020_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001))) begin
        add_ln33_2_reg_1138 <= add_ln33_2_fu_816_p2;
        add_ln33_reg_1131 <= add_ln33_fu_795_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln19_reg_1020 == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001))) begin
        empty_73_reg_1109 <= empty_73_fu_730_p1;
        select_ln20_7_reg_1101 <= select_ln20_7_fu_634_p3;
        select_ln20_reg_1089 <= select_ln20_fu_617_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_11001))) begin
        empty_73_reg_1109_pp0_iter1_reg <= empty_73_reg_1109;
        select_ln20_7_reg_1101_pp0_iter1_reg <= select_ln20_7_reg_1101;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state1)) begin
        empty_reg_972 <= empty_fu_285_p1;
        indices_01_read_reg_957 <= indices_01_dout;
        indices_12_read_reg_967 <= indices_12_dout;
        trunc_ln250_reg_962 <= trunc_ln250_fu_280_p1;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        icmp_ln19_reg_1020 <= icmp_ln19_fu_405_p2;
        icmp_ln19_reg_1020_pp0_iter1_reg <= icmp_ln19_reg_1020;
        icmp_ln19_reg_1020_pp0_iter2_reg <= icmp_ln19_reg_1020_pp0_iter1_reg;
        is_padding_reg_1013 <= is_padding_fu_399_p2;
        p_cast5_i_i_reg_1007 <= p_cast5_i_i_fu_359_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        or_ln23_6_reg_997 <= or_ln23_6_fu_335_p2;
        p_cast_i_i_reg_979 <= p_cast_i_i_fu_302_p1;
        p_cast_reg_991 <= p_cast_fu_316_p2;
        p_mid137_reg_1002 <= p_mid137_fu_341_p2;
        sext_ln22_reg_985 <= sext_ln22_fu_312_p1;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln19_reg_1020 == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001))) begin
        select_ln19_7_reg_1082 <= select_ln19_7_fu_553_p3;
        select_ln20_10_reg_1121 <= select_ln20_10_fu_757_p3;
        select_ln20_6_reg_1095 <= select_ln20_6_fu_625_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (icmp_ln19_reg_1020_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        select_ln33_8_reg_1143 <= select_ln33_8_fu_895_p3;
        select_ln33_9_reg_1148 <= select_ln33_9_fu_916_p3;
    end
end

always @ (*) begin
    if ((icmp_ln19_reg_1020 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state4 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state4 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state9)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln19_reg_1020 == 1'd0) & (1'b0 == ap_block_pp0_stage0))) begin
        ap_phi_mux_ii_phi_fu_238_p4 = select_ln19_7_reg_1082;
    end else begin
        ap_phi_mux_ii_phi_fu_238_p4 = ii_reg_234;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln19_reg_1020 == 1'd0) & (1'b0 == ap_block_pp0_stage0))) begin
        ap_phi_mux_indvar_flatten47_phi_fu_226_p4 = add_ln19_2_reg_1077;
    end else begin
        ap_phi_mux_indvar_flatten47_phi_fu_226_p4 = indvar_flatten47_reg_222;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln19_reg_1020 == 1'd0) & (1'b0 == ap_block_pp0_stage0))) begin
        ap_phi_mux_indvar_flatten_phi_fu_250_p4 = select_ln20_10_reg_1121;
    end else begin
        ap_phi_mux_indvar_flatten_phi_fu_250_p4 = indvar_flatten_reg_246;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln19_reg_1020 == 1'd0) & (1'b0 == ap_block_pp0_stage0))) begin
        ap_phi_mux_jj_phi_fu_261_p4 = select_ln20_6_reg_1095;
    end else begin
        ap_phi_mux_jj_phi_fu_261_p4 = jj_reg_257;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln19_reg_1020_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage1))) begin
        ap_phi_mux_kk_0_i_i_phi_fu_273_p4 = add_ln25_reg_1126;
    end else begin
        ap_phi_mux_kk_0_i_i_phi_fu_273_p4 = kk_0_i_i_reg_269;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state9)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((ap_enable_reg_pp0_iter2 == 1'b1)) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ifmap_vec_address0 = sext_ln33_4_fu_952_p1;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0))) begin
            ifmap_vec_address0 = sext_ln33_fu_854_p1;
        end else begin
            ifmap_vec_address0 = 'bx;
        end
    end else begin
        ifmap_vec_address0 = 'bx;
    end
end

always @ (*) begin
    if ((ap_enable_reg_pp0_iter2 == 1'b1)) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ifmap_vec_address1 = sext_ln33_3_fu_935_p1;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0))) begin
            ifmap_vec_address1 = zext_ln33_9_fu_822_p1;
        end else begin
            ifmap_vec_address1 = 'bx;
        end
    end else begin
        ifmap_vec_address1 = 'bx;
    end
end

always @ (*) begin
    if ((((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_11001)) | ((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
        ifmap_vec_ce0 = 1'b1;
    end else begin
        ifmap_vec_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1_11001)) | ((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
        ifmap_vec_ce1 = 1'b1;
    end else begin
        ifmap_vec_ce1 = 1'b0;
    end
end

always @ (*) begin
    if ((ap_enable_reg_pp0_iter2 == 1'b1)) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ifmap_vec_d0 = select_ln33_9_reg_1148;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0))) begin
            ifmap_vec_d0 = select_ln33_7_fu_873_p3;
        end else begin
            ifmap_vec_d0 = 'bx;
        end
    end else begin
        ifmap_vec_d0 = 'bx;
    end
end

always @ (*) begin
    if ((ap_enable_reg_pp0_iter2 == 1'b1)) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage1) & (1'b0 == ap_block_pp0_stage1))) begin
            ifmap_vec_d1 = select_ln33_8_reg_1143;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0))) begin
            ifmap_vec_d1 = select_ln33_fu_834_p3;
        end else begin
            ifmap_vec_d1 = 'bx;
        end
    end else begin
        ifmap_vec_d1 = 'bx;
    end
end

always @ (*) begin
    if ((((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln19_reg_1020_pp0_iter2_reg == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001)) | ((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (icmp_ln19_reg_1020_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
        ifmap_vec_we0 = 1'b1;
    end else begin
        ifmap_vec_we0 = 1'b0;
    end
end

always @ (*) begin
    if ((((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln19_reg_1020_pp0_iter2_reg == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001)) | ((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (icmp_ln19_reg_1020_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
        ifmap_vec_we1 = 1'b1;
    end else begin
        ifmap_vec_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001)) | ((1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b0 == ap_block_pp0_stage1_11001)) | ((1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage1_11001)) | ((1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001)))) begin
        in_data_ce0 = 1'b1;
    end else begin
        in_data_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_01_blk_n = indices_01_empty_n;
    end else begin
        indices_01_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_01_out_blk_n = indices_01_out_full_n;
    end else begin
        indices_01_out_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((indices_12_out_full_n == 1'b0) | (indices_01_out_full_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_01_out_write = 1'b1;
    end else begin
        indices_01_out_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((indices_12_out_full_n == 1'b0) | (indices_01_out_full_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_01_read = 1'b1;
    end else begin
        indices_01_read = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_12_blk_n = indices_12_empty_n;
    end else begin
        indices_12_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_12_out_blk_n = indices_12_out_full_n;
    end else begin
        indices_12_out_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((indices_12_out_full_n == 1'b0) | (indices_01_out_full_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_12_out_write = 1'b1;
    end else begin
        indices_12_out_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((indices_12_out_full_n == 1'b0) | (indices_01_out_full_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_12_read = 1'b1;
    end else begin
        indices_12_read = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((indices_12_out_full_n == 1'b0) | (indices_01_out_full_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_state2 : begin
            ap_NS_fsm = ap_ST_fsm_pp0_stage0;
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_pp0_stage1 : begin
            if ((~((ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln19_reg_1020 == 1'd1) & (1'b0 == ap_block_pp0_stage1_subdone)) & ~((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b0) & (1'b0 == ap_block_pp0_stage1_subdone)) & (1'b0 == ap_block_pp0_stage1_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if ((((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b0) & (1'b0 == ap_block_pp0_stage1_subdone)) | ((ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln19_reg_1020 == 1'd1) & (1'b0 == ap_block_pp0_stage1_subdone)))) begin
                ap_NS_fsm = ap_ST_fsm_state9;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end
        end
        ap_ST_fsm_state9 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln19_2_fu_515_p2 = (indvar_flatten47_reg_222 + 7'd1);

assign add_ln19_fu_411_p2 = (ap_phi_mux_ii_phi_fu_238_p4 + 2'd1);

assign add_ln20_2_fu_509_p2 = (ap_phi_mux_indvar_flatten_phi_fu_250_p4 + 6'd1);

assign add_ln20_fu_468_p2 = (select_ln19_fu_423_p3 + 2'd1);

assign add_ln22_2_fu_374_p2 = ((sext_ln22_reg_985) + (zext_ln20_fu_370_p1));

assign add_ln22_3_fu_478_p2 = ((sext_ln22_reg_985) + (zext_ln20_2_fu_474_p1));

assign add_ln22_fu_306_p2 = ((j_cast_i_i_fu_290_p1) + (17'd131071));

assign add_ln25_fu_763_p2 = (select_ln20_reg_1089 + 6'd4);

assign add_ln32_fu_724_p2 = ((sext_ln20_fu_708_p1) + (zext_ln32_10_fu_720_p1));

assign add_ln33_2_fu_816_p2 = (tmp_30_cast_fu_805_p3 + zext_ln33_8_fu_813_p1);

assign add_ln33_fu_795_p2 = ((sub_ln33_cast_fu_788_p1) + (zext_ln33_7_fu_792_p1));

assign and_ln19_fu_606_p2 = (xor_ln19_fu_595_p2 & icmp_ln25_fu_600_p2);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_pp0_stage1 = ap_CS_fsm[32'd3];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state9 = ap_CS_fsm[32'd4];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((indices_12_out_full_n == 1'b0) | (indices_01_out_full_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0));
end

assign ap_block_state3_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage1_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage1_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage1_iter2 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign bitcast_ln32_7_fu_869_p1 = tmp_17_i_i_fu_859_p4;

assign bitcast_ln32_8_fu_891_p1 = tmp_18_i_i_fu_881_p4;

assign bitcast_ln32_9_fu_912_p1 = tmp_19_i_i_fu_902_p4;

assign bitcast_ln32_fu_830_p1 = trunc_ln32_fu_826_p1;

assign col_coord_int_fu_546_p3 = ((is_padding_reg_1013[0:0] == 1'b1) ? 10'd0 : empty_71_fu_541_p2);

assign col_coord_int_mid139_fu_575_p3 = ((or_ln23_8_reg_1052[0:0] == 1'b1) ? 10'd0 : p_mid137_reg_1002);

assign col_coord_int_mid1_fu_663_p3 = ((or_ln23_10_reg_1065[0:0] == 1'b1) ? 10'd0 : p_mid1_fu_658_p2);

assign empty_68_fu_296_p2 = ((zext_ln19_fu_293_p1) + (17'd131071));

assign empty_69_fu_354_p2 = ((p_cast_i_i_reg_979) + (ii_cast_i_i_fu_346_p1));

assign empty_70_fu_364_p2 = ((empty_69_fu_354_p2 > 18'd27) ? 1'b1 : 1'b0);

assign empty_71_fu_541_p2 = ((tmp1_cast_fu_537_p1) + (empty_reg_972));

assign empty_73_fu_730_p1 = select_ln20_fu_617_p3[4:0];

assign empty_fu_285_p1 = indices_12_dout[9:0];

assign icmp_ln19_fu_405_p2 = ((ap_phi_mux_indvar_flatten47_phi_fu_226_p4 == 7'd72) ? 1'b1 : 1'b0);

assign icmp_ln20_fu_417_p2 = ((ap_phi_mux_indvar_flatten_phi_fu_250_p4 == 6'd24) ? 1'b1 : 1'b0);

assign icmp_ln24_2_fu_387_p2 = (((add_ln22_2_fu_374_p2) > (18'd27)) ? 1'b1 : 1'b0);

assign icmp_ln24_3_fu_491_p2 = (((add_ln22_3_fu_478_p2) > (18'd27)) ? 1'b1 : 1'b0);

assign icmp_ln24_fu_329_p2 = (((add_ln22_fu_306_p2) > (17'd27)) ? 1'b1 : 1'b0);

assign icmp_ln25_fu_600_p2 = ((ap_phi_mux_kk_0_i_i_phi_fu_273_p4 == 6'd32) ? 1'b1 : 1'b0);

assign ii_cast_fu_350_p1 = ap_phi_mux_ii_phi_fu_238_p4;

assign ii_cast_i_i_fu_346_p1 = ap_phi_mux_ii_phi_fu_238_p4;

assign ii_cast_i_i_mid1_fu_431_p1 = add_ln19_fu_411_p2;

assign ii_cast_mid1_fu_435_p1 = add_ln19_fu_411_p2;

assign in_data_address0 = sext_ln32_fu_752_p1;

assign indices_01_out_din = indices_01_dout[4:0];

assign indices_12_out_din = indices_12_dout[9:0];

assign is_padding_fu_399_p2 = (or_ln23_fu_393_p2 | empty_70_fu_364_p2);

assign j_cast_i_i_fu_290_p1 = indices_12_read_reg_967;

assign lshr_ln_fu_734_p4 = {{select_ln20_fu_617_p3[4:2]}};

assign or_ln20_fu_612_p2 = (icmp_ln20_reg_1029 | and_ln19_fu_606_p2);

assign or_ln23_10_fu_503_p2 = (select_ln19_9_fu_455_p3 | or_ln23_9_fu_497_p2);

assign or_ln23_6_fu_335_p2 = (tmp_9_fu_321_p3 | icmp_ln24_fu_329_p2);

assign or_ln23_8_fu_463_p2 = (p_mid113_fu_449_p2 | or_ln23_6_reg_997);

assign or_ln23_9_fu_497_p2 = (tmp_11_fu_483_p3 | icmp_ln24_3_fu_491_p2);

assign or_ln23_fu_393_p2 = (tmp_10_fu_379_p3 | icmp_ln24_2_fu_387_p2);

assign or_ln25_5_fu_923_p2 = (empty_73_reg_1109_pp0_iter1_reg | 5'd2);

assign or_ln25_6_fu_940_p2 = (empty_73_reg_1109_pp0_iter1_reg | 5'd3);

assign or_ln25_fu_842_p2 = (empty_73_reg_1109_pp0_iter1_reg | 5'd1);

assign p_cast5_i_i_fu_359_p2 = (p_cast_reg_991 + ii_cast_fu_350_p1);

assign p_cast5_i_i_mid1_fu_444_p2 = (p_cast_reg_991 + ii_cast_mid1_fu_435_p1);

assign p_cast_fu_316_p2 = ((trunc_ln250_reg_962) + (5'd31));

assign p_cast_i_i_fu_302_p1 = (empty_68_fu_296_p2);

assign p_mid111_fu_439_p2 = ((p_cast_i_i_reg_979) + (ii_cast_i_i_mid1_fu_431_p1));

assign p_mid113_fu_449_p2 = ((p_mid111_fu_439_p2 > 18'd27) ? 1'b1 : 1'b0);

assign p_mid137_fu_341_p2 = ((empty_reg_972) + (10'd1023));

assign p_mid1_fu_658_p2 = ((tmp1_cast_mid1_fu_654_p1) + (empty_reg_972));

assign row_coord_int_fu_525_p3 = ((is_padding_reg_1013[0:0] == 1'b1) ? 5'd0 : p_cast5_i_i_reg_1007);

assign row_coord_int_mid131_fu_569_p3 = ((or_ln23_8_reg_1052[0:0] == 1'b1) ? 5'd0 : p_cast5_i_i_mid1_reg_1046);

assign row_coord_int_mid1_fu_641_p3 = ((or_ln23_10_reg_1065[0:0] == 1'b1) ? 5'd0 : select_ln19_8_fu_559_p3);

assign select_ln19_10_fu_564_p3 = ((icmp_ln20_reg_1029[0:0] == 1'b1) ? or_ln23_8_reg_1052 : is_padding_reg_1013);

assign select_ln19_11_fu_581_p3 = ((icmp_ln20_reg_1029[0:0] == 1'b1) ? row_coord_int_mid131_fu_569_p3 : row_coord_int_fu_525_p3);

assign select_ln19_12_fu_588_p3 = ((icmp_ln20_reg_1029[0:0] == 1'b1) ? col_coord_int_mid139_fu_575_p3 : col_coord_int_fu_546_p3);

assign select_ln19_7_fu_553_p3 = ((icmp_ln20_reg_1029[0:0] == 1'b1) ? add_ln19_reg_1024 : ii_reg_234);

assign select_ln19_8_fu_559_p3 = ((icmp_ln20_reg_1029[0:0] == 1'b1) ? p_cast5_i_i_mid1_reg_1046 : p_cast5_i_i_reg_1007);

assign select_ln19_9_fu_455_p3 = ((icmp_ln20_fu_417_p2[0:0] == 1'b1) ? p_mid113_fu_449_p2 : empty_70_fu_364_p2);

assign select_ln19_fu_423_p3 = ((icmp_ln20_fu_417_p2[0:0] == 1'b1) ? 2'd0 : ap_phi_mux_jj_phi_fu_261_p4);

assign select_ln20_10_fu_757_p3 = ((icmp_ln20_reg_1029[0:0] == 1'b1) ? 6'd1 : add_ln20_2_reg_1072);

assign select_ln20_6_fu_625_p3 = ((and_ln19_fu_606_p2[0:0] == 1'b1) ? add_ln20_reg_1059 : select_ln19_reg_1041);

assign select_ln20_7_fu_634_p3 = ((and_ln19_fu_606_p2[0:0] == 1'b1) ? or_ln23_10_reg_1065 : select_ln19_10_fu_564_p3);

assign select_ln20_8_fu_670_p3 = ((and_ln19_fu_606_p2[0:0] == 1'b1) ? row_coord_int_mid1_fu_641_p3 : select_ln19_11_fu_581_p3);

assign select_ln20_9_fu_712_p3 = ((and_ln19_fu_606_p2[0:0] == 1'b1) ? col_coord_int_mid1_fu_663_p3 : select_ln19_12_fu_588_p3);

assign select_ln20_fu_617_p3 = ((or_ln20_fu_612_p2[0:0] == 1'b1) ? 6'd0 : ap_phi_mux_kk_0_i_i_phi_fu_273_p4);

assign select_ln33_7_fu_873_p3 = ((select_ln20_7_reg_1101_pp0_iter1_reg[0:0] == 1'b1) ? 16'd0 : bitcast_ln32_7_fu_869_p1);

assign select_ln33_8_fu_895_p3 = ((select_ln20_7_reg_1101_pp0_iter1_reg[0:0] == 1'b1) ? 16'd0 : bitcast_ln32_8_fu_891_p1);

assign select_ln33_9_fu_916_p3 = ((select_ln20_7_reg_1101_pp0_iter1_reg[0:0] == 1'b1) ? 16'd0 : bitcast_ln32_9_fu_912_p1);

assign select_ln33_fu_834_p3 = ((select_ln20_7_reg_1101_pp0_iter1_reg[0:0] == 1'b1) ? 16'd0 : bitcast_ln32_fu_830_p1);

assign sext_ln20_fu_708_p1 = (sub_ln32_fu_702_p2);

assign sext_ln22_fu_312_p1 = add_ln22_fu_306_p2;

assign sext_ln32_fu_752_p1 = (tmp_12_fu_744_p3);

assign sext_ln33_3_fu_935_p1 = (tmp_14_fu_928_p3);

assign sext_ln33_4_fu_952_p1 = (tmp_15_fu_945_p3);

assign sext_ln33_fu_854_p1 = (tmp_13_fu_847_p3);

assign sub_ln32_fu_702_p2 = (zext_ln32_fu_686_p1 - zext_ln32_9_fu_698_p1);

assign sub_ln33_cast_fu_788_p1 = (sub_ln33_fu_782_p2);

assign sub_ln33_fu_782_p2 = (zext_ln33_6_fu_778_p1 - zext_ln33_fu_768_p1);

assign tmp1_cast_fu_537_p1 = (tmp1_fu_531_p2);

assign tmp1_cast_mid1_fu_654_p1 = (tmp1_mid1_fu_648_p2);

assign tmp1_fu_531_p2 = ((zext_ln22_fu_521_p1) + (3'd7));

assign tmp1_mid1_fu_648_p2 = ((zext_ln22_2_fu_631_p1) + (3'd7));

assign tmp_10_fu_379_p3 = add_ln22_2_fu_374_p2[32'd17];

assign tmp_11_fu_483_p3 = add_ln22_3_fu_478_p2[32'd17];

assign tmp_12_fu_744_p3 = {{add_ln32_fu_724_p2}, {lshr_ln_fu_734_p4}};

assign tmp_13_fu_847_p3 = {{add_ln33_reg_1131}, {or_ln25_fu_842_p2}};

assign tmp_14_fu_928_p3 = {{add_ln33_reg_1131}, {or_ln25_5_fu_923_p2}};

assign tmp_15_fu_945_p3 = {{add_ln33_reg_1131}, {or_ln25_6_fu_940_p2}};

assign tmp_17_i_i_fu_859_p4 = {{in_data_q0[31:16]}};

assign tmp_18_i_i_fu_881_p4 = {{in_data_q0[47:32]}};

assign tmp_19_i_i_fu_902_p4 = {{in_data_q0[63:48]}};

assign tmp_30_cast_fu_805_p3 = {{trunc_ln33_fu_801_p1}, {5'd0}};

assign tmp_3_fu_690_p3 = {{select_ln20_8_fu_670_p3}, {2'd0}};

assign tmp_9_fu_321_p3 = add_ln22_fu_306_p2[32'd16];

assign tmp_fu_771_p3 = {{select_ln19_7_reg_1082}, {2'd0}};

assign tmp_s_fu_678_p3 = {{select_ln20_8_fu_670_p3}, {5'd0}};

assign trunc_ln250_fu_280_p1 = indices_01_dout[4:0];

assign trunc_ln32_fu_826_p1 = in_data_q0[15:0];

assign trunc_ln33_fu_801_p1 = add_ln33_fu_795_p2[3:0];

assign xor_ln19_fu_595_p2 = (icmp_ln20_reg_1029 ^ 1'd1);

assign zext_ln19_fu_293_p1 = indices_01_read_reg_957;

assign zext_ln20_2_fu_474_p1 = add_ln20_fu_468_p2;

assign zext_ln20_fu_370_p1 = ap_phi_mux_jj_phi_fu_261_p4;

assign zext_ln22_2_fu_631_p1 = add_ln20_reg_1059;

assign zext_ln22_fu_521_p1 = jj_reg_257;

assign zext_ln32_10_fu_720_p1 = select_ln20_9_fu_712_p3;

assign zext_ln32_9_fu_698_p1 = tmp_3_fu_690_p3;

assign zext_ln32_fu_686_p1 = tmp_s_fu_678_p3;

assign zext_ln33_6_fu_778_p1 = tmp_fu_771_p3;

assign zext_ln33_7_fu_792_p1 = select_ln20_6_reg_1095;

assign zext_ln33_8_fu_813_p1 = select_ln20_reg_1089;

assign zext_ln33_9_fu_822_p1 = add_ln33_2_reg_1138;

assign zext_ln33_fu_768_p1 = select_ln19_7_reg_1082;

endmodule //td_fused_top_tdf7_readInputs53
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf8_17 (
        in_data_address0,
        in_data_ce0,
        in_data_d0,
        in_data_q0,
        in_data_we0,
        in_data_address1,
        in_data_ce1,
        in_data_d1,
        in_data_q1,
        in_data_we1,
        out_data_address0,
        out_data_ce0,
        out_data_d0,
        out_data_q0,
        out_data_we0,
        out_data_address1,
        out_data_ce1,
        out_data_d1,
        out_data_q1,
        out_data_we1,
        filter_data_address0,
        filter_data_ce0,
        filter_data_d0,
        filter_data_q0,
        filter_data_we0,
        filter_data_address1,
        filter_data_ce1,
        filter_data_d1,
        filter_data_q1,
        filter_data_we1,
        adjustments_address0,
        adjustments_ce0,
        adjustments_d0,
        adjustments_q0,
        adjustments_we0,
        adjustments_address1,
        adjustments_ce1,
        adjustments_d1,
        adjustments_q1,
        adjustments_we1,
        ap_clk,
        ap_rst,
        in_data_empty_n,
        in_data_read,
        out_data_full_n,
        out_data_write,
        ap_start,
        ap_done,
        ap_ready,
        ap_idle,
        ap_continue
);


output  [12:0] in_data_address0;
output   in_data_ce0;
output  [63:0] in_data_d0;
input  [63:0] in_data_q0;
output   in_data_we0;
output  [12:0] in_data_address1;
output   in_data_ce1;
output  [63:0] in_data_d1;
input  [63:0] in_data_q1;
output   in_data_we1;
output  [13:0] out_data_address0;
output   out_data_ce0;
output  [63:0] out_data_d0;
input  [63:0] out_data_q0;
output   out_data_we0;
output  [13:0] out_data_address1;
output   out_data_ce1;
output  [63:0] out_data_d1;
input  [63:0] out_data_q1;
output   out_data_we1;
output  [16:0] filter_data_address0;
output   filter_data_ce0;
output  [15:0] filter_data_d0;
input  [15:0] filter_data_q0;
output   filter_data_we0;
output  [16:0] filter_data_address1;
output   filter_data_ce1;
output  [15:0] filter_data_d1;
input  [15:0] filter_data_q1;
output   filter_data_we1;
output  [7:0] adjustments_address0;
output   adjustments_ce0;
output  [47:0] adjustments_d0;
input  [47:0] adjustments_q0;
output   adjustments_we0;
output  [7:0] adjustments_address1;
output   adjustments_ce1;
output  [47:0] adjustments_d1;
input  [47:0] adjustments_q1;
output   adjustments_we1;
input   ap_clk;
input   ap_rst;
input   in_data_empty_n;
output   in_data_read;
input   out_data_full_n;
output   out_data_write;
input   ap_start;
output   ap_done;
output   ap_ready;
output   ap_idle;
input   ap_continue;

reg ap_done;
reg ap_ready;
reg ap_idle;

wire   [12:0] dataflow_in_loop_TOP_LOOP37454_U0_in_data_address0;
wire    dataflow_in_loop_TOP_LOOP37454_U0_in_data_ce0;
wire   [63:0] dataflow_in_loop_TOP_LOOP37454_U0_in_data_d0;
wire    dataflow_in_loop_TOP_LOOP37454_U0_in_data_we0;
wire   [12:0] dataflow_in_loop_TOP_LOOP37454_U0_in_data_address1;
wire    dataflow_in_loop_TOP_LOOP37454_U0_in_data_ce1;
wire   [63:0] dataflow_in_loop_TOP_LOOP37454_U0_in_data_d1;
wire    dataflow_in_loop_TOP_LOOP37454_U0_in_data_we1;
wire   [16:0] dataflow_in_loop_TOP_LOOP37454_U0_filter_data_address0;
wire    dataflow_in_loop_TOP_LOOP37454_U0_filter_data_ce0;
wire   [15:0] dataflow_in_loop_TOP_LOOP37454_U0_filter_data_d0;
wire    dataflow_in_loop_TOP_LOOP37454_U0_filter_data_we0;
wire   [16:0] dataflow_in_loop_TOP_LOOP37454_U0_filter_data_address1;
wire    dataflow_in_loop_TOP_LOOP37454_U0_filter_data_ce1;
wire   [15:0] dataflow_in_loop_TOP_LOOP37454_U0_filter_data_d1;
wire    dataflow_in_loop_TOP_LOOP37454_U0_filter_data_we1;
wire   [7:0] dataflow_in_loop_TOP_LOOP37454_U0_adjustments_address0;
wire    dataflow_in_loop_TOP_LOOP37454_U0_adjustments_ce0;
wire   [47:0] dataflow_in_loop_TOP_LOOP37454_U0_adjustments_d0;
wire    dataflow_in_loop_TOP_LOOP37454_U0_adjustments_we0;
wire   [7:0] dataflow_in_loop_TOP_LOOP37454_U0_adjustments_address1;
wire    dataflow_in_loop_TOP_LOOP37454_U0_adjustments_ce1;
wire   [47:0] dataflow_in_loop_TOP_LOOP37454_U0_adjustments_d1;
wire    dataflow_in_loop_TOP_LOOP37454_U0_adjustments_we1;
wire   [13:0] dataflow_in_loop_TOP_LOOP37454_U0_out_data_address0;
wire    dataflow_in_loop_TOP_LOOP37454_U0_out_data_ce0;
wire   [63:0] dataflow_in_loop_TOP_LOOP37454_U0_out_data_d0;
wire    dataflow_in_loop_TOP_LOOP37454_U0_out_data_we0;
wire   [13:0] dataflow_in_loop_TOP_LOOP37454_U0_out_data_address1;
wire    dataflow_in_loop_TOP_LOOP37454_U0_out_data_ce1;
wire   [63:0] dataflow_in_loop_TOP_LOOP37454_U0_out_data_d1;
wire    dataflow_in_loop_TOP_LOOP37454_U0_out_data_we1;
wire    dataflow_in_loop_TOP_LOOP37454_U0_ap_start;
wire    dataflow_in_loop_TOP_LOOP37454_U0_in_data_read;
wire    dataflow_in_loop_TOP_LOOP37454_U0_out_data_write;
wire    dataflow_in_loop_TOP_LOOP37454_U0_ap_done;
wire    dataflow_in_loop_TOP_LOOP37454_U0_ap_ready;
wire    dataflow_in_loop_TOP_LOOP37454_U0_ap_idle;
reg    dataflow_in_loop_TOP_LOOP37454_U0_ap_continue;
wire    dataflow_in_loop_TOP_LOOP37454_U0_in_data_full_n;
wire    dataflow_in_loop_TOP_LOOP37454_U0_in_data_write;
wire    ap_sync_continue;
wire    ap_sync_done;
wire    ap_sync_ready;
reg   [17:0] loop_dataflow_input_count;
reg   [17:0] loop_dataflow_output_count;
wire   [17:0] bound_minus_1;
wire    dataflow_in_loop_TOP_LOOP37454_U0_start_full_n;
wire    dataflow_in_loop_TOP_LOOP37454_U0_start_write;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 loop_dataflow_input_count = 18'd0;
#0 loop_dataflow_output_count = 18'd0;
end

td_fused_top_dataflow_in_loop_TOP_LOOP37454 dataflow_in_loop_TOP_LOOP37454_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .in_data_address0(dataflow_in_loop_TOP_LOOP37454_U0_in_data_address0),
    .in_data_ce0(dataflow_in_loop_TOP_LOOP37454_U0_in_data_ce0),
    .in_data_d0(dataflow_in_loop_TOP_LOOP37454_U0_in_data_d0),
    .in_data_q0(in_data_q0),
    .in_data_we0(dataflow_in_loop_TOP_LOOP37454_U0_in_data_we0),
    .in_data_address1(dataflow_in_loop_TOP_LOOP37454_U0_in_data_address1),
    .in_data_ce1(dataflow_in_loop_TOP_LOOP37454_U0_in_data_ce1),
    .in_data_d1(dataflow_in_loop_TOP_LOOP37454_U0_in_data_d1),
    .in_data_q1(64'd0),
    .in_data_we1(dataflow_in_loop_TOP_LOOP37454_U0_in_data_we1),
    .filter_data_address0(dataflow_in_loop_TOP_LOOP37454_U0_filter_data_address0),
    .filter_data_ce0(dataflow_in_loop_TOP_LOOP37454_U0_filter_data_ce0),
    .filter_data_d0(dataflow_in_loop_TOP_LOOP37454_U0_filter_data_d0),
    .filter_data_q0(filter_data_q0),
    .filter_data_we0(dataflow_in_loop_TOP_LOOP37454_U0_filter_data_we0),
    .filter_data_address1(dataflow_in_loop_TOP_LOOP37454_U0_filter_data_address1),
    .filter_data_ce1(dataflow_in_loop_TOP_LOOP37454_U0_filter_data_ce1),
    .filter_data_d1(dataflow_in_loop_TOP_LOOP37454_U0_filter_data_d1),
    .filter_data_q1(16'd0),
    .filter_data_we1(dataflow_in_loop_TOP_LOOP37454_U0_filter_data_we1),
    .adjustments_address0(dataflow_in_loop_TOP_LOOP37454_U0_adjustments_address0),
    .adjustments_ce0(dataflow_in_loop_TOP_LOOP37454_U0_adjustments_ce0),
    .adjustments_d0(dataflow_in_loop_TOP_LOOP37454_U0_adjustments_d0),
    .adjustments_q0(adjustments_q0),
    .adjustments_we0(dataflow_in_loop_TOP_LOOP37454_U0_adjustments_we0),
    .adjustments_address1(dataflow_in_loop_TOP_LOOP37454_U0_adjustments_address1),
    .adjustments_ce1(dataflow_in_loop_TOP_LOOP37454_U0_adjustments_ce1),
    .adjustments_d1(dataflow_in_loop_TOP_LOOP37454_U0_adjustments_d1),
    .adjustments_q1(48'd0),
    .adjustments_we1(dataflow_in_loop_TOP_LOOP37454_U0_adjustments_we1),
    .out_data_address0(dataflow_in_loop_TOP_LOOP37454_U0_out_data_address0),
    .out_data_ce0(dataflow_in_loop_TOP_LOOP37454_U0_out_data_ce0),
    .out_data_d0(dataflow_in_loop_TOP_LOOP37454_U0_out_data_d0),
    .out_data_q0(64'd0),
    .out_data_we0(dataflow_in_loop_TOP_LOOP37454_U0_out_data_we0),
    .out_data_address1(dataflow_in_loop_TOP_LOOP37454_U0_out_data_address1),
    .out_data_ce1(dataflow_in_loop_TOP_LOOP37454_U0_out_data_ce1),
    .out_data_d1(dataflow_in_loop_TOP_LOOP37454_U0_out_data_d1),
    .out_data_q1(64'd0),
    .out_data_we1(dataflow_in_loop_TOP_LOOP37454_U0_out_data_we1),
    .ap_start(dataflow_in_loop_TOP_LOOP37454_U0_ap_start),
    .in_data_empty_n(1'b0),
    .in_data_read(dataflow_in_loop_TOP_LOOP37454_U0_in_data_read),
    .out_data_full_n(out_data_full_n),
    .out_data_write(dataflow_in_loop_TOP_LOOP37454_U0_out_data_write),
    .ap_done(dataflow_in_loop_TOP_LOOP37454_U0_ap_done),
    .ap_ready(dataflow_in_loop_TOP_LOOP37454_U0_ap_ready),
    .ap_idle(dataflow_in_loop_TOP_LOOP37454_U0_ap_idle),
    .ap_continue(dataflow_in_loop_TOP_LOOP37454_U0_ap_continue)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        loop_dataflow_input_count <= 18'd0;
    end else begin
        if ((~(loop_dataflow_input_count == bound_minus_1) & (dataflow_in_loop_TOP_LOOP37454_U0_ap_ready == 1'b1) & (ap_start == 1'b1))) begin
            loop_dataflow_input_count <= (loop_dataflow_input_count + 18'd1);
        end else if (((dataflow_in_loop_TOP_LOOP37454_U0_ap_ready == 1'b1) & (loop_dataflow_input_count == bound_minus_1) & (ap_start == 1'b1))) begin
            loop_dataflow_input_count <= 18'd0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        loop_dataflow_output_count <= 18'd0;
    end else begin
        if ((~(loop_dataflow_output_count == bound_minus_1) & (dataflow_in_loop_TOP_LOOP37454_U0_ap_done == 1'b1) & (dataflow_in_loop_TOP_LOOP37454_U0_ap_continue == 1'b1))) begin
            loop_dataflow_output_count <= (loop_dataflow_output_count + 18'd1);
        end else if (((dataflow_in_loop_TOP_LOOP37454_U0_ap_done == 1'b1) & (loop_dataflow_output_count == bound_minus_1) & (dataflow_in_loop_TOP_LOOP37454_U0_ap_continue == 1'b1))) begin
            loop_dataflow_output_count <= 18'd0;
        end
    end
end

always @ (*) begin
    if (((dataflow_in_loop_TOP_LOOP37454_U0_ap_done == 1'b1) & (loop_dataflow_output_count == bound_minus_1))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = 1'b0;
    end
end

always @ (*) begin
    if (((dataflow_in_loop_TOP_LOOP37454_U0_ap_idle == 1'b1) & (loop_dataflow_output_count == 18'd0) & (ap_start == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((dataflow_in_loop_TOP_LOOP37454_U0_ap_ready == 1'b1) & (loop_dataflow_input_count == bound_minus_1) & (ap_start == 1'b1))) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((~(loop_dataflow_output_count == bound_minus_1) | (ap_continue == 1'b1))) begin
        dataflow_in_loop_TOP_LOOP37454_U0_ap_continue = 1'b1;
    end else begin
        dataflow_in_loop_TOP_LOOP37454_U0_ap_continue = 1'b0;
    end
end

assign adjustments_address0 = dataflow_in_loop_TOP_LOOP37454_U0_adjustments_address0;

assign adjustments_address1 = 8'd0;

assign adjustments_ce0 = dataflow_in_loop_TOP_LOOP37454_U0_adjustments_ce0;

assign adjustments_ce1 = 1'b0;

assign adjustments_d0 = 48'd0;

assign adjustments_d1 = 48'd0;

assign adjustments_we0 = 1'b0;

assign adjustments_we1 = 1'b0;

assign ap_sync_continue = ap_continue;

assign ap_sync_done = dataflow_in_loop_TOP_LOOP37454_U0_ap_done;

assign ap_sync_ready = dataflow_in_loop_TOP_LOOP37454_U0_ap_ready;

assign bound_minus_1 = (18'd200704 - 18'd1);

assign dataflow_in_loop_TOP_LOOP37454_U0_ap_start = ap_start;

assign dataflow_in_loop_TOP_LOOP37454_U0_in_data_full_n = in_data_empty_n;

assign dataflow_in_loop_TOP_LOOP37454_U0_in_data_write = 1'b0;

assign dataflow_in_loop_TOP_LOOP37454_U0_start_full_n = 1'b1;

assign dataflow_in_loop_TOP_LOOP37454_U0_start_write = 1'b0;

assign filter_data_address0 = dataflow_in_loop_TOP_LOOP37454_U0_filter_data_address0;

assign filter_data_address1 = 17'd0;

assign filter_data_ce0 = dataflow_in_loop_TOP_LOOP37454_U0_filter_data_ce0;

assign filter_data_ce1 = 1'b0;

assign filter_data_d0 = 16'd0;

assign filter_data_d1 = 16'd0;

assign filter_data_we0 = 1'b0;

assign filter_data_we1 = 1'b0;

assign in_data_address0 = dataflow_in_loop_TOP_LOOP37454_U0_in_data_address0;

assign in_data_address1 = 13'd0;

assign in_data_ce0 = dataflow_in_loop_TOP_LOOP37454_U0_in_data_ce0;

assign in_data_ce1 = 1'b0;

assign in_data_d0 = 64'd0;

assign in_data_d1 = 64'd0;

assign in_data_read = dataflow_in_loop_TOP_LOOP37454_U0_in_data_write;

assign in_data_we0 = 1'b0;

assign in_data_we1 = 1'b0;

assign out_data_address0 = 14'd0;

assign out_data_address1 = dataflow_in_loop_TOP_LOOP37454_U0_out_data_address1;

assign out_data_ce0 = 1'b0;

assign out_data_ce1 = dataflow_in_loop_TOP_LOOP37454_U0_out_data_ce1;

assign out_data_d0 = 64'd0;

assign out_data_d1 = dataflow_in_loop_TOP_LOOP37454_U0_out_data_d1;

assign out_data_we0 = 1'b0;

assign out_data_we1 = dataflow_in_loop_TOP_LOOP37454_U0_out_data_we1;

assign out_data_write = dataflow_in_loop_TOP_LOOP37454_U0_out_data_write;

endmodule //td_fused_top_tdf8_17
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf8_accum_1 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        accum_in_0_address0,
        accum_in_0_ce0,
        accum_in_0_q0,
        accum_in_0_address1,
        accum_in_0_ce1,
        accum_in_0_q1,
        accum_out_address0,
        accum_out_ce0,
        accum_out_we0,
        accum_out_d0,
        accum_out_address1,
        accum_out_ce1,
        accum_out_we1,
        accum_out_d1
);

parameter    ap_ST_fsm_state1 = 8'd1;
parameter    ap_ST_fsm_pp0_stage0 = 8'd2;
parameter    ap_ST_fsm_pp0_stage1 = 8'd4;
parameter    ap_ST_fsm_pp0_stage2 = 8'd8;
parameter    ap_ST_fsm_pp0_stage3 = 8'd16;
parameter    ap_ST_fsm_state12 = 8'd32;
parameter    ap_ST_fsm_state13 = 8'd64;
parameter    ap_ST_fsm_state14 = 8'd128;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [8:0] accum_in_0_address0;
output   accum_in_0_ce0;
input  [15:0] accum_in_0_q0;
output  [8:0] accum_in_0_address1;
output   accum_in_0_ce1;
input  [15:0] accum_in_0_q1;
output  [2:0] accum_out_address0;
output   accum_out_ce0;
output   accum_out_we0;
output  [15:0] accum_out_d0;
output  [2:0] accum_out_address1;
output   accum_out_ce1;
output   accum_out_we1;
output  [15:0] accum_out_d1;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg[8:0] accum_in_0_address0;
reg accum_in_0_ce0;
reg[8:0] accum_in_0_address1;
reg accum_in_0_ce1;
reg accum_out_ce0;
reg accum_out_we0;
reg accum_out_ce1;
reg accum_out_we1;

reg    ap_done_reg;
  reg   [7:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg   [8:0] x_reg_168;
reg   [15:0] psum_7_08_reg_180;
reg   [15:0] psum_6_07_reg_192;
reg   [15:0] psum_5_06_reg_204;
reg   [15:0] psum_4_05_reg_216;
reg   [15:0] psum_3_04_reg_228;
reg   [15:0] psum_2_03_reg_240;
reg   [15:0] psum_1_02_reg_252;
reg   [15:0] psum_0_01_reg_264;
wire   [0:0] icmp_ln49_fu_321_p2;
reg   [0:0] icmp_ln49_reg_492;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state6_pp0_stage0_iter1;
wire    ap_block_state10_pp0_stage0_iter2;
wire    ap_block_pp0_stage0_11001;
reg   [0:0] icmp_ln49_reg_492_pp0_iter1_reg;
reg   [0:0] icmp_ln49_reg_492_pp0_iter2_reg;
reg   [15:0] accum_in_0_load_reg_506;
wire    ap_CS_fsm_pp0_stage1;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_state3_pp0_stage1_iter0;
wire    ap_block_state7_pp0_stage1_iter1;
wire    ap_block_state11_pp0_stage1_iter2;
wire    ap_block_pp0_stage1_11001;
reg   [15:0] accum_in_0_load_8_reg_511;
reg   [15:0] accum_in_0_load_9_reg_526;
wire    ap_CS_fsm_pp0_stage2;
wire    ap_block_state4_pp0_stage2_iter0;
wire    ap_block_state8_pp0_stage2_iter1;
wire    ap_block_pp0_stage2_11001;
reg   [15:0] accum_in_0_load_10_reg_531;
wire   [8:0] add_ln49_fu_387_p2;
reg   [8:0] add_ln49_reg_546;
wire    ap_CS_fsm_pp0_stage3;
wire    ap_block_state5_pp0_stage3_iter0;
wire    ap_block_state9_pp0_stage3_iter1;
wire    ap_block_pp0_stage3_11001;
reg   [15:0] accum_in_0_load_11_reg_551;
reg   [15:0] accum_in_0_load_12_reg_556;
reg   [15:0] accum_in_0_load_13_reg_571;
reg    ap_enable_reg_pp0_iter1;
reg   [15:0] accum_in_0_load_14_reg_576;
wire   [15:0] grp_fu_305_p2;
wire   [15:0] grp_fu_310_p2;
reg    ap_enable_reg_pp0_iter2;
wire   [3:0] add_ln57_fu_432_p2;
wire    ap_CS_fsm_state13;
wire   [0:0] tmp_fu_415_p3;
reg    ap_block_state1;
wire    ap_block_pp0_stage2_subdone;
reg    ap_condition_pp0_exit_iter0_state4;
wire    ap_block_pp0_stage3_subdone;
wire    ap_block_pp0_stage1_subdone;
reg   [8:0] ap_phi_mux_x_phi_fu_172_p4;
wire    ap_block_pp0_stage0;
wire   [15:0] ap_phi_mux_psum_7_08_phi_fu_184_p4;
wire    ap_block_pp0_stage1;
wire   [15:0] ap_phi_mux_psum_6_07_phi_fu_196_p4;
wire   [15:0] ap_phi_mux_psum_5_06_phi_fu_208_p4;
wire   [15:0] ap_phi_mux_psum_4_05_phi_fu_220_p4;
wire   [15:0] ap_phi_mux_psum_3_04_phi_fu_232_p4;
wire    ap_block_pp0_stage3;
wire   [15:0] ap_phi_mux_psum_2_03_phi_fu_244_p4;
wire    ap_block_pp0_stage2;
reg   [3:0] q_reg_276;
wire    ap_CS_fsm_state12;
reg   [15:0] ap_phi_mux_phi_ln69_phi_fu_290_p8;
wire   [2:0] trunc_ln57_fu_428_p1;
wire   [63:0] zext_ln49_fu_327_p1;
wire   [63:0] zext_ln53_fu_338_p1;
wire   [63:0] zext_ln53_1_fu_349_p1;
wire   [63:0] zext_ln53_2_fu_360_p1;
wire   [63:0] zext_ln53_3_fu_371_p1;
wire   [63:0] zext_ln53_4_fu_382_p1;
wire   [63:0] zext_ln53_5_fu_399_p1;
wire   [63:0] zext_ln53_6_fu_410_p1;
wire   [63:0] zext_ln57_fu_423_p1;
wire   [63:0] zext_ln57_1_fu_444_p1;
reg   [15:0] grp_fu_305_p0;
reg   [15:0] grp_fu_305_p1;
reg   [15:0] grp_fu_310_p0;
reg   [15:0] grp_fu_310_p1;
wire   [8:0] or_ln53_fu_332_p2;
wire   [8:0] or_ln53_1_fu_343_p2;
wire   [8:0] or_ln53_2_fu_354_p2;
wire   [8:0] or_ln53_3_fu_365_p2;
wire   [8:0] or_ln53_4_fu_376_p2;
wire   [8:0] or_ln53_5_fu_393_p2;
wire   [8:0] or_ln53_6_fu_404_p2;
wire   [2:0] or_ln57_fu_438_p2;
wire   [0:0] icmp_ln69_fu_449_p2;
wire   [0:0] icmp_ln69_1_fu_463_p2;
wire   [15:0] select_ln69_fu_455_p3;
wire   [0:0] icmp_ln69_2_fu_477_p2;
wire   [15:0] select_ln69_1_fu_469_p3;
wire    ap_CS_fsm_state14;
reg   [7:0] ap_NS_fsm;
wire    ap_block_pp0_stage0_subdone;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
reg    ap_condition_514;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 8'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
end

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U498(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(grp_fu_305_p0),
    .din1(grp_fu_305_p1),
    .dout(grp_fu_305_p2)
);

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U499(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(grp_fu_310_p0),
    .din1(grp_fu_310_p1),
    .dout(grp_fu_310_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state14)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage2_subdone) & (1'b1 == ap_condition_pp0_exit_iter0_state4) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage3_subdone) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b0)) | ((1'b0 == ap_block_pp0_stage3_subdone) & (1'b1 == ap_CS_fsm_pp0_stage3)))) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end else if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter2 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state12)) begin
        q_reg_276 <= 4'd0;
    end else if (((tmp_fu_415_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state13))) begin
        q_reg_276 <= add_ln57_fu_432_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln49_reg_492 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        x_reg_168 <= add_ln49_reg_546;
    end else if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        x_reg_168 <= 9'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2_11001) & (icmp_ln49_reg_492 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
        accum_in_0_load_10_reg_531 <= accum_in_0_q0;
        accum_in_0_load_9_reg_526 <= accum_in_0_q1;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage3_11001) & (icmp_ln49_reg_492 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
        accum_in_0_load_11_reg_551 <= accum_in_0_q1;
        accum_in_0_load_12_reg_556 <= accum_in_0_q0;
        add_ln49_reg_546 <= add_ln49_fu_387_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (icmp_ln49_reg_492 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        accum_in_0_load_13_reg_571 <= accum_in_0_q1;
        accum_in_0_load_14_reg_576 <= accum_in_0_q0;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage1_11001) & (icmp_ln49_reg_492 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
        accum_in_0_load_8_reg_511 <= accum_in_0_q0;
        accum_in_0_load_reg_506 <= accum_in_0_q1;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln49_reg_492 <= icmp_ln49_fu_321_p2;
        icmp_ln49_reg_492_pp0_iter1_reg <= icmp_ln49_reg_492;
        icmp_ln49_reg_492_pp0_iter2_reg <= icmp_ln49_reg_492_pp0_iter1_reg;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln49_reg_492_pp0_iter1_reg == 1'd1) & (1'b0 == ap_block_pp0_stage2_11001) & (1'b1 == ap_CS_fsm_pp0_stage2) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        psum_0_01_reg_264 <= grp_fu_305_p2;
        psum_1_02_reg_252 <= grp_fu_310_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln49_reg_492_pp0_iter1_reg == 1'd1) & (1'b0 == ap_block_pp0_stage3_11001) & (1'b1 == ap_CS_fsm_pp0_stage3) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        psum_2_03_reg_240 <= grp_fu_305_p2;
        psum_3_04_reg_228 <= grp_fu_310_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln49_reg_492_pp0_iter1_reg == 1'd1) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        psum_4_05_reg_216 <= grp_fu_305_p2;
        psum_5_06_reg_204 <= grp_fu_310_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln49_reg_492_pp0_iter2_reg == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        psum_6_07_reg_192 <= grp_fu_305_p2;
        psum_7_08_reg_180 <= grp_fu_310_p2;
    end
end

always @ (*) begin
    if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
        if (((1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            accum_in_0_address0 = zext_ln53_6_fu_410_p1;
        end else if (((1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            accum_in_0_address0 = zext_ln53_4_fu_382_p1;
        end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            accum_in_0_address0 = zext_ln53_2_fu_360_p1;
        end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            accum_in_0_address0 = zext_ln53_fu_338_p1;
        end else begin
            accum_in_0_address0 = 'bx;
        end
    end else begin
        accum_in_0_address0 = 'bx;
    end
end

always @ (*) begin
    if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
        if (((1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            accum_in_0_address1 = zext_ln53_5_fu_399_p1;
        end else if (((1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            accum_in_0_address1 = zext_ln53_3_fu_371_p1;
        end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            accum_in_0_address1 = zext_ln53_1_fu_349_p1;
        end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            accum_in_0_address1 = zext_ln49_fu_327_p1;
        end else begin
            accum_in_0_address1 = 'bx;
        end
    end else begin
        accum_in_0_address1 = 'bx;
    end
end

always @ (*) begin
    if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage3_11001) & (1'b1 == ap_CS_fsm_pp0_stage3)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2_11001) & (1'b1 == ap_CS_fsm_pp0_stage2)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1)))) begin
        accum_in_0_ce0 = 1'b1;
    end else begin
        accum_in_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage3_11001) & (1'b1 == ap_CS_fsm_pp0_stage3)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2_11001) & (1'b1 == ap_CS_fsm_pp0_stage2)) | ((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1)))) begin
        accum_in_0_ce1 = 1'b1;
    end else begin
        accum_in_0_ce1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state13)) begin
        accum_out_ce0 = 1'b1;
    end else begin
        accum_out_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state13)) begin
        accum_out_ce1 = 1'b1;
    end else begin
        accum_out_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((tmp_fu_415_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state13))) begin
        accum_out_we0 = 1'b1;
    end else begin
        accum_out_we0 = 1'b0;
    end
end

always @ (*) begin
    if (((tmp_fu_415_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state13))) begin
        accum_out_we1 = 1'b1;
    end else begin
        accum_out_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((icmp_ln49_reg_492 == 1'd0)) begin
        ap_condition_pp0_exit_iter0_state4 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state4 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state14)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((tmp_fu_415_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state13))) begin
        if ((trunc_ln57_fu_428_p1 == 3'd0)) begin
            ap_phi_mux_phi_ln69_phi_fu_290_p8 = psum_0_01_reg_264;
        end else if ((1'b1 == ap_condition_514)) begin
            ap_phi_mux_phi_ln69_phi_fu_290_p8 = psum_6_07_reg_192;
        end else if ((trunc_ln57_fu_428_p1 == 3'd4)) begin
            ap_phi_mux_phi_ln69_phi_fu_290_p8 = psum_4_05_reg_216;
        end else if ((trunc_ln57_fu_428_p1 == 3'd2)) begin
            ap_phi_mux_phi_ln69_phi_fu_290_p8 = psum_2_03_reg_240;
        end else begin
            ap_phi_mux_phi_ln69_phi_fu_290_p8 = 'bx;
        end
    end else begin
        ap_phi_mux_phi_ln69_phi_fu_290_p8 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0) & (icmp_ln49_reg_492 == 1'd1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_x_phi_fu_172_p4 = add_ln49_reg_546;
    end else begin
        ap_phi_mux_x_phi_fu_172_p4 = x_reg_168;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state14)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_305_p0 = ap_phi_mux_psum_6_07_phi_fu_196_p4;
    end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_305_p0 = ap_phi_mux_psum_4_05_phi_fu_220_p4;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
        grp_fu_305_p0 = ap_phi_mux_psum_2_03_phi_fu_244_p4;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
        grp_fu_305_p0 = grp_fu_305_p2;
    end else begin
        grp_fu_305_p0 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_305_p1 = accum_in_0_load_13_reg_571;
    end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_305_p1 = accum_in_0_load_11_reg_551;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
        grp_fu_305_p1 = accum_in_0_load_9_reg_526;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
        grp_fu_305_p1 = accum_in_0_load_reg_506;
    end else begin
        grp_fu_305_p1 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_310_p0 = ap_phi_mux_psum_7_08_phi_fu_184_p4;
    end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_310_p0 = ap_phi_mux_psum_5_06_phi_fu_208_p4;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
        grp_fu_310_p0 = ap_phi_mux_psum_3_04_phi_fu_232_p4;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
        grp_fu_310_p0 = grp_fu_310_p2;
    end else begin
        grp_fu_310_p0 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_310_p1 = accum_in_0_load_14_reg_576;
    end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_310_p1 = accum_in_0_load_12_reg_556;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
        grp_fu_310_p1 = accum_in_0_load_10_reg_531;
    end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
        grp_fu_310_p1 = accum_in_0_load_8_reg_511;
    end else begin
        grp_fu_310_p1 = 'bx;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_pp0_stage1 : begin
            if ((~((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter2 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0)) & (1'b0 == ap_block_pp0_stage1_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage2;
            end else if (((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter2 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
                ap_NS_fsm = ap_ST_fsm_state12;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end
        end
        ap_ST_fsm_pp0_stage2 : begin
            if ((~((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2_subdone) & (icmp_ln49_reg_492 == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b0)) & (1'b0 == ap_block_pp0_stage2_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage3;
            end else if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage2_subdone) & (icmp_ln49_reg_492 == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
                ap_NS_fsm = ap_ST_fsm_state12;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage2;
            end
        end
        ap_ST_fsm_pp0_stage3 : begin
            if ((1'b0 == ap_block_pp0_stage3_subdone)) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage3;
            end
        end
        ap_ST_fsm_state12 : begin
            ap_NS_fsm = ap_ST_fsm_state13;
        end
        ap_ST_fsm_state13 : begin
            if (((tmp_fu_415_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state13))) begin
                ap_NS_fsm = ap_ST_fsm_state13;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state14;
            end
        end
        ap_ST_fsm_state14 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign accum_out_address0 = zext_ln57_1_fu_444_p1;

assign accum_out_address1 = zext_ln57_fu_423_p1;

assign accum_out_d0 = ((icmp_ln69_2_fu_477_p2[0:0] == 1'b1) ? psum_5_06_reg_204 : select_ln69_1_fu_469_p3);

assign accum_out_d1 = ap_phi_mux_phi_ln69_phi_fu_290_p8;

assign add_ln49_fu_387_p2 = (x_reg_168 + 9'd8);

assign add_ln57_fu_432_p2 = (q_reg_276 + 4'd2);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_pp0_stage1 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_pp0_stage2 = ap_CS_fsm[32'd3];

assign ap_CS_fsm_pp0_stage3 = ap_CS_fsm[32'd4];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state12 = ap_CS_fsm[32'd5];

assign ap_CS_fsm_state13 = ap_CS_fsm[32'd6];

assign ap_CS_fsm_state14 = ap_CS_fsm[32'd7];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1_subdone = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage2 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage2_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage2_subdone = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage3 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage3_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage3_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((ap_done_reg == 1'b1) | (ap_start == 1'b0));
end

assign ap_block_state10_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state11_pp0_stage1_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage1_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage2_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage3_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage1_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage2_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state9_pp0_stage3_iter1 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_condition_514 = (~(trunc_ln57_fu_428_p1 == 3'd0) & ~(trunc_ln57_fu_428_p1 == 3'd4) & ~(trunc_ln57_fu_428_p1 == 3'd2));
end

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign ap_phi_mux_psum_2_03_phi_fu_244_p4 = grp_fu_305_p2;

assign ap_phi_mux_psum_3_04_phi_fu_232_p4 = grp_fu_310_p2;

assign ap_phi_mux_psum_4_05_phi_fu_220_p4 = grp_fu_305_p2;

assign ap_phi_mux_psum_5_06_phi_fu_208_p4 = grp_fu_310_p2;

assign ap_phi_mux_psum_6_07_phi_fu_196_p4 = grp_fu_305_p2;

assign ap_phi_mux_psum_7_08_phi_fu_184_p4 = grp_fu_310_p2;

assign icmp_ln49_fu_321_p2 = ((ap_phi_mux_x_phi_fu_172_p4 < 9'd288) ? 1'b1 : 1'b0);

assign icmp_ln69_1_fu_463_p2 = ((or_ln57_fu_438_p2 == 3'd3) ? 1'b1 : 1'b0);

assign icmp_ln69_2_fu_477_p2 = ((or_ln57_fu_438_p2 == 3'd5) ? 1'b1 : 1'b0);

assign icmp_ln69_fu_449_p2 = ((or_ln57_fu_438_p2 == 3'd1) ? 1'b1 : 1'b0);

assign or_ln53_1_fu_343_p2 = (x_reg_168 | 9'd2);

assign or_ln53_2_fu_354_p2 = (x_reg_168 | 9'd3);

assign or_ln53_3_fu_365_p2 = (x_reg_168 | 9'd4);

assign or_ln53_4_fu_376_p2 = (x_reg_168 | 9'd5);

assign or_ln53_5_fu_393_p2 = (x_reg_168 | 9'd6);

assign or_ln53_6_fu_404_p2 = (x_reg_168 | 9'd7);

assign or_ln53_fu_332_p2 = (ap_phi_mux_x_phi_fu_172_p4 | 9'd1);

assign or_ln57_fu_438_p2 = (trunc_ln57_fu_428_p1 | 3'd1);

assign select_ln69_1_fu_469_p3 = ((icmp_ln69_1_fu_463_p2[0:0] == 1'b1) ? psum_3_04_reg_228 : select_ln69_fu_455_p3);

assign select_ln69_fu_455_p3 = ((icmp_ln69_fu_449_p2[0:0] == 1'b1) ? psum_1_02_reg_252 : psum_7_08_reg_180);

assign tmp_fu_415_p3 = q_reg_276[32'd3];

assign trunc_ln57_fu_428_p1 = q_reg_276[2:0];

assign zext_ln49_fu_327_p1 = ap_phi_mux_x_phi_fu_172_p4;

assign zext_ln53_1_fu_349_p1 = or_ln53_1_fu_343_p2;

assign zext_ln53_2_fu_360_p1 = or_ln53_2_fu_354_p2;

assign zext_ln53_3_fu_371_p1 = or_ln53_3_fu_365_p2;

assign zext_ln53_4_fu_382_p1 = or_ln53_4_fu_376_p2;

assign zext_ln53_5_fu_399_p1 = or_ln53_5_fu_393_p2;

assign zext_ln53_6_fu_410_p1 = or_ln53_6_fu_404_p2;

assign zext_ln53_fu_338_p1 = or_ln53_fu_332_p2;

assign zext_ln57_1_fu_444_p1 = or_ln57_fu_438_p2;

assign zext_ln57_fu_423_p1 = q_reg_276;

endmodule //td_fused_top_tdf8_accum_1
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf8_accum_2 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        accum_in_4,
        accum_in_4_ap_vld,
        accum_in_address0,
        accum_in_ce0,
        accum_in_q0
);

parameter    ap_ST_fsm_state1 = 7'd1;
parameter    ap_ST_fsm_state2 = 7'd2;
parameter    ap_ST_fsm_state3 = 7'd4;
parameter    ap_ST_fsm_state4 = 7'd8;
parameter    ap_ST_fsm_state5 = 7'd16;
parameter    ap_ST_fsm_state6 = 7'd32;
parameter    ap_ST_fsm_state7 = 7'd64;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [15:0] accum_in_4;
output   accum_in_4_ap_vld;
output  [2:0] accum_in_address0;
output   accum_in_ce0;
input  [15:0] accum_in_q0;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg[15:0] accum_in_4;
reg accum_in_4_ap_vld;
reg accum_in_ce0;

reg    ap_done_reg;
  reg   [6:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
wire   [3:0] add_ln81_fu_74_p2;
reg   [3:0] add_ln81_reg_91;
wire    ap_CS_fsm_state2;
wire   [0:0] icmp_ln81_fu_85_p2;
wire    ap_CS_fsm_state3;
wire   [15:0] grp_fu_68_p2;
wire    ap_CS_fsm_state7;
reg   [3:0] i_1_1_reg_44;
reg    ap_block_state1;
reg   [15:0] sum_01_reg_55;
wire   [63:0] zext_ln81_fu_80_p1;
reg   [15:0] accum_in_4_preg;
reg   [6:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 7'd1;
#0 accum_in_4_preg = 16'd0;
end

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U502(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(sum_01_reg_55),
    .din1(accum_in_q0),
    .dout(grp_fu_68_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        accum_in_4_preg <= 16'd0;
    end else begin
        if (((icmp_ln81_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
            accum_in_4_preg <= sum_01_reg_55;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if (((icmp_ln81_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        i_1_1_reg_44 <= 4'd0;
    end else if ((1'b1 == ap_CS_fsm_state7)) begin
        i_1_1_reg_44 <= add_ln81_reg_91;
    end
end

always @ (posedge ap_clk) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        sum_01_reg_55 <= 16'd0;
    end else if ((1'b1 == ap_CS_fsm_state7)) begin
        sum_01_reg_55 <= grp_fu_68_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        add_ln81_reg_91 <= add_ln81_fu_74_p2;
    end
end

always @ (*) begin
    if (((icmp_ln81_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        accum_in_4 = sum_01_reg_55;
    end else begin
        accum_in_4 = accum_in_4_preg;
    end
end

always @ (*) begin
    if (((icmp_ln81_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        accum_in_4_ap_vld = 1'b1;
    end else begin
        accum_in_4_ap_vld = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        accum_in_ce0 = 1'b1;
    end else begin
        accum_in_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln81_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln81_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_state2 : begin
            if (((icmp_ln81_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end
        end
        ap_ST_fsm_state3 : begin
            ap_NS_fsm = ap_ST_fsm_state4;
        end
        ap_ST_fsm_state4 : begin
            ap_NS_fsm = ap_ST_fsm_state5;
        end
        ap_ST_fsm_state5 : begin
            ap_NS_fsm = ap_ST_fsm_state6;
        end
        ap_ST_fsm_state6 : begin
            ap_NS_fsm = ap_ST_fsm_state7;
        end
        ap_ST_fsm_state7 : begin
            ap_NS_fsm = ap_ST_fsm_state2;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign accum_in_address0 = zext_ln81_fu_80_p1;

assign add_ln81_fu_74_p2 = (i_1_1_reg_44 + 4'd1);

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state7 = ap_CS_fsm[32'd6];

always @ (*) begin
    ap_block_state1 = ((ap_done_reg == 1'b1) | (ap_start == 1'b0));
end

assign icmp_ln81_fu_85_p2 = ((i_1_1_reg_44 == 4'd8) ? 1'b1 : 1'b0);

assign zext_ln81_fu_80_p1 = i_1_1_reg_44;

endmodule //td_fused_top_tdf8_accum_2
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf8_adjust (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        sums_read,
        adjustments_address0,
        adjustments_ce0,
        adjustments_q0,
        input_indices_23_dout,
        input_indices_23_empty_n,
        input_indices_23_read,
        ap_return
);

parameter    ap_ST_fsm_state1 = 17'd1;
parameter    ap_ST_fsm_state2 = 17'd2;
parameter    ap_ST_fsm_state3 = 17'd4;
parameter    ap_ST_fsm_state4 = 17'd8;
parameter    ap_ST_fsm_state5 = 17'd16;
parameter    ap_ST_fsm_state6 = 17'd32;
parameter    ap_ST_fsm_state7 = 17'd64;
parameter    ap_ST_fsm_state8 = 17'd128;
parameter    ap_ST_fsm_state9 = 17'd256;
parameter    ap_ST_fsm_state10 = 17'd512;
parameter    ap_ST_fsm_state11 = 17'd1024;
parameter    ap_ST_fsm_state12 = 17'd2048;
parameter    ap_ST_fsm_state13 = 17'd4096;
parameter    ap_ST_fsm_state14 = 17'd8192;
parameter    ap_ST_fsm_state15 = 17'd16384;
parameter    ap_ST_fsm_state16 = 17'd32768;
parameter    ap_ST_fsm_state17 = 17'd65536;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
input  [15:0] sums_read;
output  [7:0] adjustments_address0;
output   adjustments_ce0;
input  [47:0] adjustments_q0;
input  [7:0] input_indices_23_dout;
input   input_indices_23_empty_n;
output   input_indices_23_read;
output  [15:0] ap_return;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg adjustments_ce0;
reg input_indices_23_read;

reg    ap_done_reg;
  reg   [16:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    input_indices_23_blk_n;
wire    ap_CS_fsm_state4;
reg   [15:0] tmp_15_i_i_reg_167;
reg   [15:0] tmp_16_i_i_reg_172;
wire   [15:0] grp_fu_81_p2;
reg   [15:0] sub_i_i_i_reg_177;
wire    ap_CS_fsm_state8;
wire    ap_CS_fsm_state9;
wire   [15:0] grp_fu_86_p2;
reg   [15:0] mul_i_i_i_reg_187;
wire    ap_CS_fsm_state12;
wire    ap_CS_fsm_state13;
wire   [63:0] zext_ln220_fu_90_p1;
reg    ap_block_state1;
wire    ap_CS_fsm_state2;
wire    ap_CS_fsm_state3;
wire   [15:0] grp_fu_77_p1;
wire   [15:0] grp_fu_81_p1;
wire   [15:0] grp_fu_86_p1;
wire   [15:0] trunc_ln220_fu_95_p1;
wire   [15:0] grp_fu_77_p2;
wire    ap_CS_fsm_state17;
wire   [15:0] bitcast_ln648_fu_132_p1;
wire   [0:0] tmp_fu_136_p3;
reg   [16:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 17'd1;
end

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U506(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(mul_i_i_i_reg_187),
    .din1(grp_fu_77_p1),
    .dout(grp_fu_77_p2)
);

td_fused_top_hsub_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hsub_16ns_16ns_16_5_full_dsp_1_U507(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(sums_read),
    .din1(grp_fu_81_p1),
    .dout(grp_fu_81_p2)
);

td_fused_top_hmul_16ns_16ns_16_4_max_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hmul_16ns_16ns_16_4_max_dsp_1_U508(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(sub_i_i_i_reg_177),
    .din1(grp_fu_86_p1),
    .dout(grp_fu_86_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state17)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state12)) begin
        mul_i_i_i_reg_187 <= grp_fu_86_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state8)) begin
        sub_i_i_i_reg_177 <= grp_fu_81_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        tmp_15_i_i_reg_167 <= {{adjustments_q0[31:16]}};
        tmp_16_i_i_reg_172 <= {{adjustments_q0[47:32]}};
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state2) | (~((input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1)))) begin
        adjustments_ce0 = 1'b1;
    end else begin
        adjustments_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state17)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state17)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        input_indices_23_blk_n = input_indices_23_empty_n;
    end else begin
        input_indices_23_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        input_indices_23_read = 1'b1;
    end else begin
        input_indices_23_read = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_state2 : begin
            ap_NS_fsm = ap_ST_fsm_state3;
        end
        ap_ST_fsm_state3 : begin
            ap_NS_fsm = ap_ST_fsm_state4;
        end
        ap_ST_fsm_state4 : begin
            ap_NS_fsm = ap_ST_fsm_state5;
        end
        ap_ST_fsm_state5 : begin
            ap_NS_fsm = ap_ST_fsm_state6;
        end
        ap_ST_fsm_state6 : begin
            ap_NS_fsm = ap_ST_fsm_state7;
        end
        ap_ST_fsm_state7 : begin
            ap_NS_fsm = ap_ST_fsm_state8;
        end
        ap_ST_fsm_state8 : begin
            ap_NS_fsm = ap_ST_fsm_state9;
        end
        ap_ST_fsm_state9 : begin
            ap_NS_fsm = ap_ST_fsm_state10;
        end
        ap_ST_fsm_state10 : begin
            ap_NS_fsm = ap_ST_fsm_state11;
        end
        ap_ST_fsm_state11 : begin
            ap_NS_fsm = ap_ST_fsm_state12;
        end
        ap_ST_fsm_state12 : begin
            ap_NS_fsm = ap_ST_fsm_state13;
        end
        ap_ST_fsm_state13 : begin
            ap_NS_fsm = ap_ST_fsm_state14;
        end
        ap_ST_fsm_state14 : begin
            ap_NS_fsm = ap_ST_fsm_state15;
        end
        ap_ST_fsm_state15 : begin
            ap_NS_fsm = ap_ST_fsm_state16;
        end
        ap_ST_fsm_state16 : begin
            ap_NS_fsm = ap_ST_fsm_state17;
        end
        ap_ST_fsm_state17 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign adjustments_address0 = zext_ln220_fu_90_p1;

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state12 = ap_CS_fsm[32'd11];

assign ap_CS_fsm_state13 = ap_CS_fsm[32'd12];

assign ap_CS_fsm_state17 = ap_CS_fsm[32'd16];

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

assign ap_CS_fsm_state8 = ap_CS_fsm[32'd7];

assign ap_CS_fsm_state9 = ap_CS_fsm[32'd8];

always @ (*) begin
    ap_block_state1 = ((input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0));
end

assign ap_return = ((tmp_fu_136_p3[0:0] == 1'b1) ? 16'd0 : grp_fu_77_p2);

assign bitcast_ln648_fu_132_p1 = grp_fu_77_p2;

assign grp_fu_77_p1 = tmp_16_i_i_reg_172;

assign grp_fu_81_p1 = trunc_ln220_fu_95_p1;

assign grp_fu_86_p1 = tmp_15_i_i_reg_167;

assign tmp_fu_136_p3 = bitcast_ln648_fu_132_p1[32'd15];

assign trunc_ln220_fu_95_p1 = adjustments_q0[15:0];

assign zext_ln220_fu_90_p1 = input_indices_23_dout;

endmodule //td_fused_top_tdf8_adjust
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf8_dot_product (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        ifmap_vec_address0,
        ifmap_vec_ce0,
        ifmap_vec_q0,
        weight_vecs_0_address0,
        weight_vecs_0_ce0,
        weight_vecs_0_q0,
        products_0_address0,
        products_0_ce0,
        products_0_we0,
        products_0_d0
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state10 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [8:0] ifmap_vec_address0;
output   ifmap_vec_ce0;
input  [15:0] ifmap_vec_q0;
output  [8:0] weight_vecs_0_address0;
output   weight_vecs_0_ce0;
input  [15:0] weight_vecs_0_q0;
output  [8:0] products_0_address0;
output   products_0_ce0;
output   products_0_we0;
output  [15:0] products_0_d0;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg ifmap_vec_ce0;
reg weight_vecs_0_ce0;
reg products_0_ce0;
reg products_0_we0;

reg    ap_done_reg;
  reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg   [8:0] indvar_flatten17_reg_97;
reg   [7:0] indvar_flatten_reg_108;
reg   [1:0] jj_reg_119;
reg   [5:0] ic_reg_131;
reg   [1:0] ii_reg_142;
wire   [8:0] add_ln147_1_fu_157_p2;
wire    ap_CS_fsm_pp0_stage0;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
wire    ap_block_state4_pp0_stage0_iter2;
wire    ap_block_state5_pp0_stage0_iter3;
wire    ap_block_state6_pp0_stage0_iter4;
wire    ap_block_state7_pp0_stage0_iter5;
wire    ap_block_state8_pp0_stage0_iter6;
wire    ap_block_state9_pp0_stage0_iter7;
wire    ap_block_pp0_stage0_11001;
wire   [0:0] icmp_ln147_fu_163_p2;
reg   [0:0] icmp_ln147_reg_408;
reg   [0:0] icmp_ln147_reg_408_pp0_iter1_reg;
reg   [0:0] icmp_ln147_reg_408_pp0_iter2_reg;
reg   [0:0] icmp_ln147_reg_408_pp0_iter3_reg;
reg   [0:0] icmp_ln147_reg_408_pp0_iter4_reg;
reg   [0:0] icmp_ln147_reg_408_pp0_iter5_reg;
reg   [0:0] icmp_ln147_reg_408_pp0_iter6_reg;
wire   [0:0] icmp_ln148_fu_169_p2;
reg   [0:0] icmp_ln148_reg_412;
wire   [0:0] and_ln147_fu_195_p2;
reg   [0:0] and_ln147_reg_419;
wire   [1:0] add_ln148_fu_201_p2;
reg   [1:0] add_ln148_reg_424;
wire   [5:0] select_ln148_fu_213_p3;
reg   [5:0] select_ln148_reg_429;
wire   [1:0] select_ln148_1_fu_221_p3;
reg   [1:0] select_ln148_1_reg_434;
wire   [4:0] trunc_ln150_fu_229_p1;
reg   [4:0] trunc_ln150_reg_440;
reg   [4:0] trunc_ln150_reg_440_pp0_iter1_reg;
reg   [4:0] trunc_ln150_reg_440_pp0_iter2_reg;
reg   [4:0] trunc_ln150_reg_440_pp0_iter3_reg;
reg   [4:0] trunc_ln150_reg_440_pp0_iter4_reg;
reg   [4:0] trunc_ln150_reg_440_pp0_iter5_reg;
reg   [4:0] trunc_ln150_reg_440_pp0_iter6_reg;
wire   [5:0] add_ln149_fu_233_p2;
wire   [7:0] select_ln148_3_fu_245_p3;
wire   [1:0] select_ln147_2_fu_287_p3;
reg   [1:0] select_ln147_2_reg_455;
reg    ap_enable_reg_pp0_iter1;
wire   [3:0] select_ln148_2_fu_370_p3;
reg   [3:0] select_ln148_2_reg_460;
reg   [3:0] select_ln148_2_reg_460_pp0_iter2_reg;
reg   [3:0] select_ln148_2_reg_460_pp0_iter3_reg;
reg   [3:0] select_ln148_2_reg_460_pp0_iter4_reg;
reg   [3:0] select_ln148_2_reg_460_pp0_iter5_reg;
reg   [3:0] select_ln148_2_reg_460_pp0_iter6_reg;
reg   [15:0] ifmap_vec_load_reg_475;
reg   [15:0] weight_vecs_0_load_reg_480;
wire   [15:0] grp_fu_153_p2;
reg   [15:0] mul_reg_485;
reg    ap_block_state1;
wire    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_flush_enable;
reg    ap_enable_reg_pp0_iter2;
reg    ap_condition_pp0_exit_iter1_state3;
reg    ap_enable_reg_pp0_iter3;
reg    ap_enable_reg_pp0_iter4;
reg    ap_enable_reg_pp0_iter5;
reg    ap_enable_reg_pp0_iter6;
reg    ap_enable_reg_pp0_iter7;
reg   [1:0] ap_phi_mux_jj_phi_fu_123_p4;
wire    ap_block_pp0_stage0;
reg   [1:0] ap_phi_mux_ii_phi_fu_146_p4;
wire   [63:0] p_cast25_fu_386_p1;
wire   [63:0] idxprom30_fu_398_p1;
wire   [0:0] icmp_ln149_fu_189_p2;
wire   [0:0] xor_ln147_fu_183_p2;
wire   [1:0] select_ln147_fu_175_p3;
wire   [0:0] or_ln148_fu_207_p2;
wire   [7:0] add_ln148_1_fu_239_p2;
wire   [3:0] shl_ln_fu_257_p3;
wire   [3:0] zext_ln150_fu_253_p1;
wire   [3:0] sub_ln150_fu_265_p2;
wire   [3:0] zext_ln150_1_fu_271_p1;
wire   [1:0] add_ln147_fu_281_p2;
wire   [3:0] tmp_fu_298_p3;
wire   [3:0] select_ln147_2_cast_fu_294_p1;
wire   [3:0] shl_ln150_mid1_fu_316_p3;
wire   [3:0] zext_ln150_2_fu_312_p1;
wire   [3:0] sub_ln150_1_fu_324_p2;
wire   [3:0] add_ln150_fu_275_p2;
wire   [3:0] empty_64_fu_306_p2;
wire   [3:0] select_ln148_1_cast_fu_344_p1;
wire   [3:0] empty_65_fu_347_p2;
wire   [3:0] select_ln147_3_fu_330_p3;
wire   [3:0] zext_ln150_3_fu_361_p1;
wire   [3:0] add_ln150_1_fu_364_p2;
wire   [3:0] select_ln147_4_fu_337_p3;
wire   [8:0] tmp_28_cast_fu_353_p3;
wire   [8:0] select_ln148_cast_fu_377_p1;
wire   [8:0] empty_66_fu_380_p2;
wire   [8:0] p_fu_392_p3;
wire    ap_CS_fsm_state10;
reg   [2:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
#0 ap_enable_reg_pp0_iter4 = 1'b0;
#0 ap_enable_reg_pp0_iter5 = 1'b0;
#0 ap_enable_reg_pp0_iter6 = 1'b0;
#0 ap_enable_reg_pp0_iter7 = 1'b0;
end

td_fused_top_hmul_16ns_16ns_16_4_max_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hmul_16ns_16ns_16_4_max_dsp_1_U494(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(ifmap_vec_load_reg_475),
    .din1(weight_vecs_0_load_reg_480),
    .dout(grp_fu_153_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state10)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if ((1'b1 == ap_condition_pp0_flush_enable)) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            if ((1'b1 == ap_condition_pp0_exit_iter1_state3)) begin
                ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter0;
            end else if ((1'b1 == 1'b1)) begin
                ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
            end
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter4 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter5 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter5 <= ap_enable_reg_pp0_iter4;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter6 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter6 <= ap_enable_reg_pp0_iter5;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter7 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter7 <= ap_enable_reg_pp0_iter6;
        end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter7 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_fu_163_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ic_reg_131 <= add_ln149_fu_233_p2;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ic_reg_131 <= 6'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_reg_408_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        ii_reg_142 <= select_ln147_2_reg_455;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ii_reg_142 <= 2'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_fu_163_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        indvar_flatten17_reg_97 <= add_ln147_1_fu_157_p2;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indvar_flatten17_reg_97 <= 9'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_fu_163_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        indvar_flatten_reg_108 <= select_ln148_3_fu_245_p3;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indvar_flatten_reg_108 <= 8'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_reg_408 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        jj_reg_119 <= select_ln148_1_reg_434;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        jj_reg_119 <= 2'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_fu_163_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        add_ln148_reg_424 <= add_ln148_fu_201_p2;
        and_ln147_reg_419 <= and_ln147_fu_195_p2;
        icmp_ln148_reg_412 <= icmp_ln148_fu_169_p2;
        select_ln148_reg_429 <= select_ln148_fu_213_p3;
        trunc_ln150_reg_440 <= trunc_ln150_fu_229_p1;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln147_reg_408 <= icmp_ln147_fu_163_p2;
        icmp_ln147_reg_408_pp0_iter1_reg <= icmp_ln147_reg_408;
        trunc_ln150_reg_440_pp0_iter1_reg <= trunc_ln150_reg_440;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        icmp_ln147_reg_408_pp0_iter2_reg <= icmp_ln147_reg_408_pp0_iter1_reg;
        icmp_ln147_reg_408_pp0_iter3_reg <= icmp_ln147_reg_408_pp0_iter2_reg;
        icmp_ln147_reg_408_pp0_iter4_reg <= icmp_ln147_reg_408_pp0_iter3_reg;
        icmp_ln147_reg_408_pp0_iter5_reg <= icmp_ln147_reg_408_pp0_iter4_reg;
        icmp_ln147_reg_408_pp0_iter6_reg <= icmp_ln147_reg_408_pp0_iter5_reg;
        select_ln148_2_reg_460_pp0_iter2_reg <= select_ln148_2_reg_460;
        select_ln148_2_reg_460_pp0_iter3_reg <= select_ln148_2_reg_460_pp0_iter2_reg;
        select_ln148_2_reg_460_pp0_iter4_reg <= select_ln148_2_reg_460_pp0_iter3_reg;
        select_ln148_2_reg_460_pp0_iter5_reg <= select_ln148_2_reg_460_pp0_iter4_reg;
        select_ln148_2_reg_460_pp0_iter6_reg <= select_ln148_2_reg_460_pp0_iter5_reg;
        trunc_ln150_reg_440_pp0_iter2_reg <= trunc_ln150_reg_440_pp0_iter1_reg;
        trunc_ln150_reg_440_pp0_iter3_reg <= trunc_ln150_reg_440_pp0_iter2_reg;
        trunc_ln150_reg_440_pp0_iter4_reg <= trunc_ln150_reg_440_pp0_iter3_reg;
        trunc_ln150_reg_440_pp0_iter5_reg <= trunc_ln150_reg_440_pp0_iter4_reg;
        trunc_ln150_reg_440_pp0_iter6_reg <= trunc_ln150_reg_440_pp0_iter5_reg;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_reg_408_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        ifmap_vec_load_reg_475 <= ifmap_vec_q0;
        weight_vecs_0_load_reg_480 <= weight_vecs_0_q0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_reg_408_pp0_iter5_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        mul_reg_485 <= grp_fu_153_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_reg_408 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        select_ln147_2_reg_455 <= select_ln147_2_fu_287_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_fu_163_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        select_ln148_1_reg_434 <= select_ln148_1_fu_221_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln147_reg_408 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        select_ln148_2_reg_460 <= select_ln148_2_fu_370_p3;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_condition_pp0_exit_iter1_state3 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter1_state3 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln147_fu_163_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_condition_pp0_flush_enable = 1'b1;
    end else begin
        ap_condition_pp0_flush_enable = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state10)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter7 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln147_reg_408_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        ap_phi_mux_ii_phi_fu_146_p4 = select_ln147_2_reg_455;
    end else begin
        ap_phi_mux_ii_phi_fu_146_p4 = ii_reg_142;
    end
end

always @ (*) begin
    if (((icmp_ln147_reg_408 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_jj_phi_fu_123_p4 = select_ln148_1_reg_434;
    end else begin
        ap_phi_mux_jj_phi_fu_123_p4 = jj_reg_119;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state10)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ifmap_vec_ce0 = 1'b1;
    end else begin
        ifmap_vec_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter7 == 1'b1))) begin
        products_0_ce0 = 1'b1;
    end else begin
        products_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln147_reg_408_pp0_iter6_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter7 == 1'b1))) begin
        products_0_we0 = 1'b1;
    end else begin
        products_0_we0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        weight_vecs_0_ce0 = 1'b1;
    end else begin
        weight_vecs_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((~((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b1)) & ~((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter7 == 1'b1) & (ap_enable_reg_pp0_iter6 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if ((((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter7 == 1'b1) & (ap_enable_reg_pp0_iter6 == 1'b0)) | ((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b1)))) begin
                ap_NS_fsm = ap_ST_fsm_state10;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state10 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln147_1_fu_157_p2 = (indvar_flatten17_reg_97 + 9'd1);

assign add_ln147_fu_281_p2 = (ap_phi_mux_ii_phi_fu_146_p4 + 2'd1);

assign add_ln148_1_fu_239_p2 = (indvar_flatten_reg_108 + 8'd1);

assign add_ln148_fu_201_p2 = (select_ln147_fu_175_p3 + 2'd1);

assign add_ln149_fu_233_p2 = (select_ln148_fu_213_p3 + 6'd1);

assign add_ln150_1_fu_364_p2 = (select_ln147_3_fu_330_p3 + zext_ln150_3_fu_361_p1);

assign add_ln150_fu_275_p2 = (sub_ln150_fu_265_p2 + zext_ln150_1_fu_271_p1);

assign and_ln147_fu_195_p2 = (xor_ln147_fu_183_p2 & icmp_ln149_fu_189_p2);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state10 = ap_CS_fsm[32'd2];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (ap_done_reg == 1'b1));
end

assign ap_block_state2_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter4 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage0_iter5 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage0_iter6 = ~(1'b1 == 1'b1);

assign ap_block_state9_pp0_stage0_iter7 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign empty_64_fu_306_p2 = (tmp_fu_298_p3 - select_ln147_2_cast_fu_294_p1);

assign empty_65_fu_347_p2 = (empty_64_fu_306_p2 + select_ln148_1_cast_fu_344_p1);

assign empty_66_fu_380_p2 = (tmp_28_cast_fu_353_p3 + select_ln148_cast_fu_377_p1);

assign icmp_ln147_fu_163_p2 = ((indvar_flatten17_reg_97 == 9'd288) ? 1'b1 : 1'b0);

assign icmp_ln148_fu_169_p2 = ((indvar_flatten_reg_108 == 8'd96) ? 1'b1 : 1'b0);

assign icmp_ln149_fu_189_p2 = ((ic_reg_131 == 6'd32) ? 1'b1 : 1'b0);

assign idxprom30_fu_398_p1 = p_fu_392_p3;

assign ifmap_vec_address0 = p_cast25_fu_386_p1;

assign or_ln148_fu_207_p2 = (icmp_ln148_fu_169_p2 | and_ln147_fu_195_p2);

assign p_cast25_fu_386_p1 = empty_66_fu_380_p2;

assign p_fu_392_p3 = {{select_ln148_2_reg_460_pp0_iter6_reg}, {trunc_ln150_reg_440_pp0_iter6_reg}};

assign products_0_address0 = idxprom30_fu_398_p1;

assign products_0_d0 = mul_reg_485;

assign select_ln147_2_cast_fu_294_p1 = select_ln147_2_fu_287_p3;

assign select_ln147_2_fu_287_p3 = ((icmp_ln148_reg_412[0:0] == 1'b1) ? add_ln147_fu_281_p2 : ap_phi_mux_ii_phi_fu_146_p4);

assign select_ln147_3_fu_330_p3 = ((icmp_ln148_reg_412[0:0] == 1'b1) ? sub_ln150_1_fu_324_p2 : sub_ln150_fu_265_p2);

assign select_ln147_4_fu_337_p3 = ((icmp_ln148_reg_412[0:0] == 1'b1) ? sub_ln150_1_fu_324_p2 : add_ln150_fu_275_p2);

assign select_ln147_fu_175_p3 = ((icmp_ln148_fu_169_p2[0:0] == 1'b1) ? 2'd0 : ap_phi_mux_jj_phi_fu_123_p4);

assign select_ln148_1_cast_fu_344_p1 = select_ln148_1_reg_434;

assign select_ln148_1_fu_221_p3 = ((and_ln147_fu_195_p2[0:0] == 1'b1) ? add_ln148_fu_201_p2 : select_ln147_fu_175_p3);

assign select_ln148_2_fu_370_p3 = ((and_ln147_reg_419[0:0] == 1'b1) ? add_ln150_1_fu_364_p2 : select_ln147_4_fu_337_p3);

assign select_ln148_3_fu_245_p3 = ((icmp_ln148_fu_169_p2[0:0] == 1'b1) ? 8'd1 : add_ln148_1_fu_239_p2);

assign select_ln148_cast_fu_377_p1 = select_ln148_reg_429;

assign select_ln148_fu_213_p3 = ((or_ln148_fu_207_p2[0:0] == 1'b1) ? 6'd0 : ic_reg_131);

assign shl_ln150_mid1_fu_316_p3 = {{add_ln147_fu_281_p2}, {2'd0}};

assign shl_ln_fu_257_p3 = {{ap_phi_mux_ii_phi_fu_146_p4}, {2'd0}};

assign sub_ln150_1_fu_324_p2 = (shl_ln150_mid1_fu_316_p3 - zext_ln150_2_fu_312_p1);

assign sub_ln150_fu_265_p2 = (shl_ln_fu_257_p3 - zext_ln150_fu_253_p1);

assign tmp_28_cast_fu_353_p3 = {{empty_65_fu_347_p2}, {5'd0}};

assign tmp_fu_298_p3 = {{select_ln147_2_fu_287_p3}, {2'd0}};

assign trunc_ln150_fu_229_p1 = select_ln148_fu_213_p3[4:0];

assign weight_vecs_0_address0 = p_cast25_fu_386_p1;

assign xor_ln147_fu_183_p2 = (icmp_ln148_fu_169_p2 ^ 1'd1);

assign zext_ln150_1_fu_271_p1 = jj_reg_119;

assign zext_ln150_2_fu_312_p1 = add_ln147_fu_281_p2;

assign zext_ln150_3_fu_361_p1 = add_ln148_reg_424;

assign zext_ln150_fu_253_p1 = ap_phi_mux_ii_phi_fu_146_p4;

endmodule //td_fused_top_tdf8_dot_product
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf8_get_next_ijk (
        ap_clk,
        ap_rst,
        ap_start,
        start_full_n,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        start_out,
        start_write,
        input_indices_2_out_din,
        input_indices_2_out_full_n,
        input_indices_2_out_write,
        input_indices_2_out1_din,
        input_indices_2_out1_full_n,
        input_indices_2_out1_write,
        output_indices_0_din,
        output_indices_0_full_n,
        output_indices_0_write,
        output_indices_1_din,
        output_indices_1_full_n,
        output_indices_1_write,
        resetMaximum_din,
        resetMaximum_full_n,
        resetMaximum_write,
        storeOutput_din,
        storeOutput_full_n,
        storeOutput_write,
        ap_return_0,
        ap_return_1
);

parameter    ap_ST_fsm_state1 = 1'd1;

input   ap_clk;
input   ap_rst;
input   ap_start;
input   start_full_n;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output   start_out;
output   start_write;
output  [7:0] input_indices_2_out_din;
input   input_indices_2_out_full_n;
output   input_indices_2_out_write;
output  [7:0] input_indices_2_out1_din;
input   input_indices_2_out1_full_n;
output   input_indices_2_out1_write;
output  [3:0] output_indices_0_din;
input   output_indices_0_full_n;
output   output_indices_0_write;
output  [7:0] output_indices_1_din;
input   output_indices_1_full_n;
output   output_indices_1_write;
output   resetMaximum_din;
input   resetMaximum_full_n;
output   resetMaximum_write;
output   storeOutput_din;
input   storeOutput_full_n;
output   storeOutput_write;
output  [15:0] ap_return_0;
output  [15:0] ap_return_1;

reg ap_done;
reg ap_idle;
reg start_write;
reg input_indices_2_out_write;
reg input_indices_2_out1_write;
reg output_indices_0_write;
reg output_indices_1_write;
reg resetMaximum_write;
reg storeOutput_write;

reg    real_start;
reg    start_once_reg;
reg    ap_done_reg;
  reg   [0:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    internal_ap_ready;
reg   [1:0] i_p;
reg   [1:0] j_p;
reg   [15:0] i_8;
reg   [15:0] j_8;
reg   [15:0] k_8;
reg   [15:0] i_out;
reg   [15:0] j_out;
reg    input_indices_2_out_blk_n;
reg    input_indices_2_out1_blk_n;
reg    output_indices_0_blk_n;
reg    output_indices_1_blk_n;
reg    resetMaximum_blk_n;
reg    storeOutput_blk_n;
wire   [1:0] select_ln142_fu_336_p3;
reg    ap_block_state1;
wire   [0:0] or_ln142_fu_310_p2;
wire   [1:0] select_ln142_1_fu_344_p3;
wire   [15:0] select_ln147_fu_276_p3;
wire   [0:0] and_ln142_1_fu_304_p2;
wire   [15:0] select_ln142_2_fu_358_p3;
wire   [0:0] and_ln132_fu_352_p2;
wire   [15:0] select_ln142_3_fu_386_p3;
wire   [0:0] and_ln135_fu_292_p2;
wire   [15:0] select_ln147_1_fu_284_p3;
wire   [15:0] select_ln142_4_fu_394_p3;
wire   [7:0] trunc_ln128_fu_180_p1;
wire   [1:0] or_ln124_fu_124_p2;
wire   [0:0] icmp_ln125_fu_137_p2;
wire   [0:0] icmp_ln125_1_fu_143_p2;
wire   [15:0] zext_ln126_fu_112_p1;
wire   [15:0] zext_ln127_fu_120_p1;
wire   [1:0] add_ln131_fu_204_p2;
wire   [1:0] add_ln134_fu_216_p2;
wire   [15:0] add_ln137_fu_228_p2;
wire   [15:0] add_ln141_fu_246_p2;
wire   [15:0] add_ln146_fu_264_p2;
wire   [0:0] icmp_ln147_fu_270_p2;
wire   [15:0] add_ln145_fu_258_p2;
wire   [0:0] icmp_ln132_fu_210_p2;
wire   [0:0] icmp_ln135_fu_222_p2;
wire   [0:0] icmp_ln138_fu_234_p2;
wire   [0:0] icmp_ln142_fu_252_p2;
wire   [0:0] and_ln142_fu_298_p2;
wire   [0:0] xor_ln135_fu_316_p2;
wire   [0:0] and_ln135_1_fu_322_p2;
wire   [1:0] select_ln135_fu_328_p3;
wire   [15:0] add_ln140_fu_240_p2;
wire   [0:0] xor_ln138_fu_366_p2;
wire   [0:0] and_ln138_fu_372_p2;
wire   [15:0] select_ln138_fu_378_p3;
wire   [15:0] add_ln126_fu_160_p2;
wire   [15:0] add_ln127_fu_170_p2;
reg   [0:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 start_once_reg = 1'b0;
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 1'd1;
#0 i_p = 2'd0;
#0 j_p = 2'd0;
#0 i_8 = 16'd0;
#0 j_8 = 16'd0;
#0 k_8 = 16'd0;
#0 i_out = 16'd0;
#0 j_out = 16'd0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        start_once_reg <= 1'b0;
    end else begin
        if (((real_start == 1'b1) & (internal_ap_ready == 1'b0))) begin
            start_once_reg <= 1'b1;
        end else if ((internal_ap_ready == 1'b1)) begin
            start_once_reg <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1) & (1'd1 == and_ln142_1_fu_304_p2))) begin
        i_8 <= select_ln147_fu_276_p3;
        i_out <= select_ln147_1_fu_284_p3;
    end
end

always @ (posedge ap_clk) begin
    if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (or_ln142_fu_310_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1))) begin
        i_p <= select_ln142_fu_336_p3;
    end
end

always @ (posedge ap_clk) begin
    if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1) & (1'd1 == and_ln132_fu_352_p2))) begin
        j_8 <= select_ln142_2_fu_358_p3;
        j_out <= select_ln142_4_fu_394_p3;
    end
end

always @ (posedge ap_clk) begin
    if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        j_p <= select_ln142_1_fu_344_p3;
    end
end

always @ (posedge ap_clk) begin
    if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1) & (1'd1 == and_ln135_fu_292_p2))) begin
        k_8 <= select_ln142_3_fu_386_p3;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((real_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        input_indices_2_out1_blk_n = input_indices_2_out1_full_n;
    end else begin
        input_indices_2_out1_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        input_indices_2_out1_write = 1'b1;
    end else begin
        input_indices_2_out1_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        input_indices_2_out_blk_n = input_indices_2_out_full_n;
    end else begin
        input_indices_2_out_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        input_indices_2_out_write = 1'b1;
    end else begin
        input_indices_2_out_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        internal_ap_ready = 1'b1;
    end else begin
        internal_ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        output_indices_0_blk_n = output_indices_0_full_n;
    end else begin
        output_indices_0_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        output_indices_0_write = 1'b1;
    end else begin
        output_indices_0_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        output_indices_1_blk_n = output_indices_1_full_n;
    end else begin
        output_indices_1_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        output_indices_1_write = 1'b1;
    end else begin
        output_indices_1_write = 1'b0;
    end
end

always @ (*) begin
    if (((start_full_n == 1'b0) & (start_once_reg == 1'b0))) begin
        real_start = 1'b0;
    end else begin
        real_start = ap_start;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        resetMaximum_blk_n = resetMaximum_full_n;
    end else begin
        resetMaximum_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        resetMaximum_write = 1'b1;
    end else begin
        resetMaximum_write = 1'b0;
    end
end

always @ (*) begin
    if (((real_start == 1'b1) & (start_once_reg == 1'b0))) begin
        start_write = 1'b1;
    end else begin
        start_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        storeOutput_blk_n = storeOutput_full_n;
    end else begin
        storeOutput_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        storeOutput_write = 1'b1;
    end else begin
        storeOutput_write = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln126_fu_160_p2 = (i_8 + zext_ln126_fu_112_p1);

assign add_ln127_fu_170_p2 = (j_8 + zext_ln127_fu_120_p1);

assign add_ln131_fu_204_p2 = (j_p + 2'd1);

assign add_ln134_fu_216_p2 = (i_p + 2'd1);

assign add_ln137_fu_228_p2 = (k_8 + 16'd1);

assign add_ln140_fu_240_p2 = (j_8 + 16'd2);

assign add_ln141_fu_246_p2 = (j_out + 16'd1);

assign add_ln145_fu_258_p2 = (i_8 + 16'd2);

assign add_ln146_fu_264_p2 = (i_out + 16'd1);

assign and_ln132_fu_352_p2 = (icmp_ln138_fu_234_p2 & and_ln135_fu_292_p2);

assign and_ln135_1_fu_322_p2 = (xor_ln135_fu_316_p2 & icmp_ln132_fu_210_p2);

assign and_ln135_fu_292_p2 = (icmp_ln135_fu_222_p2 & icmp_ln132_fu_210_p2);

assign and_ln138_fu_372_p2 = (xor_ln138_fu_366_p2 & and_ln135_fu_292_p2);

assign and_ln142_1_fu_304_p2 = (and_ln142_fu_298_p2 & and_ln135_fu_292_p2);

assign and_ln142_fu_298_p2 = (icmp_ln142_fu_252_p2 & icmp_ln138_fu_234_p2);

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

always @ (*) begin
    ap_block_state1 = ((real_start == 1'b0) | (storeOutput_full_n == 1'b0) | (resetMaximum_full_n == 1'b0) | (output_indices_1_full_n == 1'b0) | (output_indices_0_full_n == 1'b0) | (input_indices_2_out1_full_n == 1'b0) | (input_indices_2_out_full_n == 1'b0) | (ap_done_reg == 1'b1));
end

assign ap_ready = internal_ap_ready;

assign ap_return_0 = add_ln126_fu_160_p2;

assign ap_return_1 = add_ln127_fu_170_p2;

assign icmp_ln125_1_fu_143_p2 = ((j_p == 2'd1) ? 1'b1 : 1'b0);

assign icmp_ln125_fu_137_p2 = ((i_p == 2'd1) ? 1'b1 : 1'b0);

assign icmp_ln132_fu_210_p2 = ((add_ln131_fu_204_p2 == 2'd2) ? 1'b1 : 1'b0);

assign icmp_ln135_fu_222_p2 = ((add_ln134_fu_216_p2 == 2'd2) ? 1'b1 : 1'b0);

assign icmp_ln138_fu_234_p2 = ((add_ln137_fu_228_p2 == 16'd256) ? 1'b1 : 1'b0);

assign icmp_ln142_fu_252_p2 = ((add_ln141_fu_246_p2 == 16'd14) ? 1'b1 : 1'b0);

assign icmp_ln147_fu_270_p2 = ((add_ln146_fu_264_p2 == 16'd14) ? 1'b1 : 1'b0);

assign input_indices_2_out1_din = trunc_ln128_fu_180_p1;

assign input_indices_2_out_din = trunc_ln128_fu_180_p1;

assign or_ln124_fu_124_p2 = (j_p | i_p);

assign or_ln142_fu_310_p2 = (icmp_ln132_fu_210_p2 | and_ln142_1_fu_304_p2);

assign output_indices_0_din = i_out[3:0];

assign output_indices_1_din = j_out[7:0];

assign resetMaximum_din = ((or_ln124_fu_124_p2 == 2'd0) ? 1'b1 : 1'b0);

assign select_ln135_fu_328_p3 = ((and_ln135_1_fu_322_p2[0:0] == 1'b1) ? add_ln134_fu_216_p2 : 2'd0);

assign select_ln138_fu_378_p3 = ((and_ln138_fu_372_p2[0:0] == 1'b1) ? add_ln137_fu_228_p2 : 16'd0);

assign select_ln142_1_fu_344_p3 = ((or_ln142_fu_310_p2[0:0] == 1'b1) ? 2'd0 : add_ln131_fu_204_p2);

assign select_ln142_2_fu_358_p3 = ((and_ln142_1_fu_304_p2[0:0] == 1'b1) ? 16'd0 : add_ln140_fu_240_p2);

assign select_ln142_3_fu_386_p3 = ((and_ln142_1_fu_304_p2[0:0] == 1'b1) ? 16'd0 : select_ln138_fu_378_p3);

assign select_ln142_4_fu_394_p3 = ((and_ln142_1_fu_304_p2[0:0] == 1'b1) ? 16'd0 : add_ln141_fu_246_p2);

assign select_ln142_fu_336_p3 = ((and_ln142_1_fu_304_p2[0:0] == 1'b1) ? 2'd0 : select_ln135_fu_328_p3);

assign select_ln147_1_fu_284_p3 = ((icmp_ln147_fu_270_p2[0:0] == 1'b1) ? 16'd0 : add_ln146_fu_264_p2);

assign select_ln147_fu_276_p3 = ((icmp_ln147_fu_270_p2[0:0] == 1'b1) ? 16'd0 : add_ln145_fu_258_p2);

assign start_out = real_start;

assign storeOutput_din = (icmp_ln125_fu_137_p2 & icmp_ln125_1_fu_143_p2);

assign trunc_ln128_fu_180_p1 = k_8[7:0];

assign xor_ln135_fu_316_p2 = (icmp_ln135_fu_222_p2 ^ 1'd1);

assign xor_ln138_fu_366_p2 = (icmp_ln138_fu_234_p2 ^ 1'd1);

assign zext_ln126_fu_112_p1 = i_p;

assign zext_ln127_fu_120_p1 = j_p;

endmodule //td_fused_top_tdf8_get_next_ijk
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf8_poolOutputs (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        output_indices_04_dout,
        output_indices_04_empty_n,
        output_indices_04_read,
        output_indices_15_dout,
        output_indices_15_empty_n,
        output_indices_15_read,
        resetMaximum6_dout,
        resetMaximum6_empty_n,
        resetMaximum6_read,
        storeOutput7_dout,
        storeOutput7_empty_n,
        storeOutput7_read,
        p_read,
        out_data_address1,
        out_data_ce1,
        out_data_we1,
        out_data_d1
);

parameter    ap_ST_fsm_state1 = 4'd1;
parameter    ap_ST_fsm_state2 = 4'd2;
parameter    ap_ST_fsm_state3 = 4'd4;
parameter    ap_ST_fsm_state4 = 4'd8;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
input  [3:0] output_indices_04_dout;
input   output_indices_04_empty_n;
output   output_indices_04_read;
input  [7:0] output_indices_15_dout;
input   output_indices_15_empty_n;
output   output_indices_15_read;
input  [0:0] resetMaximum6_dout;
input   resetMaximum6_empty_n;
output   resetMaximum6_read;
input  [0:0] storeOutput7_dout;
input   storeOutput7_empty_n;
output   storeOutput7_read;
input  [15:0] p_read;
output  [13:0] out_data_address1;
output   out_data_ce1;
output   out_data_we1;
output  [63:0] out_data_d1;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg output_indices_04_read;
reg output_indices_15_read;
reg resetMaximum6_read;
reg storeOutput7_read;

reg    ap_done_reg;
  reg   [3:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg   [15:0] max_vals_0;
reg    output_indices_04_blk_n;
wire    ap_CS_fsm_state2;
reg    output_indices_15_blk_n;
reg    resetMaximum6_blk_n;
reg    storeOutput7_blk_n;
reg   [3:0] output_indices_04_read_reg_147;
reg   [7:0] output_indices_15_read_reg_152;
wire   [0:0] storeOutput7_read_read_fu_82_p2;
reg   [0:0] storeOutput7_read_reg_157;
wire    grp_tdf8_writeOutputs_unaligned_fu_88_ap_start;
wire    grp_tdf8_writeOutputs_unaligned_fu_88_ap_done;
wire    grp_tdf8_writeOutputs_unaligned_fu_88_ap_idle;
wire    grp_tdf8_writeOutputs_unaligned_fu_88_ap_ready;
wire   [13:0] grp_tdf8_writeOutputs_unaligned_fu_88_out_data_address1;
wire    grp_tdf8_writeOutputs_unaligned_fu_88_out_data_ce1;
wire    grp_tdf8_writeOutputs_unaligned_fu_88_out_data_we1;
wire   [63:0] grp_tdf8_writeOutputs_unaligned_fu_88_out_data_d1;
reg    grp_tdf8_writeOutputs_unaligned_fu_88_ap_start_reg;
wire    ap_CS_fsm_state3;
wire    ap_CS_fsm_state4;
reg    ap_block_state4_on_subcall_done;
wire   [15:0] select_ln24_fu_126_p3;
reg    ap_block_state2;
reg    ap_block_state1;
wire   [0:0] grp_fu_110_p2;
wire   [0:0] or_ln24_fu_120_p2;
reg    grp_fu_110_ce;
reg   [3:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 4'd1;
#0 max_vals_0 = 16'd0;
#0 grp_tdf8_writeOutputs_unaligned_fu_88_ap_start_reg = 1'b0;
end

td_fused_top_tdf8_writeOutputs_unaligned grp_tdf8_writeOutputs_unaligned_fu_88(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(grp_tdf8_writeOutputs_unaligned_fu_88_ap_start),
    .ap_done(grp_tdf8_writeOutputs_unaligned_fu_88_ap_done),
    .ap_idle(grp_tdf8_writeOutputs_unaligned_fu_88_ap_idle),
    .ap_ready(grp_tdf8_writeOutputs_unaligned_fu_88_ap_ready),
    .i(output_indices_04_read_reg_147),
    .j(output_indices_15_read_reg_152),
    .out_data_address1(grp_tdf8_writeOutputs_unaligned_fu_88_out_data_address1),
    .out_data_ce1(grp_tdf8_writeOutputs_unaligned_fu_88_out_data_ce1),
    .out_data_we1(grp_tdf8_writeOutputs_unaligned_fu_88_out_data_we1),
    .out_data_d1(grp_tdf8_writeOutputs_unaligned_fu_88_out_data_d1),
    .max_vals_0(max_vals_0)
);

td_fused_top_hcmp_16ns_16ns_1_2_no_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 2 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 1 ))
hcmp_16ns_16ns_1_2_no_dsp_1_U516(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(grp_fu_110_ce),
    .din0(max_vals_0),
    .din1(p_read),
    .opcode(5'd4),
    .dout(grp_fu_110_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_state4) & (1'b0 == ap_block_state4_on_subcall_done))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        grp_tdf8_writeOutputs_unaligned_fu_88_ap_start_reg <= 1'b0;
    end else begin
        if ((1'b1 == ap_CS_fsm_state3)) begin
            grp_tdf8_writeOutputs_unaligned_fu_88_ap_start_reg <= 1'b1;
        end else if ((grp_tdf8_writeOutputs_unaligned_fu_88_ap_ready == 1'b1)) begin
            grp_tdf8_writeOutputs_unaligned_fu_88_ap_start_reg <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((~((storeOutput7_empty_n == 1'b0) | (resetMaximum6_empty_n == 1'b0) | (output_indices_15_empty_n == 1'b0) | (output_indices_04_empty_n == 1'b0)) & (1'b1 == ap_CS_fsm_state2))) begin
        max_vals_0 <= select_ln24_fu_126_p3;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        output_indices_04_read_reg_147 <= output_indices_04_dout;
        output_indices_15_read_reg_152 <= output_indices_15_dout;
        storeOutput7_read_reg_157 <= storeOutput7_dout;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state4) & (1'b0 == ap_block_state4_on_subcall_done))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state4) & (1'b0 == ap_block_state4_on_subcall_done))) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1)) | (~((storeOutput7_empty_n == 1'b0) | (resetMaximum6_empty_n == 1'b0) | (output_indices_15_empty_n == 1'b0) | (output_indices_04_empty_n == 1'b0)) & (1'b1 == ap_CS_fsm_state2)))) begin
        grp_fu_110_ce = 1'b1;
    end else begin
        grp_fu_110_ce = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        output_indices_04_blk_n = output_indices_04_empty_n;
    end else begin
        output_indices_04_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((storeOutput7_empty_n == 1'b0) | (resetMaximum6_empty_n == 1'b0) | (output_indices_15_empty_n == 1'b0) | (output_indices_04_empty_n == 1'b0)) & (1'b1 == ap_CS_fsm_state2))) begin
        output_indices_04_read = 1'b1;
    end else begin
        output_indices_04_read = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        output_indices_15_blk_n = output_indices_15_empty_n;
    end else begin
        output_indices_15_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((storeOutput7_empty_n == 1'b0) | (resetMaximum6_empty_n == 1'b0) | (output_indices_15_empty_n == 1'b0) | (output_indices_04_empty_n == 1'b0)) & (1'b1 == ap_CS_fsm_state2))) begin
        output_indices_15_read = 1'b1;
    end else begin
        output_indices_15_read = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        resetMaximum6_blk_n = resetMaximum6_empty_n;
    end else begin
        resetMaximum6_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((storeOutput7_empty_n == 1'b0) | (resetMaximum6_empty_n == 1'b0) | (output_indices_15_empty_n == 1'b0) | (output_indices_04_empty_n == 1'b0)) & (1'b1 == ap_CS_fsm_state2))) begin
        resetMaximum6_read = 1'b1;
    end else begin
        resetMaximum6_read = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        storeOutput7_blk_n = storeOutput7_empty_n;
    end else begin
        storeOutput7_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((storeOutput7_empty_n == 1'b0) | (resetMaximum6_empty_n == 1'b0) | (output_indices_15_empty_n == 1'b0) | (output_indices_04_empty_n == 1'b0)) & (1'b1 == ap_CS_fsm_state2))) begin
        storeOutput7_read = 1'b1;
    end else begin
        storeOutput7_read = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_state2 : begin
            if ((~((storeOutput7_empty_n == 1'b0) | (resetMaximum6_empty_n == 1'b0) | (output_indices_15_empty_n == 1'b0) | (output_indices_04_empty_n == 1'b0)) & (storeOutput7_read_read_fu_82_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state2))) begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end else if ((~((storeOutput7_empty_n == 1'b0) | (resetMaximum6_empty_n == 1'b0) | (output_indices_15_empty_n == 1'b0) | (output_indices_04_empty_n == 1'b0)) & (storeOutput7_read_read_fu_82_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end
        end
        ap_ST_fsm_state3 : begin
            ap_NS_fsm = ap_ST_fsm_state4;
        end
        ap_ST_fsm_state4 : begin
            if (((1'b1 == ap_CS_fsm_state4) & (1'b0 == ap_block_state4_on_subcall_done))) begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (ap_done_reg == 1'b1));
end

always @ (*) begin
    ap_block_state2 = ((storeOutput7_empty_n == 1'b0) | (resetMaximum6_empty_n == 1'b0) | (output_indices_15_empty_n == 1'b0) | (output_indices_04_empty_n == 1'b0));
end

always @ (*) begin
    ap_block_state4_on_subcall_done = ((grp_tdf8_writeOutputs_unaligned_fu_88_ap_done == 1'b0) & (storeOutput7_read_reg_157 == 1'd1));
end

assign grp_tdf8_writeOutputs_unaligned_fu_88_ap_start = grp_tdf8_writeOutputs_unaligned_fu_88_ap_start_reg;

assign or_ln24_fu_120_p2 = (resetMaximum6_dout | grp_fu_110_p2);

assign out_data_address1 = grp_tdf8_writeOutputs_unaligned_fu_88_out_data_address1;

assign out_data_ce1 = grp_tdf8_writeOutputs_unaligned_fu_88_out_data_ce1;

assign out_data_d1 = grp_tdf8_writeOutputs_unaligned_fu_88_out_data_d1;

assign out_data_we1 = grp_tdf8_writeOutputs_unaligned_fu_88_out_data_we1;

assign select_ln24_fu_126_p3 = ((or_ln24_fu_120_p2[0:0] == 1'b1) ? p_read : max_vals_0);

assign storeOutput7_read_read_fu_82_p2 = storeOutput7_dout;

endmodule //td_fused_top_tdf8_poolOutputs
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf8_readFilters56 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        filter_data_address0,
        filter_data_ce0,
        filter_data_q0,
        input_indices_23_dout,
        input_indices_23_empty_n,
        input_indices_23_read,
        weight_vecs_0_address0,
        weight_vecs_0_ce0,
        weight_vecs_0_we0,
        weight_vecs_0_d0
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state7 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [16:0] filter_data_address0;
output   filter_data_ce0;
input  [15:0] filter_data_q0;
input  [7:0] input_indices_23_dout;
input   input_indices_23_empty_n;
output   input_indices_23_read;
output  [8:0] weight_vecs_0_address0;
output   weight_vecs_0_ce0;
output   weight_vecs_0_we0;
output  [15:0] weight_vecs_0_d0;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg filter_data_ce0;
reg input_indices_23_read;
reg weight_vecs_0_ce0;
reg weight_vecs_0_we0;

reg    ap_done_reg;
  reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    input_indices_23_blk_n;
reg   [8:0] indvar_flatten13_reg_123;
reg   [1:0] ii_reg_134;
reg   [7:0] indvar_flatten_reg_145;
reg   [1:0] jj_reg_156;
reg   [5:0] kk_reg_167;
wire   [11:0] sext_ln47_fu_200_p1;
reg   [11:0] sext_ln47_reg_408;
wire   [8:0] add_ln47_1_fu_204_p2;
wire    ap_CS_fsm_pp0_stage0;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
wire    ap_block_state4_pp0_stage0_iter2;
wire    ap_block_state5_pp0_stage0_iter3;
wire    ap_block_state6_pp0_stage0_iter4;
wire    ap_block_pp0_stage0_11001;
wire   [0:0] icmp_ln47_fu_210_p2;
reg   [0:0] icmp_ln47_reg_418;
reg   [0:0] icmp_ln47_reg_418_pp0_iter1_reg;
reg   [0:0] icmp_ln47_reg_418_pp0_iter2_reg;
reg   [0:0] icmp_ln47_reg_418_pp0_iter3_reg;
wire   [0:0] icmp_ln48_fu_222_p2;
reg   [0:0] icmp_ln48_reg_422;
wire   [1:0] select_ln47_1_fu_228_p3;
reg   [1:0] select_ln47_1_reg_429;
wire   [7:0] select_ln48_2_fu_242_p3;
wire   [1:0] select_ln48_1_fu_329_p3;
reg   [1:0] select_ln48_1_reg_442;
reg    ap_enable_reg_pp0_iter1;
wire   [8:0] add_ln55_4_fu_392_p2;
reg   [8:0] add_ln55_4_reg_452;
reg   [8:0] add_ln55_4_reg_452_pp0_iter2_reg;
reg   [8:0] add_ln55_4_reg_452_pp0_iter3_reg;
wire   [5:0] add_ln49_fu_398_p2;
reg    ap_block_state1;
wire    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_flush_enable;
reg    ap_enable_reg_pp0_iter2;
reg    ap_condition_pp0_exit_iter1_state3;
reg    ap_enable_reg_pp0_iter3;
reg    ap_enable_reg_pp0_iter4;
reg   [1:0] ap_phi_mux_ii_phi_fu_138_p4;
wire    ap_block_pp0_stage0;
reg   [1:0] ap_phi_mux_jj_phi_fu_160_p4;
wire   [63:0] zext_ln55_9_fu_387_p1;
wire   [63:0] zext_ln55_10_fu_404_p1;
wire   [9:0] tmp_fu_182_p3;
wire   [10:0] zext_ln55_2_fu_190_p1;
wire   [10:0] zext_ln55_fu_178_p1;
wire   [10:0] sub_ln55_fu_194_p2;
wire   [1:0] add_ln47_fu_216_p2;
wire   [7:0] add_ln48_1_fu_236_p2;
wire   [11:0] zext_ln55_4_fu_260_p1;
wire   [11:0] add_ln55_fu_263_p2;
wire   [11:0] shl_ln55_fu_268_p2;
wire   [3:0] tmp_s_fu_280_p3;
wire   [3:0] zext_ln55_3_fu_257_p1;
wire   [0:0] icmp_ln49_fu_298_p2;
wire   [0:0] xor_ln47_fu_293_p2;
wire   [1:0] select_ln47_fu_250_p3;
wire   [0:0] and_ln47_fu_304_p2;
wire   [0:0] or_ln48_fu_316_p2;
wire   [1:0] add_ln48_fu_310_p2;
wire   [11:0] sub_ln55_1_fu_274_p2;
wire   [11:0] zext_ln55_6_fu_341_p1;
wire   [11:0] add_ln55_1_fu_345_p2;
wire   [3:0] sub_ln55_2_fu_287_p2;
wire   [3:0] zext_ln55_5_fu_337_p1;
wire   [3:0] add_ln55_2_fu_359_p2;
wire   [5:0] select_ln48_fu_321_p3;
wire   [16:0] tmp_24_cast_fu_351_p3;
wire   [16:0] zext_ln55_8_fu_377_p1;
wire   [16:0] add_ln55_3_fu_381_p2;
wire   [8:0] tmp_26_cast_fu_365_p3;
wire   [8:0] zext_ln55_7_fu_373_p1;
wire    ap_CS_fsm_state7;
reg   [2:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
#0 ap_enable_reg_pp0_iter4 = 1'b0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state7)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if ((1'b1 == ap_condition_pp0_flush_enable)) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((~((ap_start == 1'b0) | (input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            if ((1'b1 == ap_condition_pp0_exit_iter1_state3)) begin
                ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter0;
            end else if ((1'b1 == 1'b1)) begin
                ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
            end
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter4 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
        end else if ((~((ap_start == 1'b0) | (input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter4 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln47_reg_418 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ii_reg_134 <= select_ln47_1_reg_429;
    end else if ((~((ap_start == 1'b0) | (input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ii_reg_134 <= 2'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_fu_210_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        indvar_flatten13_reg_123 <= add_ln47_1_fu_204_p2;
    end else if ((~((ap_start == 1'b0) | (input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indvar_flatten13_reg_123 <= 9'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_fu_210_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        indvar_flatten_reg_145 <= select_ln48_2_fu_242_p3;
    end else if ((~((ap_start == 1'b0) | (input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indvar_flatten_reg_145 <= 8'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_reg_418_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        jj_reg_156 <= select_ln48_1_reg_442;
    end else if ((~((ap_start == 1'b0) | (input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        jj_reg_156 <= 2'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln47_reg_418 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        kk_reg_167 <= add_ln49_fu_398_p2;
    end else if ((~((ap_start == 1'b0) | (input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        kk_reg_167 <= 6'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_reg_418 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        add_ln55_4_reg_452 <= add_ln55_4_fu_392_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        add_ln55_4_reg_452_pp0_iter2_reg <= add_ln55_4_reg_452;
        add_ln55_4_reg_452_pp0_iter3_reg <= add_ln55_4_reg_452_pp0_iter2_reg;
        icmp_ln47_reg_418_pp0_iter2_reg <= icmp_ln47_reg_418_pp0_iter1_reg;
        icmp_ln47_reg_418_pp0_iter3_reg <= icmp_ln47_reg_418_pp0_iter2_reg;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln47_reg_418 <= icmp_ln47_fu_210_p2;
        icmp_ln47_reg_418_pp0_iter1_reg <= icmp_ln47_reg_418;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_fu_210_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln48_reg_422 <= icmp_ln48_fu_222_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln47_fu_210_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        select_ln47_1_reg_429 <= select_ln47_1_fu_228_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln47_reg_418 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        select_ln48_1_reg_442 <= select_ln48_1_fu_329_p3;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state1)) begin
        sext_ln47_reg_408 <= sext_ln47_fu_200_p1;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_condition_pp0_exit_iter1_state3 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter1_state3 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln47_fu_210_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_condition_pp0_flush_enable = 1'b1;
    end else begin
        ap_condition_pp0_flush_enable = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state7)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln47_reg_418 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_phi_mux_ii_phi_fu_138_p4 = select_ln47_1_reg_429;
    end else begin
        ap_phi_mux_ii_phi_fu_138_p4 = ii_reg_134;
    end
end

always @ (*) begin
    if (((icmp_ln47_reg_418_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        ap_phi_mux_jj_phi_fu_160_p4 = select_ln48_1_reg_442;
    end else begin
        ap_phi_mux_jj_phi_fu_160_p4 = jj_reg_156;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state7)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter3 == 1'b1)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter4 == 1'b1)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1)))) begin
        filter_data_ce0 = 1'b1;
    end else begin
        filter_data_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        input_indices_23_blk_n = input_indices_23_empty_n;
    end else begin
        input_indices_23_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        input_indices_23_read = 1'b1;
    end else begin
        input_indices_23_read = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter4 == 1'b1))) begin
        weight_vecs_0_ce0 = 1'b1;
    end else begin
        weight_vecs_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln47_reg_418_pp0_iter3_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter4 == 1'b1))) begin
        weight_vecs_0_we0 = 1'b1;
    end else begin
        weight_vecs_0_we0 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_start == 1'b0) | (input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((~((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b0)) & ~((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter4 == 1'b1) & (ap_enable_reg_pp0_iter3 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if ((((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b0)) | ((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter4 == 1'b1) & (ap_enable_reg_pp0_iter3 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_state7;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state7 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln47_1_fu_204_p2 = (indvar_flatten13_reg_123 + 9'd1);

assign add_ln47_fu_216_p2 = (ap_phi_mux_ii_phi_fu_138_p4 + 2'd1);

assign add_ln48_1_fu_236_p2 = (indvar_flatten_reg_145 + 8'd1);

assign add_ln48_fu_310_p2 = (select_ln47_fu_250_p3 + 2'd1);

assign add_ln49_fu_398_p2 = (select_ln48_fu_321_p3 + 6'd1);

assign add_ln55_1_fu_345_p2 = (sub_ln55_1_fu_274_p2 + zext_ln55_6_fu_341_p1);

assign add_ln55_2_fu_359_p2 = (sub_ln55_2_fu_287_p2 + zext_ln55_5_fu_337_p1);

assign add_ln55_3_fu_381_p2 = (tmp_24_cast_fu_351_p3 + zext_ln55_8_fu_377_p1);

assign add_ln55_4_fu_392_p2 = (tmp_26_cast_fu_365_p3 + zext_ln55_7_fu_373_p1);

assign add_ln55_fu_263_p2 = ((sext_ln47_reg_408) + (zext_ln55_4_fu_260_p1));

assign and_ln47_fu_304_p2 = (xor_ln47_fu_293_p2 & icmp_ln49_fu_298_p2);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state7 = ap_CS_fsm[32'd2];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (input_indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1));
end

assign ap_block_state2_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter4 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign filter_data_address0 = zext_ln55_9_fu_387_p1;

assign icmp_ln47_fu_210_p2 = ((indvar_flatten13_reg_123 == 9'd288) ? 1'b1 : 1'b0);

assign icmp_ln48_fu_222_p2 = ((indvar_flatten_reg_145 == 8'd96) ? 1'b1 : 1'b0);

assign icmp_ln49_fu_298_p2 = ((kk_reg_167 == 6'd32) ? 1'b1 : 1'b0);

assign or_ln48_fu_316_p2 = (icmp_ln48_reg_422 | and_ln47_fu_304_p2);

assign select_ln47_1_fu_228_p3 = ((icmp_ln48_fu_222_p2[0:0] == 1'b1) ? add_ln47_fu_216_p2 : ap_phi_mux_ii_phi_fu_138_p4);

assign select_ln47_fu_250_p3 = ((icmp_ln48_reg_422[0:0] == 1'b1) ? 2'd0 : ap_phi_mux_jj_phi_fu_160_p4);

assign select_ln48_1_fu_329_p3 = ((and_ln47_fu_304_p2[0:0] == 1'b1) ? add_ln48_fu_310_p2 : select_ln47_fu_250_p3);

assign select_ln48_2_fu_242_p3 = ((icmp_ln48_fu_222_p2[0:0] == 1'b1) ? 8'd1 : add_ln48_1_fu_236_p2);

assign select_ln48_fu_321_p3 = ((or_ln48_fu_316_p2[0:0] == 1'b1) ? 6'd0 : kk_reg_167);

assign sext_ln47_fu_200_p1 = (sub_ln55_fu_194_p2);

assign shl_ln55_fu_268_p2 = add_ln55_fu_263_p2 << 12'd2;

assign sub_ln55_1_fu_274_p2 = (shl_ln55_fu_268_p2 - add_ln55_fu_263_p2);

assign sub_ln55_2_fu_287_p2 = (tmp_s_fu_280_p3 - zext_ln55_3_fu_257_p1);

assign sub_ln55_fu_194_p2 = (zext_ln55_2_fu_190_p1 - zext_ln55_fu_178_p1);

assign tmp_24_cast_fu_351_p3 = {{add_ln55_1_fu_345_p2}, {5'd0}};

assign tmp_26_cast_fu_365_p3 = {{add_ln55_2_fu_359_p2}, {5'd0}};

assign tmp_fu_182_p3 = {{input_indices_23_dout}, {2'd0}};

assign tmp_s_fu_280_p3 = {{select_ln47_1_reg_429}, {2'd0}};

assign weight_vecs_0_address0 = zext_ln55_10_fu_404_p1;

assign weight_vecs_0_d0 = filter_data_q0;

assign xor_ln47_fu_293_p2 = (icmp_ln48_reg_422 ^ 1'd1);

assign zext_ln55_10_fu_404_p1 = add_ln55_4_reg_452_pp0_iter3_reg;

assign zext_ln55_2_fu_190_p1 = tmp_fu_182_p3;

assign zext_ln55_3_fu_257_p1 = select_ln47_1_reg_429;

assign zext_ln55_4_fu_260_p1 = select_ln47_1_reg_429;

assign zext_ln55_5_fu_337_p1 = select_ln48_1_fu_329_p3;

assign zext_ln55_6_fu_341_p1 = select_ln48_1_fu_329_p3;

assign zext_ln55_7_fu_373_p1 = select_ln48_fu_321_p3;

assign zext_ln55_8_fu_377_p1 = select_ln48_fu_321_p3;

assign zext_ln55_9_fu_387_p1 = add_ln55_3_fu_381_p2;

assign zext_ln55_fu_178_p1 = input_indices_23_dout;

endmodule //td_fused_top_tdf8_readFilters56
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf8_readInputs57 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        in_data_address0,
        in_data_ce0,
        in_data_q0,
        i_13,
        j_13,
        ifmap_vec_address0,
        ifmap_vec_ce0,
        ifmap_vec_we0,
        ifmap_vec_d0,
        ifmap_vec_address1,
        ifmap_vec_ce1,
        ifmap_vec_we1,
        ifmap_vec_d1
);

parameter    ap_ST_fsm_state1 = 4'd1;
parameter    ap_ST_fsm_pp0_stage0 = 4'd2;
parameter    ap_ST_fsm_pp0_stage1 = 4'd4;
parameter    ap_ST_fsm_state8 = 4'd8;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [12:0] in_data_address0;
output   in_data_ce0;
input  [63:0] in_data_q0;
input  [15:0] i_13;
input  [15:0] j_13;
output  [8:0] ifmap_vec_address0;
output   ifmap_vec_ce0;
output   ifmap_vec_we0;
output  [15:0] ifmap_vec_d0;
output  [8:0] ifmap_vec_address1;
output   ifmap_vec_ce1;
output   ifmap_vec_we1;
output  [15:0] ifmap_vec_d1;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg in_data_ce0;
reg[8:0] ifmap_vec_address0;
reg ifmap_vec_ce0;
reg ifmap_vec_we0;
reg[15:0] ifmap_vec_d0;
reg[8:0] ifmap_vec_address1;
reg ifmap_vec_ce1;
reg ifmap_vec_we1;
reg[15:0] ifmap_vec_d1;

reg    ap_done_reg;
  reg   [3:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg   [6:0] indvar_flatten47_reg_192;
reg   [1:0] ii_reg_204;
reg   [5:0] indvar_flatten_reg_216;
reg   [1:0] jj_reg_227;
reg   [5:0] kk_0_i_reg_239;
wire   [17:0] p_cast_i_fu_268_p1;
reg   [17:0] p_cast_i_reg_929;
wire   [9:0] trunc_ln22_fu_272_p1;
reg   [9:0] trunc_ln22_reg_935;
wire   [17:0] sext_ln22_fu_282_p1;
reg   [17:0] sext_ln22_reg_941;
wire   [4:0] p_cast_fu_286_p2;
reg   [4:0] p_cast_reg_947;
wire   [0:0] or_ln23_1_fu_306_p2;
reg   [0:0] or_ln23_1_reg_953;
wire   [9:0] p_mid137_fu_312_p2;
reg   [9:0] p_mid137_reg_958;
wire   [4:0] p_cast5_i_fu_331_p2;
reg   [4:0] p_cast5_i_reg_963;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state4_pp0_stage0_iter1;
wire    ap_block_state6_pp0_stage0_iter2;
wire    ap_block_pp0_stage0_11001;
wire   [0:0] is_padding_fu_371_p2;
reg   [0:0] is_padding_reg_969;
wire   [0:0] icmp_ln19_fu_377_p2;
reg   [0:0] icmp_ln19_reg_976;
reg   [0:0] icmp_ln19_reg_976_pp0_iter1_reg;
reg   [0:0] icmp_ln19_reg_976_pp0_iter2_reg;
wire   [1:0] add_ln19_fu_383_p2;
reg   [1:0] add_ln19_reg_980;
wire   [0:0] icmp_ln20_fu_389_p2;
reg   [0:0] icmp_ln20_reg_985;
wire   [1:0] select_ln19_fu_395_p3;
reg   [1:0] select_ln19_reg_997;
wire   [4:0] p_cast5_i_mid1_fu_416_p2;
reg   [4:0] p_cast5_i_mid1_reg_1002;
wire   [0:0] or_ln23_3_fu_435_p2;
reg   [0:0] or_ln23_3_reg_1008;
wire   [1:0] add_ln20_fu_440_p2;
reg   [1:0] add_ln20_reg_1015;
wire   [0:0] or_ln23_5_fu_475_p2;
reg   [0:0] or_ln23_5_reg_1021;
wire   [5:0] add_ln20_1_fu_481_p2;
reg   [5:0] add_ln20_1_reg_1028;
wire   [6:0] add_ln19_1_fu_487_p2;
reg   [6:0] add_ln19_1_reg_1033;
wire    ap_CS_fsm_pp0_stage1;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_state3_pp0_stage1_iter0;
wire    ap_block_state5_pp0_stage1_iter1;
wire    ap_block_state7_pp0_stage1_iter2;
wire    ap_block_pp0_stage1_11001;
wire   [1:0] select_ln19_1_fu_525_p3;
reg   [1:0] select_ln19_1_reg_1038;
wire   [5:0] select_ln20_fu_589_p3;
reg   [5:0] select_ln20_reg_1045;
wire   [1:0] select_ln20_1_fu_597_p3;
reg   [1:0] select_ln20_1_reg_1051;
wire   [0:0] select_ln20_2_fu_606_p3;
reg   [0:0] select_ln20_2_reg_1057;
reg   [0:0] select_ln20_2_reg_1057_pp0_iter1_reg;
wire   [4:0] empty_63_fu_702_p1;
reg   [4:0] empty_63_reg_1065;
reg   [4:0] empty_63_reg_1065_pp0_iter1_reg;
wire   [5:0] select_ln20_5_fu_729_p3;
reg   [5:0] select_ln20_5_reg_1077;
wire   [5:0] add_ln25_fu_735_p2;
reg   [5:0] add_ln25_reg_1082;
reg    ap_enable_reg_pp0_iter1;
wire   [5:0] add_ln33_fu_767_p2;
reg   [5:0] add_ln33_reg_1087;
wire   [8:0] add_ln33_1_fu_788_p2;
reg   [8:0] add_ln33_1_reg_1094;
wire   [15:0] select_ln33_5_fu_867_p3;
reg   [15:0] select_ln33_5_reg_1099;
wire   [15:0] select_ln33_6_fu_888_p3;
reg   [15:0] select_ln33_6_reg_1104;
reg    ap_block_state1;
wire    ap_block_pp0_stage1_subdone;
reg    ap_condition_pp0_exit_iter0_state3;
reg    ap_enable_reg_pp0_iter2;
reg   [6:0] ap_phi_mux_indvar_flatten47_phi_fu_196_p4;
wire    ap_block_pp0_stage0;
reg   [1:0] ap_phi_mux_ii_phi_fu_208_p4;
reg   [5:0] ap_phi_mux_indvar_flatten_phi_fu_220_p4;
reg   [1:0] ap_phi_mux_jj_phi_fu_231_p4;
reg   [5:0] ap_phi_mux_kk_0_i_phi_fu_243_p4;
wire    ap_block_pp0_stage1;
wire   [63:0] sext_ln32_fu_724_p1;
wire   [63:0] zext_ln33_5_fu_794_p1;
wire   [63:0] sext_ln33_fu_826_p1;
wire   [63:0] sext_ln33_1_fu_907_p1;
wire   [63:0] sext_ln33_2_fu_924_p1;
wire   [15:0] select_ln33_fu_806_p3;
wire   [15:0] select_ln33_4_fu_845_p3;
wire   [16:0] zext_ln19_fu_254_p1;
wire   [16:0] empty_58_fu_262_p2;
wire   [16:0] j_cast_i_fu_250_p1;
wire   [16:0] add_ln22_fu_276_p2;
wire   [4:0] empty_fu_258_p1;
wire   [0:0] tmp_fu_292_p3;
wire   [0:0] icmp_ln24_fu_300_p2;
wire   [17:0] ii_cast_i_fu_318_p1;
wire   [4:0] ii_cast_fu_322_p1;
wire   [17:0] empty_59_fu_326_p2;
wire   [17:0] zext_ln20_fu_342_p1;
wire   [17:0] add_ln22_1_fu_346_p2;
wire   [0:0] tmp_3_fu_351_p3;
wire   [0:0] icmp_ln24_1_fu_359_p2;
wire   [0:0] or_ln23_fu_365_p2;
wire   [0:0] empty_60_fu_336_p2;
wire   [17:0] ii_cast_i_mid1_fu_403_p1;
wire   [4:0] ii_cast_mid1_fu_407_p1;
wire   [17:0] p_mid111_fu_411_p2;
wire   [0:0] p_mid113_fu_421_p2;
wire   [17:0] zext_ln20_1_fu_446_p1;
wire   [17:0] add_ln22_2_fu_450_p2;
wire   [0:0] tmp_4_fu_455_p3;
wire   [0:0] icmp_ln24_2_fu_463_p2;
wire   [0:0] or_ln23_4_fu_469_p2;
wire   [0:0] select_ln19_3_fu_427_p3;
wire   [2:0] zext_ln22_fu_493_p1;
wire   [2:0] tmp2_fu_503_p2;
wire   [9:0] tmp2_cast_fu_509_p1;
wire   [9:0] empty_61_fu_513_p2;
wire   [4:0] row_coord_int_mid131_fu_541_p3;
wire   [4:0] row_coord_int_fu_497_p3;
wire   [9:0] col_coord_int_mid139_fu_547_p3;
wire   [9:0] col_coord_int_fu_518_p3;
wire   [0:0] icmp_ln25_fu_572_p2;
wire   [0:0] xor_ln19_fu_567_p2;
wire   [0:0] and_ln19_fu_578_p2;
wire   [0:0] or_ln20_fu_584_p2;
wire   [0:0] select_ln19_4_fu_536_p3;
wire   [4:0] select_ln19_2_fu_531_p3;
wire   [2:0] zext_ln22_1_fu_603_p1;
wire   [2:0] tmp2_mid1_fu_620_p2;
wire   [9:0] tmp2_cast_mid1_fu_626_p1;
wire   [9:0] p_mid1_fu_630_p2;
wire   [4:0] row_coord_int_mid1_fu_613_p3;
wire   [4:0] select_ln19_5_fu_553_p3;
wire   [4:0] select_ln20_3_fu_642_p3;
wire   [9:0] tmp_1_fu_650_p3;
wire   [6:0] tmp_2_fu_662_p3;
wire   [10:0] zext_ln32_fu_658_p1;
wire   [10:0] zext_ln32_7_fu_670_p1;
wire   [10:0] sub_ln32_fu_674_p2;
wire   [9:0] col_coord_int_mid1_fu_635_p3;
wire   [9:0] select_ln19_6_fu_560_p3;
wire   [9:0] select_ln20_4_fu_684_p3;
wire   [11:0] sext_ln20_fu_680_p1;
wire   [11:0] zext_ln32_8_fu_692_p1;
wire   [11:0] add_ln32_fu_696_p2;
wire   [2:0] lshr_ln_fu_706_p4;
wire   [14:0] tmp_5_fu_716_p3;
wire   [3:0] tmp_s_fu_743_p3;
wire   [4:0] zext_ln33_2_fu_750_p1;
wire   [4:0] zext_ln33_fu_740_p1;
wire   [4:0] sub_ln33_fu_754_p2;
wire   [5:0] sub_ln33_cast_fu_760_p1;
wire   [5:0] zext_ln33_3_fu_764_p1;
wire   [3:0] trunc_ln33_fu_773_p1;
wire   [8:0] tmp_13_cast_fu_777_p3;
wire   [8:0] zext_ln33_4_fu_785_p1;
wire   [15:0] trunc_ln32_fu_798_p1;
wire   [15:0] bitcast_ln32_fu_802_p1;
wire   [4:0] or_ln25_fu_814_p2;
wire   [10:0] tmp_6_fu_819_p3;
wire   [15:0] tmp_12_i_fu_831_p4;
wire   [15:0] bitcast_ln32_4_fu_841_p1;
wire   [15:0] tmp_13_i_fu_853_p4;
wire   [15:0] bitcast_ln32_5_fu_863_p1;
wire   [15:0] tmp_14_i_fu_874_p4;
wire   [15:0] bitcast_ln32_6_fu_884_p1;
wire   [4:0] or_ln25_3_fu_895_p2;
wire   [10:0] tmp_7_fu_900_p3;
wire   [4:0] or_ln25_4_fu_912_p2;
wire   [10:0] tmp_8_fu_917_p3;
wire    ap_CS_fsm_state8;
reg   [3:0] ap_NS_fsm;
wire    ap_block_pp0_stage0_subdone;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 4'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_condition_pp0_exit_iter0_state3) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            if ((1'b1 == ap_condition_pp0_exit_iter0_state3)) begin
                ap_enable_reg_pp0_iter1 <= (1'b1 ^ ap_condition_pp0_exit_iter0_state3);
            end else if ((1'b1 == 1'b1)) begin
                ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
            end
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter2 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln19_reg_976 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ii_reg_204 <= select_ln19_1_reg_1038;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ii_reg_204 <= 2'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln19_reg_976 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        indvar_flatten47_reg_192 <= add_ln19_1_reg_1033;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indvar_flatten47_reg_192 <= 7'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln19_reg_976 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        indvar_flatten_reg_216 <= select_ln20_5_reg_1077;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indvar_flatten_reg_216 <= 6'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln19_reg_976 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        jj_reg_227 <= select_ln20_1_reg_1051;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        jj_reg_227 <= 2'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln19_reg_976_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        kk_0_i_reg_239 <= add_ln25_reg_1082;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        kk_0_i_reg_239 <= 6'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
        add_ln19_1_reg_1033 <= add_ln19_1_fu_487_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln19_fu_377_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        add_ln19_reg_980 <= add_ln19_fu_383_p2;
        add_ln20_1_reg_1028 <= add_ln20_1_fu_481_p2;
        add_ln20_reg_1015 <= add_ln20_fu_440_p2;
        icmp_ln20_reg_985 <= icmp_ln20_fu_389_p2;
        or_ln23_3_reg_1008 <= or_ln23_3_fu_435_p2;
        or_ln23_5_reg_1021 <= or_ln23_5_fu_475_p2;
        p_cast5_i_mid1_reg_1002 <= p_cast5_i_mid1_fu_416_p2;
        select_ln19_reg_997 <= select_ln19_fu_395_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln19_reg_976 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        add_ln25_reg_1082 <= add_ln25_fu_735_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln19_reg_976_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
        add_ln33_1_reg_1094 <= add_ln33_1_fu_788_p2;
        add_ln33_reg_1087 <= add_ln33_fu_767_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln19_reg_976 == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
        empty_63_reg_1065 <= empty_63_fu_702_p1;
        select_ln20_2_reg_1057 <= select_ln20_2_fu_606_p3;
        select_ln20_reg_1045 <= select_ln20_fu_589_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
        empty_63_reg_1065_pp0_iter1_reg <= empty_63_reg_1065;
        select_ln20_2_reg_1057_pp0_iter1_reg <= select_ln20_2_reg_1057;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln19_reg_976 <= icmp_ln19_fu_377_p2;
        icmp_ln19_reg_976_pp0_iter1_reg <= icmp_ln19_reg_976;
        icmp_ln19_reg_976_pp0_iter2_reg <= icmp_ln19_reg_976_pp0_iter1_reg;
        is_padding_reg_969 <= is_padding_fu_371_p2;
        p_cast5_i_reg_963 <= p_cast5_i_fu_331_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state1)) begin
        or_ln23_1_reg_953 <= or_ln23_1_fu_306_p2;
        p_cast_i_reg_929 <= p_cast_i_fu_268_p1;
        p_cast_reg_947 <= p_cast_fu_286_p2;
        p_mid137_reg_958 <= p_mid137_fu_312_p2;
        sext_ln22_reg_941 <= sext_ln22_fu_282_p1;
        trunc_ln22_reg_935 <= trunc_ln22_fu_272_p1;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln19_reg_976 == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
        select_ln19_1_reg_1038 <= select_ln19_1_fu_525_p3;
        select_ln20_1_reg_1051 <= select_ln20_1_fu_597_p3;
        select_ln20_5_reg_1077 <= select_ln20_5_fu_729_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln19_reg_976_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        select_ln33_5_reg_1099 <= select_ln33_5_fu_867_p3;
        select_ln33_6_reg_1104 <= select_ln33_6_fu_888_p3;
    end
end

always @ (*) begin
    if ((icmp_ln19_reg_976 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state3 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state3 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state8)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln19_reg_976 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_ii_phi_fu_208_p4 = select_ln19_1_reg_1038;
    end else begin
        ap_phi_mux_ii_phi_fu_208_p4 = ii_reg_204;
    end
end

always @ (*) begin
    if (((icmp_ln19_reg_976 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_indvar_flatten47_phi_fu_196_p4 = add_ln19_1_reg_1033;
    end else begin
        ap_phi_mux_indvar_flatten47_phi_fu_196_p4 = indvar_flatten47_reg_192;
    end
end

always @ (*) begin
    if (((icmp_ln19_reg_976 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_indvar_flatten_phi_fu_220_p4 = select_ln20_5_reg_1077;
    end else begin
        ap_phi_mux_indvar_flatten_phi_fu_220_p4 = indvar_flatten_reg_216;
    end
end

always @ (*) begin
    if (((icmp_ln19_reg_976 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_jj_phi_fu_231_p4 = select_ln20_1_reg_1051;
    end else begin
        ap_phi_mux_jj_phi_fu_231_p4 = jj_reg_227;
    end
end

always @ (*) begin
    if (((icmp_ln19_reg_976_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_kk_0_i_phi_fu_243_p4 = add_ln25_reg_1082;
    end else begin
        ap_phi_mux_kk_0_i_phi_fu_243_p4 = kk_0_i_reg_239;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state8)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((ap_enable_reg_pp0_iter2 == 1'b1)) begin
        if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            ifmap_vec_address0 = sext_ln33_2_fu_924_p1;
        end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ifmap_vec_address0 = sext_ln33_fu_826_p1;
        end else begin
            ifmap_vec_address0 = 'bx;
        end
    end else begin
        ifmap_vec_address0 = 'bx;
    end
end

always @ (*) begin
    if ((ap_enable_reg_pp0_iter2 == 1'b1)) begin
        if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            ifmap_vec_address1 = sext_ln33_1_fu_907_p1;
        end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ifmap_vec_address1 = zext_ln33_5_fu_794_p1;
        end else begin
            ifmap_vec_address1 = 'bx;
        end
    end else begin
        ifmap_vec_address1 = 'bx;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1)) | ((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter2 == 1'b1)))) begin
        ifmap_vec_ce0 = 1'b1;
    end else begin
        ifmap_vec_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1)) | ((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter2 == 1'b1)))) begin
        ifmap_vec_ce1 = 1'b1;
    end else begin
        ifmap_vec_ce1 = 1'b0;
    end
end

always @ (*) begin
    if ((ap_enable_reg_pp0_iter2 == 1'b1)) begin
        if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            ifmap_vec_d0 = select_ln33_6_reg_1104;
        end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ifmap_vec_d0 = select_ln33_4_fu_845_p3;
        end else begin
            ifmap_vec_d0 = 'bx;
        end
    end else begin
        ifmap_vec_d0 = 'bx;
    end
end

always @ (*) begin
    if ((ap_enable_reg_pp0_iter2 == 1'b1)) begin
        if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            ifmap_vec_d1 = select_ln33_5_reg_1099;
        end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ifmap_vec_d1 = select_ln33_fu_806_p3;
        end else begin
            ifmap_vec_d1 = 'bx;
        end
    end else begin
        ifmap_vec_d1 = 'bx;
    end
end

always @ (*) begin
    if ((((icmp_ln19_reg_976_pp0_iter2_reg == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter2 == 1'b1)) | ((icmp_ln19_reg_976_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1)))) begin
        ifmap_vec_we0 = 1'b1;
    end else begin
        ifmap_vec_we0 = 1'b0;
    end
end

always @ (*) begin
    if ((((icmp_ln19_reg_976_pp0_iter2_reg == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter2 == 1'b1)) | ((icmp_ln19_reg_976_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1)))) begin
        ifmap_vec_we1 = 1'b1;
    end else begin
        ifmap_vec_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1)) | ((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1)) | ((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1)) | ((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1)))) begin
        in_data_ce0 = 1'b1;
    end else begin
        in_data_ce0 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_pp0_stage1 : begin
            if ((~((icmp_ln19_reg_976 == 1'd1) & (1'b0 == ap_block_pp0_stage1_subdone) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1)) & ~((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter2 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0)) & (1'b0 == ap_block_pp0_stage1_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if ((((icmp_ln19_reg_976 == 1'd1) & (1'b0 == ap_block_pp0_stage1_subdone) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1)) | ((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter2 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_state8;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end
        end
        ap_ST_fsm_state8 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln19_1_fu_487_p2 = (indvar_flatten47_reg_192 + 7'd1);

assign add_ln19_fu_383_p2 = (ap_phi_mux_ii_phi_fu_208_p4 + 2'd1);

assign add_ln20_1_fu_481_p2 = (ap_phi_mux_indvar_flatten_phi_fu_220_p4 + 6'd1);

assign add_ln20_fu_440_p2 = (select_ln19_fu_395_p3 + 2'd1);

assign add_ln22_1_fu_346_p2 = ((sext_ln22_reg_941) + (zext_ln20_fu_342_p1));

assign add_ln22_2_fu_450_p2 = ((sext_ln22_reg_941) + (zext_ln20_1_fu_446_p1));

assign add_ln22_fu_276_p2 = ((j_cast_i_fu_250_p1) + (17'd131071));

assign add_ln25_fu_735_p2 = (select_ln20_reg_1045 + 6'd4);

assign add_ln32_fu_696_p2 = ((sext_ln20_fu_680_p1) + (zext_ln32_8_fu_692_p1));

assign add_ln33_1_fu_788_p2 = (tmp_13_cast_fu_777_p3 + zext_ln33_4_fu_785_p1);

assign add_ln33_fu_767_p2 = ((sub_ln33_cast_fu_760_p1) + (zext_ln33_3_fu_764_p1));

assign and_ln19_fu_578_p2 = (xor_ln19_fu_567_p2 & icmp_ln25_fu_572_p2);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_pp0_stage1 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state8 = ap_CS_fsm[32'd3];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (ap_done_reg == 1'b1));
end

assign ap_block_state2_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage1_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage1_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage1_iter2 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign bitcast_ln32_4_fu_841_p1 = tmp_12_i_fu_831_p4;

assign bitcast_ln32_5_fu_863_p1 = tmp_13_i_fu_853_p4;

assign bitcast_ln32_6_fu_884_p1 = tmp_14_i_fu_874_p4;

assign bitcast_ln32_fu_802_p1 = trunc_ln32_fu_798_p1;

assign col_coord_int_fu_518_p3 = ((is_padding_reg_969[0:0] == 1'b1) ? 10'd0 : empty_61_fu_513_p2);

assign col_coord_int_mid139_fu_547_p3 = ((or_ln23_3_reg_1008[0:0] == 1'b1) ? 10'd0 : p_mid137_reg_958);

assign col_coord_int_mid1_fu_635_p3 = ((or_ln23_5_reg_1021[0:0] == 1'b1) ? 10'd0 : p_mid1_fu_630_p2);

assign empty_58_fu_262_p2 = ((zext_ln19_fu_254_p1) + (17'd131071));

assign empty_59_fu_326_p2 = ((p_cast_i_reg_929) + (ii_cast_i_fu_318_p1));

assign empty_60_fu_336_p2 = ((empty_59_fu_326_p2 > 18'd27) ? 1'b1 : 1'b0);

assign empty_61_fu_513_p2 = ((tmp2_cast_fu_509_p1) + (trunc_ln22_reg_935));

assign empty_63_fu_702_p1 = select_ln20_fu_589_p3[4:0];

assign empty_fu_258_p1 = i_13[4:0];

assign icmp_ln19_fu_377_p2 = ((ap_phi_mux_indvar_flatten47_phi_fu_196_p4 == 7'd72) ? 1'b1 : 1'b0);

assign icmp_ln20_fu_389_p2 = ((ap_phi_mux_indvar_flatten_phi_fu_220_p4 == 6'd24) ? 1'b1 : 1'b0);

assign icmp_ln24_1_fu_359_p2 = (((add_ln22_1_fu_346_p2) > (18'd27)) ? 1'b1 : 1'b0);

assign icmp_ln24_2_fu_463_p2 = (((add_ln22_2_fu_450_p2) > (18'd27)) ? 1'b1 : 1'b0);

assign icmp_ln24_fu_300_p2 = (((add_ln22_fu_276_p2) > (17'd27)) ? 1'b1 : 1'b0);

assign icmp_ln25_fu_572_p2 = ((ap_phi_mux_kk_0_i_phi_fu_243_p4 == 6'd32) ? 1'b1 : 1'b0);

assign ii_cast_fu_322_p1 = ap_phi_mux_ii_phi_fu_208_p4;

assign ii_cast_i_fu_318_p1 = ap_phi_mux_ii_phi_fu_208_p4;

assign ii_cast_i_mid1_fu_403_p1 = add_ln19_fu_383_p2;

assign ii_cast_mid1_fu_407_p1 = add_ln19_fu_383_p2;

assign in_data_address0 = sext_ln32_fu_724_p1;

assign is_padding_fu_371_p2 = (or_ln23_fu_365_p2 | empty_60_fu_336_p2);

assign j_cast_i_fu_250_p1 = j_13;

assign lshr_ln_fu_706_p4 = {{select_ln20_fu_589_p3[4:2]}};

assign or_ln20_fu_584_p2 = (icmp_ln20_reg_985 | and_ln19_fu_578_p2);

assign or_ln23_1_fu_306_p2 = (tmp_fu_292_p3 | icmp_ln24_fu_300_p2);

assign or_ln23_3_fu_435_p2 = (p_mid113_fu_421_p2 | or_ln23_1_reg_953);

assign or_ln23_4_fu_469_p2 = (tmp_4_fu_455_p3 | icmp_ln24_2_fu_463_p2);

assign or_ln23_5_fu_475_p2 = (select_ln19_3_fu_427_p3 | or_ln23_4_fu_469_p2);

assign or_ln23_fu_365_p2 = (tmp_3_fu_351_p3 | icmp_ln24_1_fu_359_p2);

assign or_ln25_3_fu_895_p2 = (empty_63_reg_1065_pp0_iter1_reg | 5'd2);

assign or_ln25_4_fu_912_p2 = (empty_63_reg_1065_pp0_iter1_reg | 5'd3);

assign or_ln25_fu_814_p2 = (empty_63_reg_1065_pp0_iter1_reg | 5'd1);

assign p_cast5_i_fu_331_p2 = (p_cast_reg_947 + ii_cast_fu_322_p1);

assign p_cast5_i_mid1_fu_416_p2 = (p_cast_reg_947 + ii_cast_mid1_fu_407_p1);

assign p_cast_fu_286_p2 = ((empty_fu_258_p1) + (5'd31));

assign p_cast_i_fu_268_p1 = (empty_58_fu_262_p2);

assign p_mid111_fu_411_p2 = ((p_cast_i_reg_929) + (ii_cast_i_mid1_fu_403_p1));

assign p_mid113_fu_421_p2 = ((p_mid111_fu_411_p2 > 18'd27) ? 1'b1 : 1'b0);

assign p_mid137_fu_312_p2 = ((trunc_ln22_fu_272_p1) + (10'd1023));

assign p_mid1_fu_630_p2 = ((tmp2_cast_mid1_fu_626_p1) + (trunc_ln22_reg_935));

assign row_coord_int_fu_497_p3 = ((is_padding_reg_969[0:0] == 1'b1) ? 5'd0 : p_cast5_i_reg_963);

assign row_coord_int_mid131_fu_541_p3 = ((or_ln23_3_reg_1008[0:0] == 1'b1) ? 5'd0 : p_cast5_i_mid1_reg_1002);

assign row_coord_int_mid1_fu_613_p3 = ((or_ln23_5_reg_1021[0:0] == 1'b1) ? 5'd0 : select_ln19_2_fu_531_p3);

assign select_ln19_1_fu_525_p3 = ((icmp_ln20_reg_985[0:0] == 1'b1) ? add_ln19_reg_980 : ii_reg_204);

assign select_ln19_2_fu_531_p3 = ((icmp_ln20_reg_985[0:0] == 1'b1) ? p_cast5_i_mid1_reg_1002 : p_cast5_i_reg_963);

assign select_ln19_3_fu_427_p3 = ((icmp_ln20_fu_389_p2[0:0] == 1'b1) ? p_mid113_fu_421_p2 : empty_60_fu_336_p2);

assign select_ln19_4_fu_536_p3 = ((icmp_ln20_reg_985[0:0] == 1'b1) ? or_ln23_3_reg_1008 : is_padding_reg_969);

assign select_ln19_5_fu_553_p3 = ((icmp_ln20_reg_985[0:0] == 1'b1) ? row_coord_int_mid131_fu_541_p3 : row_coord_int_fu_497_p3);

assign select_ln19_6_fu_560_p3 = ((icmp_ln20_reg_985[0:0] == 1'b1) ? col_coord_int_mid139_fu_547_p3 : col_coord_int_fu_518_p3);

assign select_ln19_fu_395_p3 = ((icmp_ln20_fu_389_p2[0:0] == 1'b1) ? 2'd0 : ap_phi_mux_jj_phi_fu_231_p4);

assign select_ln20_1_fu_597_p3 = ((and_ln19_fu_578_p2[0:0] == 1'b1) ? add_ln20_reg_1015 : select_ln19_reg_997);

assign select_ln20_2_fu_606_p3 = ((and_ln19_fu_578_p2[0:0] == 1'b1) ? or_ln23_5_reg_1021 : select_ln19_4_fu_536_p3);

assign select_ln20_3_fu_642_p3 = ((and_ln19_fu_578_p2[0:0] == 1'b1) ? row_coord_int_mid1_fu_613_p3 : select_ln19_5_fu_553_p3);

assign select_ln20_4_fu_684_p3 = ((and_ln19_fu_578_p2[0:0] == 1'b1) ? col_coord_int_mid1_fu_635_p3 : select_ln19_6_fu_560_p3);

assign select_ln20_5_fu_729_p3 = ((icmp_ln20_reg_985[0:0] == 1'b1) ? 6'd1 : add_ln20_1_reg_1028);

assign select_ln20_fu_589_p3 = ((or_ln20_fu_584_p2[0:0] == 1'b1) ? 6'd0 : ap_phi_mux_kk_0_i_phi_fu_243_p4);

assign select_ln33_4_fu_845_p3 = ((select_ln20_2_reg_1057_pp0_iter1_reg[0:0] == 1'b1) ? 16'd0 : bitcast_ln32_4_fu_841_p1);

assign select_ln33_5_fu_867_p3 = ((select_ln20_2_reg_1057_pp0_iter1_reg[0:0] == 1'b1) ? 16'd0 : bitcast_ln32_5_fu_863_p1);

assign select_ln33_6_fu_888_p3 = ((select_ln20_2_reg_1057_pp0_iter1_reg[0:0] == 1'b1) ? 16'd0 : bitcast_ln32_6_fu_884_p1);

assign select_ln33_fu_806_p3 = ((select_ln20_2_reg_1057_pp0_iter1_reg[0:0] == 1'b1) ? 16'd0 : bitcast_ln32_fu_802_p1);

assign sext_ln20_fu_680_p1 = (sub_ln32_fu_674_p2);

assign sext_ln22_fu_282_p1 = add_ln22_fu_276_p2;

assign sext_ln32_fu_724_p1 = (tmp_5_fu_716_p3);

assign sext_ln33_1_fu_907_p1 = (tmp_7_fu_900_p3);

assign sext_ln33_2_fu_924_p1 = (tmp_8_fu_917_p3);

assign sext_ln33_fu_826_p1 = (tmp_6_fu_819_p3);

assign sub_ln32_fu_674_p2 = (zext_ln32_fu_658_p1 - zext_ln32_7_fu_670_p1);

assign sub_ln33_cast_fu_760_p1 = (sub_ln33_fu_754_p2);

assign sub_ln33_fu_754_p2 = (zext_ln33_2_fu_750_p1 - zext_ln33_fu_740_p1);

assign tmp2_cast_fu_509_p1 = (tmp2_fu_503_p2);

assign tmp2_cast_mid1_fu_626_p1 = (tmp2_mid1_fu_620_p2);

assign tmp2_fu_503_p2 = ((zext_ln22_fu_493_p1) + (3'd7));

assign tmp2_mid1_fu_620_p2 = ((zext_ln22_1_fu_603_p1) + (3'd7));

assign tmp_12_i_fu_831_p4 = {{in_data_q0[31:16]}};

assign tmp_13_cast_fu_777_p3 = {{trunc_ln33_fu_773_p1}, {5'd0}};

assign tmp_13_i_fu_853_p4 = {{in_data_q0[47:32]}};

assign tmp_14_i_fu_874_p4 = {{in_data_q0[63:48]}};

assign tmp_1_fu_650_p3 = {{select_ln20_3_fu_642_p3}, {5'd0}};

assign tmp_2_fu_662_p3 = {{select_ln20_3_fu_642_p3}, {2'd0}};

assign tmp_3_fu_351_p3 = add_ln22_1_fu_346_p2[32'd17];

assign tmp_4_fu_455_p3 = add_ln22_2_fu_450_p2[32'd17];

assign tmp_5_fu_716_p3 = {{add_ln32_fu_696_p2}, {lshr_ln_fu_706_p4}};

assign tmp_6_fu_819_p3 = {{add_ln33_reg_1087}, {or_ln25_fu_814_p2}};

assign tmp_7_fu_900_p3 = {{add_ln33_reg_1087}, {or_ln25_3_fu_895_p2}};

assign tmp_8_fu_917_p3 = {{add_ln33_reg_1087}, {or_ln25_4_fu_912_p2}};

assign tmp_fu_292_p3 = add_ln22_fu_276_p2[32'd16];

assign tmp_s_fu_743_p3 = {{select_ln19_1_reg_1038}, {2'd0}};

assign trunc_ln22_fu_272_p1 = j_13[9:0];

assign trunc_ln32_fu_798_p1 = in_data_q0[15:0];

assign trunc_ln33_fu_773_p1 = add_ln33_fu_767_p2[3:0];

assign xor_ln19_fu_567_p2 = (icmp_ln20_reg_985 ^ 1'd1);

assign zext_ln19_fu_254_p1 = i_13;

assign zext_ln20_1_fu_446_p1 = add_ln20_fu_440_p2;

assign zext_ln20_fu_342_p1 = ap_phi_mux_jj_phi_fu_231_p4;

assign zext_ln22_1_fu_603_p1 = add_ln20_reg_1015;

assign zext_ln22_fu_493_p1 = jj_reg_227;

assign zext_ln32_7_fu_670_p1 = tmp_2_fu_662_p3;

assign zext_ln32_8_fu_692_p1 = select_ln20_4_fu_684_p3;

assign zext_ln32_fu_658_p1 = tmp_1_fu_650_p3;

assign zext_ln33_2_fu_750_p1 = tmp_s_fu_743_p3;

assign zext_ln33_3_fu_764_p1 = select_ln20_1_reg_1051;

assign zext_ln33_4_fu_785_p1 = select_ln20_reg_1045;

assign zext_ln33_5_fu_794_p1 = add_ln33_1_reg_1094;

assign zext_ln33_fu_740_p1 = select_ln19_1_reg_1038;

endmodule //td_fused_top_tdf8_readInputs57
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf8_writeOutputs_unaligned (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        i,
        j,
        out_data_address1,
        out_data_ce1,
        out_data_we1,
        out_data_d1,
        max_vals_0
);

parameter    ap_ST_fsm_state1 = 2'd1;
parameter    ap_ST_fsm_state2 = 2'd2;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
input  [3:0] i;
input  [7:0] j;
output  [13:0] out_data_address1;
output   out_data_ce1;
output   out_data_we1;
output  [63:0] out_data_d1;
input  [15:0] max_vals_0;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg out_data_ce1;
reg out_data_we1;

  reg   [1:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg   [15:0] outputCount_3;
reg   [15:0] outputChanIdx_3;
reg   [15:0] outputRow_13_0;
reg   [15:0] outputRow_13_1;
reg   [15:0] outputRow_13_2;
reg   [15:0] outputRow_13_3;
wire   [15:0] add_ln87_fu_177_p2;
wire   [0:0] icmp_ln88_fu_183_p2;
reg   [0:0] icmp_ln88_reg_297;
reg   [15:0] ap_phi_mux_empty_phi_fu_94_p4;
reg   [15:0] empty_reg_91;
wire    ap_CS_fsm_state2;
wire   [63:0] zext_ln94_4_fu_211_p1;
wire   [15:0] select_ln97_fu_269_p3;
wire   [1:0] trunc_ln86_fu_149_p1;
reg   [15:0] ap_sig_allocacmp_outputRow_13_0_load;
reg   [15:0] ap_sig_allocacmp_outputRow_13_1_load;
reg   [15:0] ap_sig_allocacmp_outputRow_13_2_load;
reg   [15:0] ap_sig_allocacmp_outputRow_13_3_load;
wire   [4:0] tmp_8_fu_109_p3;
wire   [7:0] tmp_fu_101_p3;
wire   [7:0] zext_ln94_fu_117_p1;
wire   [7:0] sub_ln94_fu_121_p2;
wire   [7:0] add_ln94_fu_127_p2;
wire   [7:0] trunc_ln94_fu_197_p1;
wire   [13:0] tmp_10_cast_fu_133_p3;
wire   [13:0] zext_ln94_3_fu_201_p1;
wire   [13:0] add_ln94_2_fu_205_p2;
wire   [15:0] bitcast_ln94_6_fu_240_p1;
wire   [15:0] bitcast_ln94_5_fu_232_p1;
wire   [15:0] bitcast_ln94_4_fu_224_p1;
wire   [15:0] bitcast_ln94_fu_216_p1;
wire   [15:0] add_ln96_fu_257_p2;
wire   [0:0] icmp_ln97_fu_263_p2;
reg   [1:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_CS_fsm = 2'd1;
#0 outputCount_3 = 16'd0;
#0 outputChanIdx_3 = 16'd0;
#0 outputRow_13_0 = 16'd0;
#0 outputRow_13_1 = 16'd0;
#0 outputRow_13_2 = 16'd0;
#0 outputRow_13_3 = 16'd0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln88_reg_297 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        empty_reg_91 <= 16'd0;
    end else if (((ap_start == 1'b1) & (icmp_ln88_fu_183_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state1))) begin
        empty_reg_91 <= add_ln87_fu_177_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state1)) begin
        icmp_ln88_reg_297 <= icmp_ln88_fu_183_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_start == 1'b1) & (icmp_ln88_fu_183_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1))) begin
        outputChanIdx_3 <= select_ln97_fu_269_p3;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        outputCount_3 <= ap_phi_mux_empty_phi_fu_94_p4;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_start == 1'b1) & (trunc_ln86_fu_149_p1 == 2'd0) & (1'b1 == ap_CS_fsm_state1))) begin
        outputRow_13_0 <= max_vals_0;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_start == 1'b1) & (trunc_ln86_fu_149_p1 == 2'd1) & (1'b1 == ap_CS_fsm_state1))) begin
        outputRow_13_1 <= max_vals_0;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_start == 1'b1) & (trunc_ln86_fu_149_p1 == 2'd2) & (1'b1 == ap_CS_fsm_state1))) begin
        outputRow_13_2 <= max_vals_0;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_start == 1'b1) & (trunc_ln86_fu_149_p1 == 2'd3) & (1'b1 == ap_CS_fsm_state1))) begin
        outputRow_13_3 <= max_vals_0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state2) | ((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1)))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = 1'b0;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln88_reg_297 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        ap_phi_mux_empty_phi_fu_94_p4 = 16'd0;
    end else begin
        ap_phi_mux_empty_phi_fu_94_p4 = empty_reg_91;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((trunc_ln86_fu_149_p1 == 2'd0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_sig_allocacmp_outputRow_13_0_load = max_vals_0;
    end else begin
        ap_sig_allocacmp_outputRow_13_0_load = outputRow_13_0;
    end
end

always @ (*) begin
    if (((trunc_ln86_fu_149_p1 == 2'd1) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_sig_allocacmp_outputRow_13_1_load = max_vals_0;
    end else begin
        ap_sig_allocacmp_outputRow_13_1_load = outputRow_13_1;
    end
end

always @ (*) begin
    if (((trunc_ln86_fu_149_p1 == 2'd2) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_sig_allocacmp_outputRow_13_2_load = max_vals_0;
    end else begin
        ap_sig_allocacmp_outputRow_13_2_load = outputRow_13_2;
    end
end

always @ (*) begin
    if (((trunc_ln86_fu_149_p1 == 2'd3) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_sig_allocacmp_outputRow_13_3_load = max_vals_0;
    end else begin
        ap_sig_allocacmp_outputRow_13_3_load = outputRow_13_3;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state2) | ((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)))) begin
        out_data_ce1 = 1'b1;
    end else begin
        out_data_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_start == 1'b1) & (icmp_ln88_fu_183_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1))) begin
        out_data_we1 = 1'b1;
    end else begin
        out_data_we1 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_state2 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln87_fu_177_p2 = (outputCount_3 + 16'd1);

assign add_ln94_2_fu_205_p2 = (tmp_10_cast_fu_133_p3 + zext_ln94_3_fu_201_p1);

assign add_ln94_fu_127_p2 = (sub_ln94_fu_121_p2 + j);

assign add_ln96_fu_257_p2 = (outputChanIdx_3 + 16'd1);

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign bitcast_ln94_4_fu_224_p1 = ap_sig_allocacmp_outputRow_13_1_load;

assign bitcast_ln94_5_fu_232_p1 = ap_sig_allocacmp_outputRow_13_2_load;

assign bitcast_ln94_6_fu_240_p1 = ap_sig_allocacmp_outputRow_13_3_load;

assign bitcast_ln94_fu_216_p1 = ap_sig_allocacmp_outputRow_13_0_load;

assign icmp_ln88_fu_183_p2 = ((add_ln87_fu_177_p2 == 16'd4) ? 1'b1 : 1'b0);

assign icmp_ln97_fu_263_p2 = ((add_ln96_fu_257_p2 == 16'd64) ? 1'b1 : 1'b0);

assign out_data_address1 = zext_ln94_4_fu_211_p1;

assign out_data_d1 = {{{{bitcast_ln94_6_fu_240_p1}, {bitcast_ln94_5_fu_232_p1}}, {bitcast_ln94_4_fu_224_p1}}, {bitcast_ln94_fu_216_p1}};

assign select_ln97_fu_269_p3 = ((icmp_ln97_fu_263_p2[0:0] == 1'b1) ? 16'd0 : add_ln96_fu_257_p2);

assign sub_ln94_fu_121_p2 = (tmp_fu_101_p3 - zext_ln94_fu_117_p1);

assign tmp_10_cast_fu_133_p3 = {{add_ln94_fu_127_p2}, {6'd0}};

assign tmp_8_fu_109_p3 = {{i}, {1'd0}};

assign tmp_fu_101_p3 = {{i}, {4'd0}};

assign trunc_ln86_fu_149_p1 = outputCount_3[1:0];

assign trunc_ln94_fu_197_p1 = outputChanIdx_3[7:0];

assign zext_ln94_3_fu_201_p1 = trunc_ln94_fu_197_p1;

assign zext_ln94_4_fu_211_p1 = add_ln94_2_fu_205_p2;

assign zext_ln94_fu_117_p1 = tmp_8_fu_109_p3;

endmodule //td_fused_top_tdf8_writeOutputs_unaligned
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf9_16 (
        in_data_address0,
        in_data_ce0,
        in_data_d0,
        in_data_q0,
        in_data_we0,
        in_data_address1,
        in_data_ce1,
        in_data_d1,
        in_data_q1,
        in_data_we1,
        out_data_address0,
        out_data_ce0,
        out_data_d0,
        out_data_q0,
        out_data_we0,
        out_data_address1,
        out_data_ce1,
        out_data_d1,
        out_data_q1,
        out_data_we1,
        filter_data_address0,
        filter_data_ce0,
        filter_data_d0,
        filter_data_q0,
        filter_data_we0,
        filter_data_address1,
        filter_data_ce1,
        filter_data_d1,
        filter_data_q1,
        filter_data_we1,
        adjustments_address0,
        adjustments_ce0,
        adjustments_d0,
        adjustments_q0,
        adjustments_we0,
        adjustments_address1,
        adjustments_ce1,
        adjustments_d1,
        adjustments_q1,
        adjustments_we1,
        ap_clk,
        ap_rst,
        in_data_empty_n,
        in_data_read,
        out_data_full_n,
        out_data_write,
        ap_start,
        ap_done,
        ap_ready,
        ap_idle,
        ap_continue
);


output  [13:0] in_data_address0;
output   in_data_ce0;
output  [63:0] in_data_d0;
input  [63:0] in_data_q0;
output   in_data_we0;
output  [13:0] in_data_address1;
output   in_data_ce1;
output  [63:0] in_data_d1;
input  [63:0] in_data_q1;
output   in_data_we1;
output  [11:0] out_data_address0;
output   out_data_ce0;
output  [63:0] out_data_d0;
input  [63:0] out_data_q0;
output   out_data_we0;
output  [11:0] out_data_address1;
output   out_data_ce1;
output  [63:0] out_data_d1;
input  [63:0] out_data_q1;
output   out_data_we1;
output  [13:0] filter_data_address0;
output   filter_data_ce0;
output  [15:0] filter_data_d0;
input  [15:0] filter_data_q0;
output   filter_data_we0;
output  [13:0] filter_data_address1;
output   filter_data_ce1;
output  [15:0] filter_data_d1;
input  [15:0] filter_data_q1;
output   filter_data_we1;
output  [5:0] adjustments_address0;
output   adjustments_ce0;
output  [47:0] adjustments_d0;
input  [47:0] adjustments_q0;
output   adjustments_we0;
output  [5:0] adjustments_address1;
output   adjustments_ce1;
output  [47:0] adjustments_d1;
input  [47:0] adjustments_q1;
output   adjustments_we1;
input   ap_clk;
input   ap_rst;
input   in_data_empty_n;
output   in_data_read;
input   out_data_full_n;
output   out_data_write;
input   ap_start;
output   ap_done;
output   ap_ready;
output   ap_idle;
input   ap_continue;

reg ap_done;
reg ap_ready;
reg ap_idle;

wire   [13:0] dataflow_in_loop_TOP_LOOP37360_U0_in_data_address0;
wire    dataflow_in_loop_TOP_LOOP37360_U0_in_data_ce0;
wire   [63:0] dataflow_in_loop_TOP_LOOP37360_U0_in_data_d0;
wire    dataflow_in_loop_TOP_LOOP37360_U0_in_data_we0;
wire   [13:0] dataflow_in_loop_TOP_LOOP37360_U0_in_data_address1;
wire    dataflow_in_loop_TOP_LOOP37360_U0_in_data_ce1;
wire   [63:0] dataflow_in_loop_TOP_LOOP37360_U0_in_data_d1;
wire    dataflow_in_loop_TOP_LOOP37360_U0_in_data_we1;
wire   [13:0] dataflow_in_loop_TOP_LOOP37360_U0_filter_data_address0;
wire    dataflow_in_loop_TOP_LOOP37360_U0_filter_data_ce0;
wire   [15:0] dataflow_in_loop_TOP_LOOP37360_U0_filter_data_d0;
wire    dataflow_in_loop_TOP_LOOP37360_U0_filter_data_we0;
wire   [13:0] dataflow_in_loop_TOP_LOOP37360_U0_filter_data_address1;
wire    dataflow_in_loop_TOP_LOOP37360_U0_filter_data_ce1;
wire   [15:0] dataflow_in_loop_TOP_LOOP37360_U0_filter_data_d1;
wire    dataflow_in_loop_TOP_LOOP37360_U0_filter_data_we1;
wire   [5:0] dataflow_in_loop_TOP_LOOP37360_U0_adjustments_address0;
wire    dataflow_in_loop_TOP_LOOP37360_U0_adjustments_ce0;
wire   [47:0] dataflow_in_loop_TOP_LOOP37360_U0_adjustments_d0;
wire    dataflow_in_loop_TOP_LOOP37360_U0_adjustments_we0;
wire   [5:0] dataflow_in_loop_TOP_LOOP37360_U0_adjustments_address1;
wire    dataflow_in_loop_TOP_LOOP37360_U0_adjustments_ce1;
wire   [47:0] dataflow_in_loop_TOP_LOOP37360_U0_adjustments_d1;
wire    dataflow_in_loop_TOP_LOOP37360_U0_adjustments_we1;
wire   [11:0] dataflow_in_loop_TOP_LOOP37360_U0_out_data_address0;
wire    dataflow_in_loop_TOP_LOOP37360_U0_out_data_ce0;
wire   [63:0] dataflow_in_loop_TOP_LOOP37360_U0_out_data_d0;
wire    dataflow_in_loop_TOP_LOOP37360_U0_out_data_we0;
wire   [11:0] dataflow_in_loop_TOP_LOOP37360_U0_out_data_address1;
wire    dataflow_in_loop_TOP_LOOP37360_U0_out_data_ce1;
wire   [63:0] dataflow_in_loop_TOP_LOOP37360_U0_out_data_d1;
wire    dataflow_in_loop_TOP_LOOP37360_U0_out_data_we1;
wire    dataflow_in_loop_TOP_LOOP37360_U0_ap_start;
wire    dataflow_in_loop_TOP_LOOP37360_U0_in_data_read;
wire    dataflow_in_loop_TOP_LOOP37360_U0_out_data_write;
wire    dataflow_in_loop_TOP_LOOP37360_U0_ap_done;
wire    dataflow_in_loop_TOP_LOOP37360_U0_ap_ready;
wire    dataflow_in_loop_TOP_LOOP37360_U0_ap_idle;
reg    dataflow_in_loop_TOP_LOOP37360_U0_ap_continue;
wire    dataflow_in_loop_TOP_LOOP37360_U0_in_data_full_n;
wire    dataflow_in_loop_TOP_LOOP37360_U0_in_data_write;
wire    ap_sync_continue;
wire    ap_sync_done;
wire    ap_sync_ready;
reg   [13:0] loop_dataflow_input_count;
reg   [13:0] loop_dataflow_output_count;
wire   [13:0] bound_minus_1;
wire    dataflow_in_loop_TOP_LOOP37360_U0_start_full_n;
wire    dataflow_in_loop_TOP_LOOP37360_U0_start_write;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 loop_dataflow_input_count = 14'd0;
#0 loop_dataflow_output_count = 14'd0;
end

td_fused_top_dataflow_in_loop_TOP_LOOP37360 dataflow_in_loop_TOP_LOOP37360_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .in_data_address0(dataflow_in_loop_TOP_LOOP37360_U0_in_data_address0),
    .in_data_ce0(dataflow_in_loop_TOP_LOOP37360_U0_in_data_ce0),
    .in_data_d0(dataflow_in_loop_TOP_LOOP37360_U0_in_data_d0),
    .in_data_q0(in_data_q0),
    .in_data_we0(dataflow_in_loop_TOP_LOOP37360_U0_in_data_we0),
    .in_data_address1(dataflow_in_loop_TOP_LOOP37360_U0_in_data_address1),
    .in_data_ce1(dataflow_in_loop_TOP_LOOP37360_U0_in_data_ce1),
    .in_data_d1(dataflow_in_loop_TOP_LOOP37360_U0_in_data_d1),
    .in_data_q1(64'd0),
    .in_data_we1(dataflow_in_loop_TOP_LOOP37360_U0_in_data_we1),
    .filter_data_address0(dataflow_in_loop_TOP_LOOP37360_U0_filter_data_address0),
    .filter_data_ce0(dataflow_in_loop_TOP_LOOP37360_U0_filter_data_ce0),
    .filter_data_d0(dataflow_in_loop_TOP_LOOP37360_U0_filter_data_d0),
    .filter_data_q0(filter_data_q0),
    .filter_data_we0(dataflow_in_loop_TOP_LOOP37360_U0_filter_data_we0),
    .filter_data_address1(dataflow_in_loop_TOP_LOOP37360_U0_filter_data_address1),
    .filter_data_ce1(dataflow_in_loop_TOP_LOOP37360_U0_filter_data_ce1),
    .filter_data_d1(dataflow_in_loop_TOP_LOOP37360_U0_filter_data_d1),
    .filter_data_q1(16'd0),
    .filter_data_we1(dataflow_in_loop_TOP_LOOP37360_U0_filter_data_we1),
    .adjustments_address0(dataflow_in_loop_TOP_LOOP37360_U0_adjustments_address0),
    .adjustments_ce0(dataflow_in_loop_TOP_LOOP37360_U0_adjustments_ce0),
    .adjustments_d0(dataflow_in_loop_TOP_LOOP37360_U0_adjustments_d0),
    .adjustments_q0(adjustments_q0),
    .adjustments_we0(dataflow_in_loop_TOP_LOOP37360_U0_adjustments_we0),
    .adjustments_address1(dataflow_in_loop_TOP_LOOP37360_U0_adjustments_address1),
    .adjustments_ce1(dataflow_in_loop_TOP_LOOP37360_U0_adjustments_ce1),
    .adjustments_d1(dataflow_in_loop_TOP_LOOP37360_U0_adjustments_d1),
    .adjustments_q1(48'd0),
    .adjustments_we1(dataflow_in_loop_TOP_LOOP37360_U0_adjustments_we1),
    .out_data_address0(dataflow_in_loop_TOP_LOOP37360_U0_out_data_address0),
    .out_data_ce0(dataflow_in_loop_TOP_LOOP37360_U0_out_data_ce0),
    .out_data_d0(dataflow_in_loop_TOP_LOOP37360_U0_out_data_d0),
    .out_data_q0(64'd0),
    .out_data_we0(dataflow_in_loop_TOP_LOOP37360_U0_out_data_we0),
    .out_data_address1(dataflow_in_loop_TOP_LOOP37360_U0_out_data_address1),
    .out_data_ce1(dataflow_in_loop_TOP_LOOP37360_U0_out_data_ce1),
    .out_data_d1(dataflow_in_loop_TOP_LOOP37360_U0_out_data_d1),
    .out_data_q1(64'd0),
    .out_data_we1(dataflow_in_loop_TOP_LOOP37360_U0_out_data_we1),
    .ap_start(dataflow_in_loop_TOP_LOOP37360_U0_ap_start),
    .in_data_empty_n(1'b0),
    .in_data_read(dataflow_in_loop_TOP_LOOP37360_U0_in_data_read),
    .out_data_full_n(out_data_full_n),
    .out_data_write(dataflow_in_loop_TOP_LOOP37360_U0_out_data_write),
    .ap_done(dataflow_in_loop_TOP_LOOP37360_U0_ap_done),
    .ap_ready(dataflow_in_loop_TOP_LOOP37360_U0_ap_ready),
    .ap_idle(dataflow_in_loop_TOP_LOOP37360_U0_ap_idle),
    .ap_continue(dataflow_in_loop_TOP_LOOP37360_U0_ap_continue)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        loop_dataflow_input_count <= 14'd0;
    end else begin
        if ((~(loop_dataflow_input_count == bound_minus_1) & (dataflow_in_loop_TOP_LOOP37360_U0_ap_ready == 1'b1) & (ap_start == 1'b1))) begin
            loop_dataflow_input_count <= (loop_dataflow_input_count + 14'd1);
        end else if (((dataflow_in_loop_TOP_LOOP37360_U0_ap_ready == 1'b1) & (loop_dataflow_input_count == bound_minus_1) & (ap_start == 1'b1))) begin
            loop_dataflow_input_count <= 14'd0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        loop_dataflow_output_count <= 14'd0;
    end else begin
        if ((~(loop_dataflow_output_count == bound_minus_1) & (dataflow_in_loop_TOP_LOOP37360_U0_ap_continue == 1'b1) & (dataflow_in_loop_TOP_LOOP37360_U0_ap_done == 1'b1))) begin
            loop_dataflow_output_count <= (loop_dataflow_output_count + 14'd1);
        end else if (((dataflow_in_loop_TOP_LOOP37360_U0_ap_continue == 1'b1) & (dataflow_in_loop_TOP_LOOP37360_U0_ap_done == 1'b1) & (loop_dataflow_output_count == bound_minus_1))) begin
            loop_dataflow_output_count <= 14'd0;
        end
    end
end

always @ (*) begin
    if (((dataflow_in_loop_TOP_LOOP37360_U0_ap_done == 1'b1) & (loop_dataflow_output_count == bound_minus_1))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = 1'b0;
    end
end

always @ (*) begin
    if (((dataflow_in_loop_TOP_LOOP37360_U0_ap_idle == 1'b1) & (loop_dataflow_output_count == 14'd0) & (ap_start == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((dataflow_in_loop_TOP_LOOP37360_U0_ap_ready == 1'b1) & (loop_dataflow_input_count == bound_minus_1) & (ap_start == 1'b1))) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((~(loop_dataflow_output_count == bound_minus_1) | (ap_continue == 1'b1))) begin
        dataflow_in_loop_TOP_LOOP37360_U0_ap_continue = 1'b1;
    end else begin
        dataflow_in_loop_TOP_LOOP37360_U0_ap_continue = 1'b0;
    end
end

assign adjustments_address0 = dataflow_in_loop_TOP_LOOP37360_U0_adjustments_address0;

assign adjustments_address1 = 6'd0;

assign adjustments_ce0 = dataflow_in_loop_TOP_LOOP37360_U0_adjustments_ce0;

assign adjustments_ce1 = 1'b0;

assign adjustments_d0 = 48'd0;

assign adjustments_d1 = 48'd0;

assign adjustments_we0 = 1'b0;

assign adjustments_we1 = 1'b0;

assign ap_sync_continue = ap_continue;

assign ap_sync_done = dataflow_in_loop_TOP_LOOP37360_U0_ap_done;

assign ap_sync_ready = dataflow_in_loop_TOP_LOOP37360_U0_ap_ready;

assign bound_minus_1 = (14'd12544 - 14'd1);

assign dataflow_in_loop_TOP_LOOP37360_U0_ap_start = ap_start;

assign dataflow_in_loop_TOP_LOOP37360_U0_in_data_full_n = in_data_empty_n;

assign dataflow_in_loop_TOP_LOOP37360_U0_in_data_write = 1'b0;

assign dataflow_in_loop_TOP_LOOP37360_U0_start_full_n = 1'b1;

assign dataflow_in_loop_TOP_LOOP37360_U0_start_write = 1'b0;

assign filter_data_address0 = dataflow_in_loop_TOP_LOOP37360_U0_filter_data_address0;

assign filter_data_address1 = 14'd0;

assign filter_data_ce0 = dataflow_in_loop_TOP_LOOP37360_U0_filter_data_ce0;

assign filter_data_ce1 = 1'b0;

assign filter_data_d0 = 16'd0;

assign filter_data_d1 = 16'd0;

assign filter_data_we0 = 1'b0;

assign filter_data_we1 = 1'b0;

assign in_data_address0 = dataflow_in_loop_TOP_LOOP37360_U0_in_data_address0;

assign in_data_address1 = 14'd0;

assign in_data_ce0 = dataflow_in_loop_TOP_LOOP37360_U0_in_data_ce0;

assign in_data_ce1 = 1'b0;

assign in_data_d0 = 64'd0;

assign in_data_d1 = 64'd0;

assign in_data_read = dataflow_in_loop_TOP_LOOP37360_U0_in_data_write;

assign in_data_we0 = 1'b0;

assign in_data_we1 = 1'b0;

assign out_data_address0 = 12'd0;

assign out_data_address1 = dataflow_in_loop_TOP_LOOP37360_U0_out_data_address1;

assign out_data_ce0 = 1'b0;

assign out_data_ce1 = dataflow_in_loop_TOP_LOOP37360_U0_out_data_ce1;

assign out_data_d0 = 64'd0;

assign out_data_d1 = dataflow_in_loop_TOP_LOOP37360_U0_out_data_d1;

assign out_data_we0 = 1'b0;

assign out_data_we1 = dataflow_in_loop_TOP_LOOP37360_U0_out_data_we1;

assign out_data_write = dataflow_in_loop_TOP_LOOP37360_U0_out_data_write;

endmodule //td_fused_top_tdf9_16
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf9_accum_1 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        accum_in_0_address0,
        accum_in_0_ce0,
        accum_in_0_q0,
        accum_in_0_address1,
        accum_in_0_ce1,
        accum_in_0_q1,
        accum_out_address0,
        accum_out_ce0,
        accum_out_we0,
        accum_out_d0,
        accum_out_address1,
        accum_out_ce1,
        accum_out_we1,
        accum_out_d1
);

parameter    ap_ST_fsm_state1 = 8'd1;
parameter    ap_ST_fsm_pp0_stage0 = 8'd2;
parameter    ap_ST_fsm_pp0_stage1 = 8'd4;
parameter    ap_ST_fsm_pp0_stage2 = 8'd8;
parameter    ap_ST_fsm_pp0_stage3 = 8'd16;
parameter    ap_ST_fsm_state12 = 8'd32;
parameter    ap_ST_fsm_state13 = 8'd64;
parameter    ap_ST_fsm_state14 = 8'd128;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [7:0] accum_in_0_address0;
output   accum_in_0_ce0;
input  [15:0] accum_in_0_q0;
output  [7:0] accum_in_0_address1;
output   accum_in_0_ce1;
input  [15:0] accum_in_0_q1;
output  [2:0] accum_out_address0;
output   accum_out_ce0;
output   accum_out_we0;
output  [15:0] accum_out_d0;
output  [2:0] accum_out_address1;
output   accum_out_ce1;
output   accum_out_we1;
output  [15:0] accum_out_d1;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg[7:0] accum_in_0_address0;
reg accum_in_0_ce0;
reg[7:0] accum_in_0_address1;
reg accum_in_0_ce1;
reg accum_out_ce0;
reg accum_out_we0;
reg accum_out_ce1;
reg accum_out_we1;

reg    ap_done_reg;
  reg   [7:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg   [8:0] x_reg_170;
reg   [15:0] psum_7_08_reg_182;
reg   [15:0] psum_6_07_reg_194;
reg   [15:0] psum_5_06_reg_206;
reg   [15:0] psum_4_05_reg_218;
reg   [15:0] psum_3_04_reg_230;
reg   [15:0] psum_2_03_reg_242;
reg   [15:0] psum_1_02_reg_254;
reg   [15:0] psum_0_01_reg_266;
wire   [0:0] tmp_fu_323_p3;
reg   [0:0] tmp_reg_494;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state6_pp0_stage0_iter1;
wire    ap_block_state10_pp0_stage0_iter2;
wire    ap_block_pp0_stage0_11001;
reg   [0:0] tmp_reg_494_pp0_iter1_reg;
reg   [0:0] tmp_reg_494_pp0_iter2_reg;
wire   [7:0] trunc_ln25_fu_336_p1;
reg   [7:0] trunc_ln25_reg_498;
reg   [15:0] accum_in_0_load_reg_518;
wire    ap_CS_fsm_pp0_stage1;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_state3_pp0_stage1_iter0;
wire    ap_block_state7_pp0_stage1_iter1;
wire    ap_block_state11_pp0_stage1_iter2;
wire    ap_block_pp0_stage1_11001;
reg   [15:0] accum_in_0_load_1_reg_523;
reg   [15:0] accum_in_0_load_2_reg_538;
wire    ap_CS_fsm_pp0_stage2;
wire    ap_block_state4_pp0_stage2_iter0;
wire    ap_block_state8_pp0_stage2_iter1;
wire    ap_block_pp0_stage2_11001;
reg   [15:0] accum_in_0_load_3_reg_543;
wire   [8:0] add_ln25_fu_391_p2;
reg   [8:0] add_ln25_reg_558;
wire    ap_CS_fsm_pp0_stage3;
wire    ap_block_state5_pp0_stage3_iter0;
wire    ap_block_state9_pp0_stage3_iter1;
wire    ap_block_pp0_stage3_11001;
reg   [15:0] accum_in_0_load_4_reg_563;
reg   [15:0] accum_in_0_load_5_reg_568;
reg   [15:0] accum_in_0_load_6_reg_583;
reg    ap_enable_reg_pp0_iter1;
reg   [15:0] accum_in_0_load_7_reg_588;
wire   [15:0] grp_fu_307_p2;
wire   [15:0] grp_fu_312_p2;
reg    ap_enable_reg_pp0_iter2;
wire   [3:0] add_ln33_fu_434_p2;
wire    ap_CS_fsm_state13;
wire   [0:0] tmp_2_fu_417_p3;
reg    ap_block_state1;
wire    ap_block_pp0_stage2_subdone;
reg    ap_condition_pp0_exit_iter0_state4;
wire    ap_block_pp0_stage3_subdone;
wire    ap_block_pp0_stage1_subdone;
reg   [8:0] ap_phi_mux_x_phi_fu_174_p4;
wire    ap_block_pp0_stage0;
wire   [15:0] ap_phi_mux_psum_7_08_phi_fu_186_p4;
wire    ap_block_pp0_stage1;
wire   [15:0] ap_phi_mux_psum_6_07_phi_fu_198_p4;
wire   [15:0] ap_phi_mux_psum_5_06_phi_fu_210_p4;
wire   [15:0] ap_phi_mux_psum_4_05_phi_fu_222_p4;
wire   [15:0] ap_phi_mux_psum_3_04_phi_fu_234_p4;
wire    ap_block_pp0_stage3;
wire   [15:0] ap_phi_mux_psum_2_03_phi_fu_246_p4;
wire    ap_block_pp0_stage2;
reg   [3:0] q_reg_278;
wire    ap_CS_fsm_state12;
reg   [15:0] ap_phi_mux_phi_ln45_phi_fu_292_p8;
wire   [2:0] trunc_ln33_fu_430_p1;
wire   [63:0] zext_ln25_fu_331_p1;
wire   [63:0] zext_ln29_fu_346_p1;
wire   [63:0] zext_ln29_1_fu_356_p1;
wire   [63:0] zext_ln29_2_fu_366_p1;
wire   [63:0] zext_ln29_3_fu_376_p1;
wire   [63:0] zext_ln29_4_fu_386_p1;
wire   [63:0] zext_ln29_5_fu_402_p1;
wire   [63:0] zext_ln29_6_fu_412_p1;
wire   [63:0] zext_ln33_fu_425_p1;
wire   [63:0] zext_ln33_1_fu_446_p1;
reg   [15:0] grp_fu_307_p0;
reg   [15:0] grp_fu_307_p1;
reg   [15:0] grp_fu_312_p0;
reg   [15:0] grp_fu_312_p1;
wire   [7:0] or_ln29_fu_340_p2;
wire   [7:0] or_ln29_1_fu_351_p2;
wire   [7:0] or_ln29_2_fu_361_p2;
wire   [7:0] or_ln29_3_fu_371_p2;
wire   [7:0] or_ln29_4_fu_381_p2;
wire   [7:0] or_ln29_5_fu_397_p2;
wire   [7:0] or_ln29_6_fu_407_p2;
wire   [2:0] or_ln33_fu_440_p2;
wire   [0:0] icmp_ln45_fu_451_p2;
wire   [0:0] icmp_ln45_1_fu_465_p2;
wire   [15:0] select_ln45_fu_457_p3;
wire   [0:0] icmp_ln45_2_fu_479_p2;
wire   [15:0] select_ln45_1_fu_471_p3;
wire    ap_CS_fsm_state14;
reg   [7:0] ap_NS_fsm;
wire    ap_block_pp0_stage0_subdone;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
reg    ap_condition_518;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 8'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
end

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U564(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(grp_fu_307_p0),
    .din1(grp_fu_307_p1),
    .dout(grp_fu_307_p2)
);

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U565(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(grp_fu_312_p0),
    .din1(grp_fu_312_p1),
    .dout(grp_fu_312_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state14)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage2_subdone) & (1'b1 == ap_condition_pp0_exit_iter0_state4) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage3_subdone) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b0)) | ((1'b0 == ap_block_pp0_stage3_subdone) & (1'b1 == ap_CS_fsm_pp0_stage3)))) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end else if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter2 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state12)) begin
        q_reg_278 <= 4'd0;
    end else if (((tmp_2_fu_417_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state13))) begin
        q_reg_278 <= add_ln33_fu_434_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (tmp_reg_494 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        x_reg_170 <= add_ln25_reg_558;
    end else if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        x_reg_170 <= 9'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage1_11001) & (tmp_reg_494 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
        accum_in_0_load_1_reg_523 <= accum_in_0_q0;
        accum_in_0_load_reg_518 <= accum_in_0_q1;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage2_11001) & (tmp_reg_494 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage2) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
        accum_in_0_load_2_reg_538 <= accum_in_0_q1;
        accum_in_0_load_3_reg_543 <= accum_in_0_q0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage3_11001) & (tmp_reg_494 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage3) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
        accum_in_0_load_4_reg_563 <= accum_in_0_q1;
        accum_in_0_load_5_reg_568 <= accum_in_0_q0;
        add_ln25_reg_558 <= add_ln25_fu_391_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (tmp_reg_494 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        accum_in_0_load_6_reg_583 <= accum_in_0_q1;
        accum_in_0_load_7_reg_588 <= accum_in_0_q0;
    end
end

always @ (posedge ap_clk) begin
    if (((tmp_reg_494_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage2_11001) & (1'b1 == ap_CS_fsm_pp0_stage2) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        psum_0_01_reg_266 <= grp_fu_307_p2;
        psum_1_02_reg_254 <= grp_fu_312_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((tmp_reg_494_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage3_11001) & (1'b1 == ap_CS_fsm_pp0_stage3) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        psum_2_03_reg_242 <= grp_fu_307_p2;
        psum_3_04_reg_230 <= grp_fu_312_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((tmp_reg_494_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        psum_4_05_reg_218 <= grp_fu_307_p2;
        psum_5_06_reg_206 <= grp_fu_312_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((tmp_reg_494_pp0_iter2_reg == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
        psum_6_07_reg_194 <= grp_fu_307_p2;
        psum_7_08_reg_182 <= grp_fu_312_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_reg_494 <= ap_phi_mux_x_phi_fu_174_p4[32'd8];
        tmp_reg_494_pp0_iter1_reg <= tmp_reg_494;
        tmp_reg_494_pp0_iter2_reg <= tmp_reg_494_pp0_iter1_reg;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (tmp_fu_323_p3 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        trunc_ln25_reg_498 <= trunc_ln25_fu_336_p1;
    end
end

always @ (*) begin
    if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
        if (((1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            accum_in_0_address0 = zext_ln29_6_fu_412_p1;
        end else if (((1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            accum_in_0_address0 = zext_ln29_4_fu_386_p1;
        end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            accum_in_0_address0 = zext_ln29_2_fu_366_p1;
        end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            accum_in_0_address0 = zext_ln29_fu_346_p1;
        end else begin
            accum_in_0_address0 = 'bx;
        end
    end else begin
        accum_in_0_address0 = 'bx;
    end
end

always @ (*) begin
    if ((ap_enable_reg_pp0_iter0 == 1'b1)) begin
        if (((1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            accum_in_0_address1 = zext_ln29_5_fu_402_p1;
        end else if (((1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            accum_in_0_address1 = zext_ln29_3_fu_376_p1;
        end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            accum_in_0_address1 = zext_ln29_1_fu_356_p1;
        end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            accum_in_0_address1 = zext_ln25_fu_331_p1;
        end else begin
            accum_in_0_address1 = 'bx;
        end
    end else begin
        accum_in_0_address1 = 'bx;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1)) | ((1'b0 == ap_block_pp0_stage3_11001) & (1'b1 == ap_CS_fsm_pp0_stage3) & (ap_enable_reg_pp0_iter0 == 1'b1)) | ((1'b0 == ap_block_pp0_stage2_11001) & (1'b1 == ap_CS_fsm_pp0_stage2) & (ap_enable_reg_pp0_iter0 == 1'b1)) | ((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1)))) begin
        accum_in_0_ce0 = 1'b1;
    end else begin
        accum_in_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1)) | ((1'b0 == ap_block_pp0_stage3_11001) & (1'b1 == ap_CS_fsm_pp0_stage3) & (ap_enable_reg_pp0_iter0 == 1'b1)) | ((1'b0 == ap_block_pp0_stage2_11001) & (1'b1 == ap_CS_fsm_pp0_stage2) & (ap_enable_reg_pp0_iter0 == 1'b1)) | ((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1)))) begin
        accum_in_0_ce1 = 1'b1;
    end else begin
        accum_in_0_ce1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state13)) begin
        accum_out_ce0 = 1'b1;
    end else begin
        accum_out_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state13)) begin
        accum_out_ce1 = 1'b1;
    end else begin
        accum_out_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((tmp_2_fu_417_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state13))) begin
        accum_out_we0 = 1'b1;
    end else begin
        accum_out_we0 = 1'b0;
    end
end

always @ (*) begin
    if (((tmp_2_fu_417_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state13))) begin
        accum_out_we1 = 1'b1;
    end else begin
        accum_out_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((tmp_reg_494 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state4 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state4 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state14)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((tmp_2_fu_417_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state13))) begin
        if ((trunc_ln33_fu_430_p1 == 3'd0)) begin
            ap_phi_mux_phi_ln45_phi_fu_292_p8 = psum_0_01_reg_266;
        end else if ((1'b1 == ap_condition_518)) begin
            ap_phi_mux_phi_ln45_phi_fu_292_p8 = psum_6_07_reg_194;
        end else if ((trunc_ln33_fu_430_p1 == 3'd4)) begin
            ap_phi_mux_phi_ln45_phi_fu_292_p8 = psum_4_05_reg_218;
        end else if ((trunc_ln33_fu_430_p1 == 3'd2)) begin
            ap_phi_mux_phi_ln45_phi_fu_292_p8 = psum_2_03_reg_242;
        end else begin
            ap_phi_mux_phi_ln45_phi_fu_292_p8 = 'bx;
        end
    end else begin
        ap_phi_mux_phi_ln45_phi_fu_292_p8 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0) & (tmp_reg_494 == 1'd0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_x_phi_fu_174_p4 = add_ln25_reg_558;
    end else begin
        ap_phi_mux_x_phi_fu_174_p4 = x_reg_170;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state14)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_307_p0 = ap_phi_mux_psum_6_07_phi_fu_198_p4;
    end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_307_p0 = ap_phi_mux_psum_4_05_phi_fu_222_p4;
    end else if (((1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
        grp_fu_307_p0 = ap_phi_mux_psum_2_03_phi_fu_246_p4;
    end else if (((1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
        grp_fu_307_p0 = grp_fu_307_p2;
    end else begin
        grp_fu_307_p0 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_307_p1 = accum_in_0_load_6_reg_583;
    end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_307_p1 = accum_in_0_load_4_reg_563;
    end else if (((1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
        grp_fu_307_p1 = accum_in_0_load_2_reg_538;
    end else if (((1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
        grp_fu_307_p1 = accum_in_0_load_reg_518;
    end else begin
        grp_fu_307_p1 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_312_p0 = ap_phi_mux_psum_7_08_phi_fu_186_p4;
    end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_312_p0 = ap_phi_mux_psum_5_06_phi_fu_210_p4;
    end else if (((1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
        grp_fu_312_p0 = ap_phi_mux_psum_3_04_phi_fu_234_p4;
    end else if (((1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
        grp_fu_312_p0 = grp_fu_312_p2;
    end else begin
        grp_fu_312_p0 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_312_p1 = accum_in_0_load_7_reg_588;
    end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        grp_fu_312_p1 = accum_in_0_load_5_reg_568;
    end else if (((1'b0 == ap_block_pp0_stage3) & (1'b1 == ap_CS_fsm_pp0_stage3) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
        grp_fu_312_p1 = accum_in_0_load_3_reg_543;
    end else if (((1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
        grp_fu_312_p1 = accum_in_0_load_1_reg_523;
    end else begin
        grp_fu_312_p1 = 'bx;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_pp0_stage1 : begin
            if ((~((1'b0 == ap_block_pp0_stage1_subdone) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b0)) & (1'b0 == ap_block_pp0_stage1_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage2;
            end else if (((1'b0 == ap_block_pp0_stage1_subdone) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
                ap_NS_fsm = ap_ST_fsm_state12;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end
        end
        ap_ST_fsm_pp0_stage2 : begin
            if ((~((1'b0 == ap_block_pp0_stage2_subdone) & (tmp_reg_494 == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1)) & (1'b0 == ap_block_pp0_stage2_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage3;
            end else if (((1'b0 == ap_block_pp0_stage2_subdone) & (tmp_reg_494 == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
                ap_NS_fsm = ap_ST_fsm_state12;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage2;
            end
        end
        ap_ST_fsm_pp0_stage3 : begin
            if ((1'b0 == ap_block_pp0_stage3_subdone)) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage3;
            end
        end
        ap_ST_fsm_state12 : begin
            ap_NS_fsm = ap_ST_fsm_state13;
        end
        ap_ST_fsm_state13 : begin
            if (((tmp_2_fu_417_p3 == 1'd0) & (1'b1 == ap_CS_fsm_state13))) begin
                ap_NS_fsm = ap_ST_fsm_state13;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state14;
            end
        end
        ap_ST_fsm_state14 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign accum_out_address0 = zext_ln33_1_fu_446_p1;

assign accum_out_address1 = zext_ln33_fu_425_p1;

assign accum_out_d0 = ((icmp_ln45_2_fu_479_p2[0:0] == 1'b1) ? psum_5_06_reg_206 : select_ln45_1_fu_471_p3);

assign accum_out_d1 = ap_phi_mux_phi_ln45_phi_fu_292_p8;

assign add_ln25_fu_391_p2 = (x_reg_170 + 9'd8);

assign add_ln33_fu_434_p2 = (q_reg_278 + 4'd2);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_pp0_stage1 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_pp0_stage2 = ap_CS_fsm[32'd3];

assign ap_CS_fsm_pp0_stage3 = ap_CS_fsm[32'd4];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state12 = ap_CS_fsm[32'd5];

assign ap_CS_fsm_state13 = ap_CS_fsm[32'd6];

assign ap_CS_fsm_state14 = ap_CS_fsm[32'd7];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1_subdone = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage2 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage2_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage2_subdone = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage3 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage3_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage3_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((ap_done_reg == 1'b1) | (ap_start == 1'b0));
end

assign ap_block_state10_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state11_pp0_stage1_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage1_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage2_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage3_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage1_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage2_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state9_pp0_stage3_iter1 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_condition_518 = (~(trunc_ln33_fu_430_p1 == 3'd0) & ~(trunc_ln33_fu_430_p1 == 3'd4) & ~(trunc_ln33_fu_430_p1 == 3'd2));
end

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign ap_phi_mux_psum_2_03_phi_fu_246_p4 = grp_fu_307_p2;

assign ap_phi_mux_psum_3_04_phi_fu_234_p4 = grp_fu_312_p2;

assign ap_phi_mux_psum_4_05_phi_fu_222_p4 = grp_fu_307_p2;

assign ap_phi_mux_psum_5_06_phi_fu_210_p4 = grp_fu_312_p2;

assign ap_phi_mux_psum_6_07_phi_fu_198_p4 = grp_fu_307_p2;

assign ap_phi_mux_psum_7_08_phi_fu_186_p4 = grp_fu_312_p2;

assign icmp_ln45_1_fu_465_p2 = ((or_ln33_fu_440_p2 == 3'd3) ? 1'b1 : 1'b0);

assign icmp_ln45_2_fu_479_p2 = ((or_ln33_fu_440_p2 == 3'd5) ? 1'b1 : 1'b0);

assign icmp_ln45_fu_451_p2 = ((or_ln33_fu_440_p2 == 3'd1) ? 1'b1 : 1'b0);

assign or_ln29_1_fu_351_p2 = (trunc_ln25_reg_498 | 8'd2);

assign or_ln29_2_fu_361_p2 = (trunc_ln25_reg_498 | 8'd3);

assign or_ln29_3_fu_371_p2 = (trunc_ln25_reg_498 | 8'd4);

assign or_ln29_4_fu_381_p2 = (trunc_ln25_reg_498 | 8'd5);

assign or_ln29_5_fu_397_p2 = (trunc_ln25_reg_498 | 8'd6);

assign or_ln29_6_fu_407_p2 = (trunc_ln25_reg_498 | 8'd7);

assign or_ln29_fu_340_p2 = (trunc_ln25_fu_336_p1 | 8'd1);

assign or_ln33_fu_440_p2 = (trunc_ln33_fu_430_p1 | 3'd1);

assign select_ln45_1_fu_471_p3 = ((icmp_ln45_1_fu_465_p2[0:0] == 1'b1) ? psum_3_04_reg_230 : select_ln45_fu_457_p3);

assign select_ln45_fu_457_p3 = ((icmp_ln45_fu_451_p2[0:0] == 1'b1) ? psum_1_02_reg_254 : psum_7_08_reg_182);

assign tmp_2_fu_417_p3 = q_reg_278[32'd3];

assign tmp_fu_323_p3 = ap_phi_mux_x_phi_fu_174_p4[32'd8];

assign trunc_ln25_fu_336_p1 = ap_phi_mux_x_phi_fu_174_p4[7:0];

assign trunc_ln33_fu_430_p1 = q_reg_278[2:0];

assign zext_ln25_fu_331_p1 = ap_phi_mux_x_phi_fu_174_p4;

assign zext_ln29_1_fu_356_p1 = or_ln29_1_fu_351_p2;

assign zext_ln29_2_fu_366_p1 = or_ln29_2_fu_361_p2;

assign zext_ln29_3_fu_376_p1 = or_ln29_3_fu_371_p2;

assign zext_ln29_4_fu_386_p1 = or_ln29_4_fu_381_p2;

assign zext_ln29_5_fu_402_p1 = or_ln29_5_fu_397_p2;

assign zext_ln29_6_fu_412_p1 = or_ln29_6_fu_407_p2;

assign zext_ln29_fu_346_p1 = or_ln29_fu_340_p2;

assign zext_ln33_1_fu_446_p1 = or_ln33_fu_440_p2;

assign zext_ln33_fu_425_p1 = q_reg_278;

endmodule //td_fused_top_tdf9_accum_1
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf9_accum_2 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        accum_in_2,
        accum_in_2_ap_vld,
        accum_in_address0,
        accum_in_ce0,
        accum_in_q0
);

parameter    ap_ST_fsm_state1 = 7'd1;
parameter    ap_ST_fsm_state2 = 7'd2;
parameter    ap_ST_fsm_state3 = 7'd4;
parameter    ap_ST_fsm_state4 = 7'd8;
parameter    ap_ST_fsm_state5 = 7'd16;
parameter    ap_ST_fsm_state6 = 7'd32;
parameter    ap_ST_fsm_state7 = 7'd64;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [15:0] accum_in_2;
output   accum_in_2_ap_vld;
output  [2:0] accum_in_address0;
output   accum_in_ce0;
input  [15:0] accum_in_q0;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg[15:0] accum_in_2;
reg accum_in_2_ap_vld;
reg accum_in_ce0;

reg    ap_done_reg;
  reg   [6:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
wire   [3:0] add_ln57_fu_74_p2;
reg   [3:0] add_ln57_reg_91;
wire    ap_CS_fsm_state2;
wire   [0:0] icmp_ln57_fu_85_p2;
wire    ap_CS_fsm_state3;
wire   [15:0] grp_fu_68_p2;
wire    ap_CS_fsm_state7;
reg   [3:0] i_1_1_reg_44;
reg    ap_block_state1;
reg   [15:0] sum_reg_55;
wire   [63:0] zext_ln57_fu_80_p1;
reg   [15:0] accum_in_2_preg;
reg   [6:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 7'd1;
#0 accum_in_2_preg = 16'd0;
end

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U568(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(sum_reg_55),
    .din1(accum_in_q0),
    .dout(grp_fu_68_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        accum_in_2_preg <= 16'd0;
    end else begin
        if (((icmp_ln57_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
            accum_in_2_preg <= sum_reg_55;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if (((icmp_ln57_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        i_1_1_reg_44 <= 4'd0;
    end else if ((1'b1 == ap_CS_fsm_state7)) begin
        i_1_1_reg_44 <= add_ln57_reg_91;
    end
end

always @ (posedge ap_clk) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        sum_reg_55 <= 16'd0;
    end else if ((1'b1 == ap_CS_fsm_state7)) begin
        sum_reg_55 <= grp_fu_68_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        add_ln57_reg_91 <= add_ln57_fu_74_p2;
    end
end

always @ (*) begin
    if (((icmp_ln57_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        accum_in_2 = sum_reg_55;
    end else begin
        accum_in_2 = accum_in_2_preg;
    end
end

always @ (*) begin
    if (((icmp_ln57_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        accum_in_2_ap_vld = 1'b1;
    end else begin
        accum_in_2_ap_vld = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        accum_in_ce0 = 1'b1;
    end else begin
        accum_in_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln57_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln57_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_state2 : begin
            if (((icmp_ln57_fu_85_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end
        end
        ap_ST_fsm_state3 : begin
            ap_NS_fsm = ap_ST_fsm_state4;
        end
        ap_ST_fsm_state4 : begin
            ap_NS_fsm = ap_ST_fsm_state5;
        end
        ap_ST_fsm_state5 : begin
            ap_NS_fsm = ap_ST_fsm_state6;
        end
        ap_ST_fsm_state6 : begin
            ap_NS_fsm = ap_ST_fsm_state7;
        end
        ap_ST_fsm_state7 : begin
            ap_NS_fsm = ap_ST_fsm_state2;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign accum_in_address0 = zext_ln57_fu_80_p1;

assign add_ln57_fu_74_p2 = (i_1_1_reg_44 + 4'd1);

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state7 = ap_CS_fsm[32'd6];

always @ (*) begin
    ap_block_state1 = ((ap_done_reg == 1'b1) | (ap_start == 1'b0));
end

assign icmp_ln57_fu_85_p2 = ((i_1_1_reg_44 == 4'd8) ? 1'b1 : 1'b0);

assign zext_ln57_fu_80_p1 = i_1_1_reg_44;

endmodule //td_fused_top_tdf9_accum_2
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_tdf9_adjustments_ram (addr0, ce0, q0, addr1, ce1, d1, we1,  clk);

parameter DWIDTH = 48;
parameter AWIDTH = 6;
parameter MEM_SIZE = 64;

input[AWIDTH-1:0] addr0;
input ce0;
output wire[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
input clk;

 reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];
wire [AWIDTH-1:0] addr0_t0; 
reg [AWIDTH-1:0] addr0_t1; 
reg [DWIDTH-1:0] q0_t0;
reg [DWIDTH-1:0] q0_t1;
wire [AWIDTH-1:0] addr1_t0; 
reg [AWIDTH-1:0] addr1_t1; 
wire [DWIDTH-1:0] d1_t0; 
wire we1_t0; 
reg [DWIDTH-1:0] d1_t1; 
reg we1_t1; 


assign addr0_t0 = addr0;
assign q0 = q0_t1;
assign addr1_t0 = addr1;
assign d1_t0 = d1;
assign we1_t0 = we1;

always @(posedge clk)  
begin
    if (ce0) 
    begin
        addr0_t1 <= addr0_t0; 
        q0_t1 <= q0_t0;
    end
    if (ce1) 
    begin
        addr1_t1 <= addr1_t0; 
        d1_t1 <= d1_t0;
        we1_t1 <= we1_t0;
    end
end


always @(posedge clk)  
begin 
    if (ce0) begin
        q0_t0 <= ram[addr0_t1];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1_t1) 
            ram[addr1_t1] <= d1_t1; 
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_tdf9_adjustments(
    reset,
    clk,
    address0,
    ce0,
    q0,
    address1,
    ce1,
    we1,
    d1);

parameter DataWidth = 32'd48;
parameter AddressRange = 32'd64;
parameter AddressWidth = 32'd6;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;



td_fused_top_tdf9_adjustments_ram td_fused_top_tdf9_adjustments_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 )
);

endmodule

// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf9_adjust (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        sums_read,
        adjustments_address0,
        adjustments_ce0,
        adjustments_q0,
        indices_23_dout,
        indices_23_empty_n,
        indices_23_read,
        ap_return
);

parameter    ap_ST_fsm_state1 = 17'd1;
parameter    ap_ST_fsm_state2 = 17'd2;
parameter    ap_ST_fsm_state3 = 17'd4;
parameter    ap_ST_fsm_state4 = 17'd8;
parameter    ap_ST_fsm_state5 = 17'd16;
parameter    ap_ST_fsm_state6 = 17'd32;
parameter    ap_ST_fsm_state7 = 17'd64;
parameter    ap_ST_fsm_state8 = 17'd128;
parameter    ap_ST_fsm_state9 = 17'd256;
parameter    ap_ST_fsm_state10 = 17'd512;
parameter    ap_ST_fsm_state11 = 17'd1024;
parameter    ap_ST_fsm_state12 = 17'd2048;
parameter    ap_ST_fsm_state13 = 17'd4096;
parameter    ap_ST_fsm_state14 = 17'd8192;
parameter    ap_ST_fsm_state15 = 17'd16384;
parameter    ap_ST_fsm_state16 = 17'd32768;
parameter    ap_ST_fsm_state17 = 17'd65536;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
input  [15:0] sums_read;
output  [5:0] adjustments_address0;
output   adjustments_ce0;
input  [47:0] adjustments_q0;
input  [5:0] indices_23_dout;
input   indices_23_empty_n;
output   indices_23_read;
output  [15:0] ap_return;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg adjustments_ce0;
reg indices_23_read;

reg    ap_done_reg;
  reg   [16:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    indices_23_blk_n;
wire    ap_CS_fsm_state4;
reg   [15:0] tmp_7_i_i_reg_167;
reg   [15:0] tmp_8_i_i_reg_172;
wire   [15:0] grp_fu_81_p2;
reg   [15:0] sub_i_i_i_reg_177;
wire    ap_CS_fsm_state8;
wire    ap_CS_fsm_state9;
wire   [15:0] grp_fu_86_p2;
reg   [15:0] mul_i_i_i_reg_187;
wire    ap_CS_fsm_state12;
wire    ap_CS_fsm_state13;
wire   [63:0] zext_ln220_fu_90_p1;
reg    ap_block_state1;
wire    ap_CS_fsm_state2;
wire    ap_CS_fsm_state3;
wire   [15:0] grp_fu_77_p1;
wire   [15:0] grp_fu_81_p1;
wire   [15:0] grp_fu_86_p1;
wire   [15:0] trunc_ln220_fu_95_p1;
wire   [15:0] grp_fu_77_p2;
wire    ap_CS_fsm_state17;
wire   [15:0] bitcast_ln648_fu_132_p1;
wire   [0:0] tmp_fu_136_p3;
reg   [16:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 17'd1;
end

td_fused_top_hadd_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hadd_16ns_16ns_16_5_full_dsp_1_U572(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(mul_i_i_i_reg_187),
    .din1(grp_fu_77_p1),
    .dout(grp_fu_77_p2)
);

td_fused_top_hsub_16ns_16ns_16_5_full_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 5 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hsub_16ns_16ns_16_5_full_dsp_1_U573(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(sums_read),
    .din1(grp_fu_81_p1),
    .dout(grp_fu_81_p2)
);

td_fused_top_hmul_16ns_16ns_16_4_max_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hmul_16ns_16ns_16_4_max_dsp_1_U574(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(sub_i_i_i_reg_177),
    .din1(grp_fu_86_p1),
    .dout(grp_fu_86_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state17)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state12)) begin
        mul_i_i_i_reg_187 <= grp_fu_86_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state8)) begin
        sub_i_i_i_reg_177 <= grp_fu_81_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        tmp_7_i_i_reg_167 <= {{adjustments_q0[31:16]}};
        tmp_8_i_i_reg_172 <= {{adjustments_q0[47:32]}};
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state2) | (~((indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1)))) begin
        adjustments_ce0 = 1'b1;
    end else begin
        adjustments_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state17)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state17)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_23_blk_n = indices_23_empty_n;
    end else begin
        indices_23_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_23_read = 1'b1;
    end else begin
        indices_23_read = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_state2 : begin
            ap_NS_fsm = ap_ST_fsm_state3;
        end
        ap_ST_fsm_state3 : begin
            ap_NS_fsm = ap_ST_fsm_state4;
        end
        ap_ST_fsm_state4 : begin
            ap_NS_fsm = ap_ST_fsm_state5;
        end
        ap_ST_fsm_state5 : begin
            ap_NS_fsm = ap_ST_fsm_state6;
        end
        ap_ST_fsm_state6 : begin
            ap_NS_fsm = ap_ST_fsm_state7;
        end
        ap_ST_fsm_state7 : begin
            ap_NS_fsm = ap_ST_fsm_state8;
        end
        ap_ST_fsm_state8 : begin
            ap_NS_fsm = ap_ST_fsm_state9;
        end
        ap_ST_fsm_state9 : begin
            ap_NS_fsm = ap_ST_fsm_state10;
        end
        ap_ST_fsm_state10 : begin
            ap_NS_fsm = ap_ST_fsm_state11;
        end
        ap_ST_fsm_state11 : begin
            ap_NS_fsm = ap_ST_fsm_state12;
        end
        ap_ST_fsm_state12 : begin
            ap_NS_fsm = ap_ST_fsm_state13;
        end
        ap_ST_fsm_state13 : begin
            ap_NS_fsm = ap_ST_fsm_state14;
        end
        ap_ST_fsm_state14 : begin
            ap_NS_fsm = ap_ST_fsm_state15;
        end
        ap_ST_fsm_state15 : begin
            ap_NS_fsm = ap_ST_fsm_state16;
        end
        ap_ST_fsm_state16 : begin
            ap_NS_fsm = ap_ST_fsm_state17;
        end
        ap_ST_fsm_state17 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign adjustments_address0 = zext_ln220_fu_90_p1;

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state12 = ap_CS_fsm[32'd11];

assign ap_CS_fsm_state13 = ap_CS_fsm[32'd12];

assign ap_CS_fsm_state17 = ap_CS_fsm[32'd16];

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

assign ap_CS_fsm_state8 = ap_CS_fsm[32'd7];

assign ap_CS_fsm_state9 = ap_CS_fsm[32'd8];

always @ (*) begin
    ap_block_state1 = ((indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0));
end

assign ap_return = ((tmp_fu_136_p3[0:0] == 1'b1) ? 16'd0 : grp_fu_77_p2);

assign bitcast_ln648_fu_132_p1 = grp_fu_77_p2;

assign grp_fu_77_p1 = tmp_8_i_i_reg_172;

assign grp_fu_81_p1 = trunc_ln220_fu_95_p1;

assign grp_fu_86_p1 = tmp_7_i_i_reg_167;

assign tmp_fu_136_p3 = bitcast_ln648_fu_132_p1[32'd15];

assign trunc_ln220_fu_95_p1 = adjustments_q0[15:0];

assign zext_ln220_fu_90_p1 = indices_23_dout;

endmodule //td_fused_top_tdf9_adjust
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf9_dot_product (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        ifmap_vec_0_0_address0,
        ifmap_vec_0_0_ce0,
        ifmap_vec_0_0_q0,
        weight_vecs_0_0_0_address0,
        weight_vecs_0_0_0_ce0,
        weight_vecs_0_0_0_q0,
        products_0_address0,
        products_0_ce0,
        products_0_we0,
        products_0_d0
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state9 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [7:0] ifmap_vec_0_0_address0;
output   ifmap_vec_0_0_ce0;
input  [15:0] ifmap_vec_0_0_q0;
output  [7:0] weight_vecs_0_0_0_address0;
output   weight_vecs_0_0_0_ce0;
input  [15:0] weight_vecs_0_0_0_q0;
output  [7:0] products_0_address0;
output   products_0_ce0;
output   products_0_we0;
output  [15:0] products_0_d0;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg ifmap_vec_0_0_ce0;
reg weight_vecs_0_0_0_ce0;
reg products_0_ce0;
reg products_0_we0;

reg    ap_done_reg;
  reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg   [8:0] ic_0_0_reg_69;
wire   [8:0] add_ln149_fu_84_p2;
wire    ap_CS_fsm_pp0_stage0;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
wire    ap_block_state4_pp0_stage0_iter2;
wire    ap_block_state5_pp0_stage0_iter3;
wire    ap_block_state6_pp0_stage0_iter4;
wire    ap_block_state7_pp0_stage0_iter5;
wire    ap_block_state8_pp0_stage0_iter6;
wire    ap_block_pp0_stage0_11001;
wire   [0:0] icmp_ln149_fu_90_p2;
reg   [0:0] icmp_ln149_reg_107;
reg   [0:0] icmp_ln149_reg_107_pp0_iter1_reg;
reg   [0:0] icmp_ln149_reg_107_pp0_iter2_reg;
reg   [0:0] icmp_ln149_reg_107_pp0_iter3_reg;
reg   [0:0] icmp_ln149_reg_107_pp0_iter4_reg;
reg   [0:0] icmp_ln149_reg_107_pp0_iter5_reg;
wire   [63:0] idxprom17_0_0_fu_96_p1;
reg   [63:0] idxprom17_0_0_reg_111;
reg   [63:0] idxprom17_0_0_reg_111_pp0_iter1_reg;
reg   [63:0] idxprom17_0_0_reg_111_pp0_iter2_reg;
reg   [63:0] idxprom17_0_0_reg_111_pp0_iter3_reg;
reg   [63:0] idxprom17_0_0_reg_111_pp0_iter4_reg;
reg   [63:0] idxprom17_0_0_reg_111_pp0_iter5_reg;
reg   [15:0] ifmap_vec_0_0_load_reg_126;
reg   [15:0] weight_vecs_0_0_0_load_reg_131;
wire   [15:0] grp_fu_80_p2;
reg   [15:0] mul_reg_136;
reg    ap_block_state1;
wire    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_exit_iter0_state2;
reg    ap_enable_reg_pp0_iter1;
reg    ap_enable_reg_pp0_iter2;
reg    ap_enable_reg_pp0_iter3;
reg    ap_enable_reg_pp0_iter4;
reg    ap_enable_reg_pp0_iter5;
reg    ap_enable_reg_pp0_iter6;
wire    ap_block_pp0_stage0;
wire    ap_CS_fsm_state9;
reg   [2:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
#0 ap_enable_reg_pp0_iter4 = 1'b0;
#0 ap_enable_reg_pp0_iter5 = 1'b0;
#0 ap_enable_reg_pp0_iter6 = 1'b0;
end

td_fused_top_hmul_16ns_16ns_16_4_max_dsp_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 16 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 16 ))
hmul_16ns_16ns_16_4_max_dsp_1_U560(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(1'b1),
    .din0(ifmap_vec_0_0_load_reg_126),
    .din1(weight_vecs_0_0_0_load_reg_131),
    .dout(grp_fu_80_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state9)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b1 == ap_condition_pp0_exit_iter0_state2))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            if ((1'b1 == ap_condition_pp0_exit_iter0_state2)) begin
                ap_enable_reg_pp0_iter1 <= (1'b1 ^ ap_condition_pp0_exit_iter0_state2);
            end else if ((1'b1 == 1'b1)) begin
                ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
            end
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter4 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter5 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter5 <= ap_enable_reg_pp0_iter4;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter6 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter6 <= ap_enable_reg_pp0_iter5;
        end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter6 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln149_fu_90_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ic_0_0_reg_69 <= add_ln149_fu_84_p2;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ic_0_0_reg_69 <= 9'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln149_reg_107 <= icmp_ln149_fu_90_p2;
        icmp_ln149_reg_107_pp0_iter1_reg <= icmp_ln149_reg_107;
        idxprom17_0_0_reg_111_pp0_iter1_reg[8 : 0] <= idxprom17_0_0_reg_111[8 : 0];
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        icmp_ln149_reg_107_pp0_iter2_reg <= icmp_ln149_reg_107_pp0_iter1_reg;
        icmp_ln149_reg_107_pp0_iter3_reg <= icmp_ln149_reg_107_pp0_iter2_reg;
        icmp_ln149_reg_107_pp0_iter4_reg <= icmp_ln149_reg_107_pp0_iter3_reg;
        icmp_ln149_reg_107_pp0_iter5_reg <= icmp_ln149_reg_107_pp0_iter4_reg;
        idxprom17_0_0_reg_111_pp0_iter2_reg[8 : 0] <= idxprom17_0_0_reg_111_pp0_iter1_reg[8 : 0];
        idxprom17_0_0_reg_111_pp0_iter3_reg[8 : 0] <= idxprom17_0_0_reg_111_pp0_iter2_reg[8 : 0];
        idxprom17_0_0_reg_111_pp0_iter4_reg[8 : 0] <= idxprom17_0_0_reg_111_pp0_iter3_reg[8 : 0];
        idxprom17_0_0_reg_111_pp0_iter5_reg[8 : 0] <= idxprom17_0_0_reg_111_pp0_iter4_reg[8 : 0];
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln149_fu_90_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        idxprom17_0_0_reg_111[8 : 0] <= idxprom17_0_0_fu_96_p1[8 : 0];
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln149_reg_107 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ifmap_vec_0_0_load_reg_126 <= ifmap_vec_0_0_q0;
        weight_vecs_0_0_0_load_reg_131 <= weight_vecs_0_0_0_q0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln149_reg_107_pp0_iter4_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        mul_reg_136 <= grp_fu_80_p2;
    end
end

always @ (*) begin
    if ((icmp_ln149_fu_90_p2 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state2 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state2 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state9)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state9)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ifmap_vec_0_0_ce0 = 1'b1;
    end else begin
        ifmap_vec_0_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter6 == 1'b1))) begin
        products_0_ce0 = 1'b1;
    end else begin
        products_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln149_reg_107_pp0_iter5_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter6 == 1'b1))) begin
        products_0_we0 = 1'b1;
    end else begin
        products_0_we0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        weight_vecs_0_0_0_ce0 = 1'b1;
    end else begin
        weight_vecs_0_0_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((~((icmp_ln149_fu_90_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0)) & ~((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter6 == 1'b1) & (ap_enable_reg_pp0_iter5 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if ((((icmp_ln149_fu_90_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0)) | ((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter6 == 1'b1) & (ap_enable_reg_pp0_iter5 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_state9;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state9 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln149_fu_84_p2 = (ic_0_0_reg_69 + 9'd1);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state9 = ap_CS_fsm[32'd2];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (ap_done_reg == 1'b1));
end

assign ap_block_state2_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter4 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage0_iter5 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage0_iter6 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign icmp_ln149_fu_90_p2 = ((ic_0_0_reg_69 == 9'd256) ? 1'b1 : 1'b0);

assign idxprom17_0_0_fu_96_p1 = ic_0_0_reg_69;

assign ifmap_vec_0_0_address0 = idxprom17_0_0_fu_96_p1;

assign products_0_address0 = idxprom17_0_0_reg_111_pp0_iter5_reg;

assign products_0_d0 = mul_reg_136;

assign weight_vecs_0_0_0_address0 = idxprom17_0_0_fu_96_p1;

always @ (posedge ap_clk) begin
    idxprom17_0_0_reg_111[63:9] <= 55'b0000000000000000000000000000000000000000000000000000000;
    idxprom17_0_0_reg_111_pp0_iter1_reg[63:9] <= 55'b0000000000000000000000000000000000000000000000000000000;
    idxprom17_0_0_reg_111_pp0_iter2_reg[63:9] <= 55'b0000000000000000000000000000000000000000000000000000000;
    idxprom17_0_0_reg_111_pp0_iter3_reg[63:9] <= 55'b0000000000000000000000000000000000000000000000000000000;
    idxprom17_0_0_reg_111_pp0_iter4_reg[63:9] <= 55'b0000000000000000000000000000000000000000000000000000000;
    idxprom17_0_0_reg_111_pp0_iter5_reg[63:9] <= 55'b0000000000000000000000000000000000000000000000000000000;
end

endmodule //td_fused_top_tdf9_dot_product
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_tdf9_filters_ram (addr0, ce0, q0, addr1, ce1, d1, we1,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 14;
parameter MEM_SIZE = 16384;

input[AWIDTH-1:0] addr0;
input ce0;
output wire[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
input clk;

 reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];
wire [AWIDTH-1:0] addr0_t0; 
reg [AWIDTH-1:0] addr0_t1; 
reg [DWIDTH-1:0] q0_t0;
reg [DWIDTH-1:0] q0_t1;
wire [AWIDTH-1:0] addr1_t0; 
reg [AWIDTH-1:0] addr1_t1; 
wire [DWIDTH-1:0] d1_t0; 
wire we1_t0; 
reg [DWIDTH-1:0] d1_t1; 
reg we1_t1; 


assign addr0_t0 = addr0;
assign q0 = q0_t1;
assign addr1_t0 = addr1;
assign d1_t0 = d1;
assign we1_t0 = we1;

always @(posedge clk)  
begin
    if (ce0) 
    begin
        addr0_t1 <= addr0_t0; 
        q0_t1 <= q0_t0;
    end
    if (ce1) 
    begin
        addr1_t1 <= addr1_t0; 
        d1_t1 <= d1_t0;
        we1_t1 <= we1_t0;
    end
end


always @(posedge clk)  
begin 
    if (ce0) begin
        q0_t0 <= ram[addr0_t1];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1_t1) 
            ram[addr1_t1] <= d1_t1; 
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_tdf9_filters(
    reset,
    clk,
    address0,
    ce0,
    q0,
    address1,
    ce1,
    we1,
    d1);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd16384;
parameter AddressWidth = 32'd14;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;



td_fused_top_tdf9_filters_ram td_fused_top_tdf9_filters_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 )
);

endmodule

// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf9_get_next_ijk (
        ap_clk,
        ap_rst,
        ap_start,
        start_full_n,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        start_out,
        start_write,
        indices_0_din,
        indices_0_full_n,
        indices_0_write,
        indices_1_din,
        indices_1_full_n,
        indices_1_write,
        indices_2_out_din,
        indices_2_out_full_n,
        indices_2_out_write,
        indices_2_out1_din,
        indices_2_out1_full_n,
        indices_2_out1_write
);

parameter    ap_ST_fsm_state1 = 1'd1;

input   ap_clk;
input   ap_rst;
input   ap_start;
input   start_full_n;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output   start_out;
output   start_write;
output  [15:0] indices_0_din;
input   indices_0_full_n;
output   indices_0_write;
output  [15:0] indices_1_din;
input   indices_1_full_n;
output   indices_1_write;
output  [5:0] indices_2_out_din;
input   indices_2_out_full_n;
output   indices_2_out_write;
output  [5:0] indices_2_out1_din;
input   indices_2_out1_full_n;
output   indices_2_out1_write;

reg ap_done;
reg ap_idle;
reg start_write;
reg indices_0_write;
reg indices_1_write;
reg indices_2_out_write;
reg indices_2_out1_write;

reg    real_start;
reg    start_once_reg;
reg    ap_done_reg;
  reg   [0:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    internal_ap_ready;
reg   [15:0] i;
reg   [15:0] j;
reg   [15:0] k;
reg    indices_0_blk_n;
reg    indices_1_blk_n;
reg    indices_2_out_blk_n;
reg    indices_2_out1_blk_n;
reg   [0:0] ap_phi_mux_j_flag_0_i_phi_fu_77_p6;
reg    ap_block_state1;
wire   [0:0] icmp_ln78_fu_141_p2;
wire   [0:0] icmp_ln81_fu_154_p2;
reg   [15:0] ap_phi_mux_j_new_0_i_phi_fu_91_p6;
wire   [15:0] add_ln80_fu_147_p2;
reg   [15:0] ap_phi_mux_k_new_0_i_phi_fu_104_p6;
wire   [15:0] add_ln77_fu_134_p2;
wire   [15:0] select_ln84_fu_172_p3;
wire   [5:0] trunc_ln76_fu_128_p1;
wire   [15:0] add_ln83_fu_160_p2;
wire   [0:0] icmp_ln84_fu_166_p2;
reg   [0:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 start_once_reg = 1'b0;
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 1'd1;
#0 i = 16'd0;
#0 j = 16'd0;
#0 k = 16'd0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((~((real_start == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        start_once_reg <= 1'b0;
    end else begin
        if (((real_start == 1'b1) & (internal_ap_ready == 1'b0))) begin
            start_once_reg <= 1'b1;
        end else if ((internal_ap_ready == 1'b1)) begin
            start_once_reg <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((~((real_start == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (icmp_ln81_fu_154_p2 == 1'd1) & (icmp_ln78_fu_141_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1))) begin
        i <= select_ln84_fu_172_p3;
    end
end

always @ (posedge ap_clk) begin
    if ((~((real_start == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (ap_phi_mux_j_flag_0_i_phi_fu_77_p6 == 1'd1) & (1'b1 == ap_CS_fsm_state1))) begin
        j <= ap_phi_mux_j_new_0_i_phi_fu_91_p6;
    end
end

always @ (posedge ap_clk) begin
    if ((~((real_start == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        k <= ap_phi_mux_k_new_0_i_phi_fu_104_p6;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((real_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln78_fu_141_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_phi_mux_j_flag_0_i_phi_fu_77_p6 = 1'd0;
    end else if ((((icmp_ln81_fu_154_p2 == 1'd0) & (icmp_ln78_fu_141_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1)) | ((icmp_ln81_fu_154_p2 == 1'd1) & (icmp_ln78_fu_141_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1)))) begin
        ap_phi_mux_j_flag_0_i_phi_fu_77_p6 = 1'd1;
    end else begin
        ap_phi_mux_j_flag_0_i_phi_fu_77_p6 = 'bx;
    end
end

always @ (*) begin
    if (((icmp_ln78_fu_141_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1))) begin
        if ((icmp_ln81_fu_154_p2 == 1'd0)) begin
            ap_phi_mux_j_new_0_i_phi_fu_91_p6 = add_ln80_fu_147_p2;
        end else if ((icmp_ln81_fu_154_p2 == 1'd1)) begin
            ap_phi_mux_j_new_0_i_phi_fu_91_p6 = 16'd0;
        end else begin
            ap_phi_mux_j_new_0_i_phi_fu_91_p6 = 'bx;
        end
    end else begin
        ap_phi_mux_j_new_0_i_phi_fu_91_p6 = 'bx;
    end
end

always @ (*) begin
    if (((icmp_ln78_fu_141_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_phi_mux_k_new_0_i_phi_fu_104_p6 = add_ln77_fu_134_p2;
    end else if ((((icmp_ln81_fu_154_p2 == 1'd0) & (icmp_ln78_fu_141_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1)) | ((icmp_ln81_fu_154_p2 == 1'd1) & (icmp_ln78_fu_141_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1)))) begin
        ap_phi_mux_k_new_0_i_phi_fu_104_p6 = 16'd0;
    end else begin
        ap_phi_mux_k_new_0_i_phi_fu_104_p6 = 'bx;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_0_blk_n = indices_0_full_n;
    end else begin
        indices_0_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_0_write = 1'b1;
    end else begin
        indices_0_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_1_blk_n = indices_1_full_n;
    end else begin
        indices_1_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_1_write = 1'b1;
    end else begin
        indices_1_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_2_out1_blk_n = indices_2_out1_full_n;
    end else begin
        indices_2_out1_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_2_out1_write = 1'b1;
    end else begin
        indices_2_out1_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_2_out_blk_n = indices_2_out_full_n;
    end else begin
        indices_2_out_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_2_out_write = 1'b1;
    end else begin
        indices_2_out_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((real_start == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        internal_ap_ready = 1'b1;
    end else begin
        internal_ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((start_full_n == 1'b0) & (start_once_reg == 1'b0))) begin
        real_start = 1'b0;
    end else begin
        real_start = ap_start;
    end
end

always @ (*) begin
    if (((real_start == 1'b1) & (start_once_reg == 1'b0))) begin
        start_write = 1'b1;
    end else begin
        start_write = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln77_fu_134_p2 = (k + 16'd1);

assign add_ln80_fu_147_p2 = (j + 16'd1);

assign add_ln83_fu_160_p2 = (i + 16'd1);

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

always @ (*) begin
    ap_block_state1 = ((real_start == 1'b0) | (indices_2_out1_full_n == 1'b0) | (indices_2_out_full_n == 1'b0) | (indices_1_full_n == 1'b0) | (indices_0_full_n == 1'b0) | (ap_done_reg == 1'b1));
end

assign ap_ready = internal_ap_ready;

assign icmp_ln78_fu_141_p2 = ((add_ln77_fu_134_p2 == 16'd64) ? 1'b1 : 1'b0);

assign icmp_ln81_fu_154_p2 = ((add_ln80_fu_147_p2 == 16'd14) ? 1'b1 : 1'b0);

assign icmp_ln84_fu_166_p2 = ((add_ln83_fu_160_p2 == 16'd14) ? 1'b1 : 1'b0);

assign indices_0_din = i;

assign indices_1_din = j;

assign indices_2_out1_din = trunc_ln76_fu_128_p1;

assign indices_2_out_din = trunc_ln76_fu_128_p1;

assign select_ln84_fu_172_p3 = ((icmp_ln84_fu_166_p2[0:0] == 1'b1) ? 16'd0 : add_ln83_fu_160_p2);

assign start_out = real_start;

assign trunc_ln76_fu_128_p1 = k[5:0];

endmodule //td_fused_top_tdf9_get_next_ijk
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf9_readFilters62 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        filter_data_address0,
        filter_data_ce0,
        filter_data_q0,
        indices_23_dout,
        indices_23_empty_n,
        indices_23_read,
        weight_vecs_0_0_0_address0,
        weight_vecs_0_0_0_ce0,
        weight_vecs_0_0_0_we0,
        weight_vecs_0_0_0_d0
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state6 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [13:0] filter_data_address0;
output   filter_data_ce0;
input  [15:0] filter_data_q0;
input  [5:0] indices_23_dout;
input   indices_23_empty_n;
output   indices_23_read;
output  [7:0] weight_vecs_0_0_0_address0;
output   weight_vecs_0_0_0_ce0;
output   weight_vecs_0_0_0_we0;
output  [15:0] weight_vecs_0_0_0_d0;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg filter_data_ce0;
reg indices_23_read;
reg weight_vecs_0_0_0_ce0;
reg weight_vecs_0_0_0_we0;

reg    ap_done_reg;
  reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    indices_23_blk_n;
reg   [8:0] kk_0_0_i_i_reg_93;
reg   [8:0] kk_0_0_i_i_reg_93_pp0_iter1_reg;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
wire    ap_block_state4_pp0_stage0_iter2;
wire    ap_block_state5_pp0_stage0_iter3;
wire    ap_block_pp0_stage0_11001;
reg   [8:0] kk_0_0_i_i_reg_93_pp0_iter2_reg;
wire   [13:0] tmp_fu_105_p3;
reg   [13:0] tmp_reg_144;
wire   [8:0] add_ln49_fu_113_p2;
reg   [8:0] add_ln49_reg_149;
reg    ap_enable_reg_pp0_iter0;
wire   [0:0] icmp_ln49_fu_119_p2;
reg   [0:0] icmp_ln49_reg_154;
reg   [0:0] icmp_ln49_reg_154_pp0_iter1_reg;
reg   [0:0] icmp_ln49_reg_154_pp0_iter2_reg;
reg    ap_block_state1;
wire    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_exit_iter0_state2;
reg    ap_enable_reg_pp0_iter1;
reg    ap_enable_reg_pp0_iter2;
reg    ap_enable_reg_pp0_iter3;
reg   [8:0] ap_phi_mux_kk_0_0_i_i_phi_fu_97_p4;
wire    ap_block_pp0_stage0;
wire   [63:0] zext_ln55_1_fu_134_p1;
wire   [63:0] idxprom16_0_0_i_i_fu_139_p1;
wire   [13:0] zext_ln55_fu_125_p1;
wire   [13:0] add_ln55_fu_129_p2;
wire    ap_CS_fsm_state6;
reg   [2:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state6)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_condition_pp0_exit_iter0_state2) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            if ((1'b1 == ap_condition_pp0_exit_iter0_state2)) begin
                ap_enable_reg_pp0_iter1 <= (1'b1 ^ ap_condition_pp0_exit_iter0_state2);
            end else if ((1'b1 == 1'b1)) begin
                ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
            end
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end else if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter3 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln49_reg_154 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        kk_0_0_i_i_reg_93 <= add_ln49_reg_149;
    end else if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        kk_0_0_i_i_reg_93 <= 9'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        add_ln49_reg_149 <= add_ln49_fu_113_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln49_reg_154 <= icmp_ln49_fu_119_p2;
        icmp_ln49_reg_154_pp0_iter1_reg <= icmp_ln49_reg_154;
        kk_0_0_i_i_reg_93_pp0_iter1_reg <= kk_0_0_i_i_reg_93;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        icmp_ln49_reg_154_pp0_iter2_reg <= icmp_ln49_reg_154_pp0_iter1_reg;
        kk_0_0_i_i_reg_93_pp0_iter2_reg <= kk_0_0_i_i_reg_93_pp0_iter1_reg;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state1)) begin
        tmp_reg_144[13 : 8] <= tmp_fu_105_p3[13 : 8];
    end
end

always @ (*) begin
    if ((icmp_ln49_fu_119_p2 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state2 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state2 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state6)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln49_reg_154 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_kk_0_0_i_i_phi_fu_97_p4 = add_ln49_reg_149;
    end else begin
        ap_phi_mux_kk_0_0_i_i_phi_fu_97_p4 = kk_0_0_i_i_reg_93;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state6)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter3 == 1'b1)))) begin
        filter_data_ce0 = 1'b1;
    end else begin
        filter_data_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_23_blk_n = indices_23_empty_n;
    end else begin
        indices_23_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_23_read = 1'b1;
    end else begin
        indices_23_read = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter3 == 1'b1))) begin
        weight_vecs_0_0_0_ce0 = 1'b1;
    end else begin
        weight_vecs_0_0_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln49_reg_154_pp0_iter2_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter3 == 1'b1))) begin
        weight_vecs_0_0_0_we0 = 1'b1;
    end else begin
        weight_vecs_0_0_0_we0 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((~((icmp_ln49_fu_119_p2 == 1'd1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter1 == 1'b0)) & ~((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter3 == 1'b1) & (ap_enable_reg_pp0_iter2 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if ((((icmp_ln49_fu_119_p2 == 1'd1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter1 == 1'b0)) | ((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter3 == 1'b1) & (ap_enable_reg_pp0_iter2 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_state6;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state6 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln49_fu_113_p2 = (ap_phi_mux_kk_0_0_i_i_phi_fu_97_p4 + 9'd1);

assign add_ln55_fu_129_p2 = (tmp_reg_144 + zext_ln55_fu_125_p1);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state6 = ap_CS_fsm[32'd2];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (indices_23_empty_n == 1'b0) | (ap_done_reg == 1'b1));
end

assign ap_block_state2_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign filter_data_address0 = zext_ln55_1_fu_134_p1;

assign icmp_ln49_fu_119_p2 = ((ap_phi_mux_kk_0_0_i_i_phi_fu_97_p4 == 9'd256) ? 1'b1 : 1'b0);

assign idxprom16_0_0_i_i_fu_139_p1 = kk_0_0_i_i_reg_93_pp0_iter2_reg;

assign tmp_fu_105_p3 = {{indices_23_dout}, {8'd0}};

assign weight_vecs_0_0_0_address0 = idxprom16_0_0_i_i_fu_139_p1;

assign weight_vecs_0_0_0_d0 = filter_data_q0;

assign zext_ln55_1_fu_134_p1 = add_ln55_fu_129_p2;

assign zext_ln55_fu_125_p1 = ap_phi_mux_kk_0_0_i_i_phi_fu_97_p4;

always @ (posedge ap_clk) begin
    tmp_reg_144[7:0] <= 8'b00000000;
end

endmodule //td_fused_top_tdf9_readFilters62
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf9_readInputs (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        in_data_address0,
        in_data_ce0,
        in_data_q0,
        indices_01_dout,
        indices_01_empty_n,
        indices_01_read,
        indices_12_dout,
        indices_12_empty_n,
        indices_12_read,
        ifmap_vec_0_0_address0,
        ifmap_vec_0_0_ce0,
        ifmap_vec_0_0_we0,
        ifmap_vec_0_0_d0,
        ifmap_vec_0_0_address1,
        ifmap_vec_0_0_ce1,
        ifmap_vec_0_0_we1,
        ifmap_vec_0_0_d1,
        indices_01_out_din,
        indices_01_out_full_n,
        indices_01_out_write,
        indices_12_out_din,
        indices_12_out_full_n,
        indices_12_out_write
);

parameter    ap_ST_fsm_state1 = 5'd1;
parameter    ap_ST_fsm_state2 = 5'd2;
parameter    ap_ST_fsm_pp0_stage0 = 5'd4;
parameter    ap_ST_fsm_pp0_stage1 = 5'd8;
parameter    ap_ST_fsm_state8 = 5'd16;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [13:0] in_data_address0;
output   in_data_ce0;
input  [63:0] in_data_q0;
input  [15:0] indices_01_dout;
input   indices_01_empty_n;
output   indices_01_read;
input  [15:0] indices_12_dout;
input   indices_12_empty_n;
output   indices_12_read;
output  [7:0] ifmap_vec_0_0_address0;
output   ifmap_vec_0_0_ce0;
output   ifmap_vec_0_0_we0;
output  [15:0] ifmap_vec_0_0_d0;
output  [7:0] ifmap_vec_0_0_address1;
output   ifmap_vec_0_0_ce1;
output   ifmap_vec_0_0_we1;
output  [15:0] ifmap_vec_0_0_d1;
output  [3:0] indices_01_out_din;
input   indices_01_out_full_n;
output   indices_01_out_write;
output  [7:0] indices_12_out_din;
input   indices_12_out_full_n;
output   indices_12_out_write;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg in_data_ce0;
reg indices_01_read;
reg indices_12_read;
reg[7:0] ifmap_vec_0_0_address0;
reg ifmap_vec_0_0_ce0;
reg ifmap_vec_0_0_we0;
reg[15:0] ifmap_vec_0_0_d0;
reg[7:0] ifmap_vec_0_0_address1;
reg ifmap_vec_0_0_ce1;
reg ifmap_vec_0_0_we1;
reg[15:0] ifmap_vec_0_0_d1;
reg indices_01_out_write;
reg indices_12_out_write;

reg    ap_done_reg;
  reg   [4:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    indices_01_blk_n;
reg    indices_12_blk_n;
reg    indices_01_out_blk_n;
reg    indices_12_out_blk_n;
reg   [8:0] kk_0_i_i_reg_180;
reg   [8:0] kk_0_i_i_reg_180_pp0_iter1_reg;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_block_state3_pp0_stage0_iter0;
wire    ap_block_state5_pp0_stage0_iter1;
wire    ap_block_state7_pp0_stage0_iter2;
wire    ap_block_pp0_stage0_11001;
wire   [3:0] trunc_ln135_fu_192_p1;
reg   [3:0] trunc_ln135_reg_434;
reg   [15:0] col_coord_reg_439;
wire   [0:0] is_padding_fu_214_p2;
reg   [0:0] is_padding_reg_444;
wire   [9:0] add_ln32_fu_274_p2;
reg   [9:0] add_ln32_reg_454;
wire    ap_CS_fsm_state2;
wire   [0:0] icmp_ln25_fu_280_p2;
reg   [0:0] icmp_ln25_reg_459;
reg   [0:0] icmp_ln25_reg_459_pp0_iter1_reg;
wire   [8:0] add_ln25_fu_308_p2;
reg   [8:0] add_ln25_reg_468;
wire    ap_CS_fsm_pp0_stage1;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_state4_pp0_stage1_iter0;
wire    ap_block_state6_pp0_stage1_iter1;
wire    ap_block_pp0_stage1_11001;
wire   [7:0] empty_56_fu_314_p1;
reg   [7:0] empty_56_reg_473;
wire   [15:0] select_ln33_2_fu_386_p3;
reg   [15:0] select_ln33_2_reg_479;
wire   [15:0] select_ln33_3_fu_407_p3;
reg   [15:0] select_ln33_3_reg_484;
wire    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_exit_iter0_state3;
reg    ap_enable_reg_pp0_iter1;
wire    ap_block_pp0_stage1_subdone;
reg    ap_enable_reg_pp0_iter2;
reg   [8:0] ap_phi_mux_kk_0_i_i_phi_fu_184_p4;
wire    ap_block_pp0_stage0;
wire   [63:0] sext_ln32_fu_303_p1;
wire   [63:0] zext_ln32_fu_318_p1;
wire    ap_block_pp0_stage1;
wire   [63:0] zext_ln32_2_fu_345_p1;
wire   [63:0] zext_ln32_3_fu_419_p1;
wire   [63:0] zext_ln32_4_fu_429_p1;
reg    ap_block_state1;
wire   [15:0] select_ln33_fu_331_p3;
wire   [15:0] select_ln33_1_fu_364_p3;
wire   [0:0] cmp7_i_i_fu_202_p2;
wire   [0:0] icmp_ln24_fu_208_p2;
wire   [3:0] empty_54_fu_220_p1;
wire   [3:0] row_coord_int_fu_223_p3;
wire   [7:0] tmp_fu_236_p3;
wire   [4:0] tmp_4_fu_248_p3;
wire   [8:0] zext_ln32_1_fu_244_p1;
wire   [8:0] zext_ln32_5_fu_256_p1;
wire   [8:0] sub_ln32_fu_260_p2;
wire   [3:0] col_coord_int_fu_229_p3;
wire   [9:0] sub_ln32_cast_fu_266_p1;
wire   [9:0] zext_ln32_6_fu_270_p1;
wire   [5:0] lshr_ln_fu_286_p4;
wire   [15:0] tmp_1_fu_296_p3;
wire   [15:0] trunc_ln32_fu_323_p1;
wire   [15:0] bitcast_ln32_fu_327_p1;
wire   [7:0] or_ln25_fu_339_p2;
wire   [15:0] tmp_4_i_i_fu_350_p4;
wire   [15:0] bitcast_ln32_1_fu_360_p1;
wire   [15:0] tmp_5_i_i_fu_372_p4;
wire   [15:0] bitcast_ln32_2_fu_382_p1;
wire   [15:0] tmp_6_i_i_fu_393_p4;
wire   [15:0] bitcast_ln32_3_fu_403_p1;
wire   [7:0] or_ln25_1_fu_414_p2;
wire   [7:0] or_ln25_2_fu_424_p2;
wire    ap_CS_fsm_state8;
reg   [4:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 5'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state8)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b1 == ap_condition_pp0_exit_iter0_state3))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1)) | ((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b0)))) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end else if ((1'b1 == ap_CS_fsm_state2)) begin
            ap_enable_reg_pp0_iter2 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln25_reg_459 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        kk_0_i_i_reg_180 <= add_ln25_reg_468;
    end else if ((1'b1 == ap_CS_fsm_state2)) begin
        kk_0_i_i_reg_180 <= 9'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln25_reg_459 == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
        add_ln25_reg_468 <= add_ln25_fu_308_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        add_ln32_reg_454 <= add_ln32_fu_274_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state1)) begin
        col_coord_reg_439 <= indices_12_dout;
        is_padding_reg_444 <= is_padding_fu_214_p2;
        trunc_ln135_reg_434 <= trunc_ln135_fu_192_p1;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln25_reg_459_pp0_iter1_reg == 1'd0))) begin
        empty_56_reg_473 <= empty_56_fu_314_p1;
        select_ln33_2_reg_479 <= select_ln33_2_fu_386_p3;
        select_ln33_3_reg_484 <= select_ln33_3_fu_407_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln25_reg_459 <= icmp_ln25_fu_280_p2;
        icmp_ln25_reg_459_pp0_iter1_reg <= icmp_ln25_reg_459;
        kk_0_i_i_reg_180_pp0_iter1_reg <= kk_0_i_i_reg_180;
    end
end

always @ (*) begin
    if ((icmp_ln25_fu_280_p2 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state3 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state3 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state8)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln25_reg_459 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ap_phi_mux_kk_0_i_i_phi_fu_184_p4 = add_ln25_reg_468;
    end else begin
        ap_phi_mux_kk_0_i_i_phi_fu_184_p4 = kk_0_i_i_reg_180;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state8)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        ifmap_vec_0_0_address0 = zext_ln32_4_fu_429_p1;
    end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ifmap_vec_0_0_address0 = zext_ln32_2_fu_345_p1;
    end else begin
        ifmap_vec_0_0_address0 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        ifmap_vec_0_0_address1 = zext_ln32_3_fu_419_p1;
    end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ifmap_vec_0_0_address1 = zext_ln32_fu_318_p1;
    end else begin
        ifmap_vec_0_0_address1 = 'bx;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1)) | ((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1)))) begin
        ifmap_vec_0_0_ce0 = 1'b1;
    end else begin
        ifmap_vec_0_0_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1)) | ((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1)))) begin
        ifmap_vec_0_0_ce1 = 1'b1;
    end else begin
        ifmap_vec_0_0_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        ifmap_vec_0_0_d0 = select_ln33_3_reg_484;
    end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ifmap_vec_0_0_d0 = select_ln33_1_fu_364_p3;
    end else begin
        ifmap_vec_0_0_d0 = 'bx;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        ifmap_vec_0_0_d1 = select_ln33_2_reg_479;
    end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        ifmap_vec_0_0_d1 = select_ln33_fu_331_p3;
    end else begin
        ifmap_vec_0_0_d1 = 'bx;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1) & (icmp_ln25_reg_459_pp0_iter1_reg == 1'd0)) | ((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln25_reg_459_pp0_iter1_reg == 1'd0)))) begin
        ifmap_vec_0_0_we0 = 1'b1;
    end else begin
        ifmap_vec_0_0_we0 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1) & (icmp_ln25_reg_459_pp0_iter1_reg == 1'd0)) | ((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln25_reg_459_pp0_iter1_reg == 1'd0)))) begin
        ifmap_vec_0_0_we1 = 1'b1;
    end else begin
        ifmap_vec_0_0_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1)) | ((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1)) | ((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1)) | ((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1)))) begin
        in_data_ce0 = 1'b1;
    end else begin
        in_data_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_01_blk_n = indices_01_empty_n;
    end else begin
        indices_01_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_01_out_blk_n = indices_01_out_full_n;
    end else begin
        indices_01_out_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((indices_12_out_full_n == 1'b0) | (indices_01_out_full_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_01_out_write = 1'b1;
    end else begin
        indices_01_out_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((indices_12_out_full_n == 1'b0) | (indices_01_out_full_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_01_read = 1'b1;
    end else begin
        indices_01_read = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_12_blk_n = indices_12_empty_n;
    end else begin
        indices_12_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_12_out_blk_n = indices_12_out_full_n;
    end else begin
        indices_12_out_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((indices_12_out_full_n == 1'b0) | (indices_01_out_full_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_12_out_write = 1'b1;
    end else begin
        indices_12_out_write = 1'b0;
    end
end

always @ (*) begin
    if ((~((indices_12_out_full_n == 1'b0) | (indices_01_out_full_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_12_read = 1'b1;
    end else begin
        indices_12_read = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((indices_12_out_full_n == 1'b0) | (indices_01_out_full_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_state2 : begin
            ap_NS_fsm = ap_ST_fsm_pp0_stage0;
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((~((icmp_ln25_fu_280_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1)) & ~((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0)) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end else if ((((icmp_ln25_fu_280_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1)) | ((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter2 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0)))) begin
                ap_NS_fsm = ap_ST_fsm_state8;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_pp0_stage1 : begin
            if ((1'b0 == ap_block_pp0_stage1_subdone)) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end
        end
        ap_ST_fsm_state8 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln25_fu_308_p2 = (kk_0_i_i_reg_180 + 9'd4);

assign add_ln32_fu_274_p2 = ((sub_ln32_cast_fu_266_p1) + (zext_ln32_6_fu_270_p1));

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_pp0_stage1 = ap_CS_fsm[32'd3];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state8 = ap_CS_fsm[32'd4];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((indices_12_out_full_n == 1'b0) | (indices_01_out_full_n == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1) | (ap_start == 1'b0));
end

assign ap_block_state3_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage1_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage1_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign bitcast_ln32_1_fu_360_p1 = tmp_4_i_i_fu_350_p4;

assign bitcast_ln32_2_fu_382_p1 = tmp_5_i_i_fu_372_p4;

assign bitcast_ln32_3_fu_403_p1 = tmp_6_i_i_fu_393_p4;

assign bitcast_ln32_fu_327_p1 = trunc_ln32_fu_323_p1;

assign cmp7_i_i_fu_202_p2 = ((indices_01_dout > 16'd13) ? 1'b1 : 1'b0);

assign col_coord_int_fu_229_p3 = ((is_padding_reg_444[0:0] == 1'b1) ? 4'd0 : empty_54_fu_220_p1);

assign empty_54_fu_220_p1 = col_coord_reg_439[3:0];

assign empty_56_fu_314_p1 = kk_0_i_i_reg_180_pp0_iter1_reg[7:0];

assign icmp_ln24_fu_208_p2 = ((indices_12_dout > 16'd13) ? 1'b1 : 1'b0);

assign icmp_ln25_fu_280_p2 = ((ap_phi_mux_kk_0_i_i_phi_fu_184_p4 == 9'd256) ? 1'b1 : 1'b0);

assign in_data_address0 = sext_ln32_fu_303_p1;

assign indices_01_out_din = indices_01_dout[3:0];

assign indices_12_out_din = indices_12_dout[7:0];

assign is_padding_fu_214_p2 = (icmp_ln24_fu_208_p2 | cmp7_i_i_fu_202_p2);

assign lshr_ln_fu_286_p4 = {{ap_phi_mux_kk_0_i_i_phi_fu_184_p4[7:2]}};

assign or_ln25_1_fu_414_p2 = (empty_56_reg_473 | 8'd2);

assign or_ln25_2_fu_424_p2 = (empty_56_reg_473 | 8'd3);

assign or_ln25_fu_339_p2 = (empty_56_fu_314_p1 | 8'd1);

assign row_coord_int_fu_223_p3 = ((is_padding_reg_444[0:0] == 1'b1) ? 4'd0 : trunc_ln135_reg_434);

assign select_ln33_1_fu_364_p3 = ((is_padding_reg_444[0:0] == 1'b1) ? 16'd0 : bitcast_ln32_1_fu_360_p1);

assign select_ln33_2_fu_386_p3 = ((is_padding_reg_444[0:0] == 1'b1) ? 16'd0 : bitcast_ln32_2_fu_382_p1);

assign select_ln33_3_fu_407_p3 = ((is_padding_reg_444[0:0] == 1'b1) ? 16'd0 : bitcast_ln32_3_fu_403_p1);

assign select_ln33_fu_331_p3 = ((is_padding_reg_444[0:0] == 1'b1) ? 16'd0 : bitcast_ln32_fu_327_p1);

assign sext_ln32_fu_303_p1 = (tmp_1_fu_296_p3);

assign sub_ln32_cast_fu_266_p1 = (sub_ln32_fu_260_p2);

assign sub_ln32_fu_260_p2 = (zext_ln32_1_fu_244_p1 - zext_ln32_5_fu_256_p1);

assign tmp_1_fu_296_p3 = {{add_ln32_reg_454}, {lshr_ln_fu_286_p4}};

assign tmp_4_fu_248_p3 = {{row_coord_int_fu_223_p3}, {1'd0}};

assign tmp_4_i_i_fu_350_p4 = {{in_data_q0[31:16]}};

assign tmp_5_i_i_fu_372_p4 = {{in_data_q0[47:32]}};

assign tmp_6_i_i_fu_393_p4 = {{in_data_q0[63:48]}};

assign tmp_fu_236_p3 = {{row_coord_int_fu_223_p3}, {4'd0}};

assign trunc_ln135_fu_192_p1 = indices_01_dout[3:0];

assign trunc_ln32_fu_323_p1 = in_data_q0[15:0];

assign zext_ln32_1_fu_244_p1 = tmp_fu_236_p3;

assign zext_ln32_2_fu_345_p1 = or_ln25_fu_339_p2;

assign zext_ln32_3_fu_419_p1 = or_ln25_1_fu_414_p2;

assign zext_ln32_4_fu_429_p1 = or_ln25_2_fu_424_p2;

assign zext_ln32_5_fu_256_p1 = tmp_4_fu_248_p3;

assign zext_ln32_6_fu_270_p1 = col_coord_int_fu_229_p3;

assign zext_ln32_fu_318_p1 = kk_0_i_i_reg_180_pp0_iter1_reg;

endmodule //td_fused_top_tdf9_readInputs
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_tdf9_writeOutputs_unaligned (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        indices_01_dout,
        indices_01_empty_n,
        indices_01_read,
        indices_12_dout,
        indices_12_empty_n,
        indices_12_read,
        p_read,
        out_data_address1,
        out_data_ce1,
        out_data_we1,
        out_data_d1
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_state2 = 3'd2;
parameter    ap_ST_fsm_state3 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
input  [3:0] indices_01_dout;
input   indices_01_empty_n;
output   indices_01_read;
input  [7:0] indices_12_dout;
input   indices_12_empty_n;
output   indices_12_read;
input  [15:0] p_read;
output  [11:0] out_data_address1;
output   out_data_ce1;
output   out_data_we1;
output  [63:0] out_data_d1;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg indices_01_read;
reg indices_12_read;
reg out_data_ce1;
reg out_data_we1;

reg    ap_done_reg;
  reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg   [15:0] outputCount;
reg   [15:0] outputChanIdx;
reg   [15:0] outputRow_0;
reg   [15:0] outputRow_1;
reg   [15:0] outputRow_2;
reg   [15:0] outputRow_3;
reg    indices_01_blk_n;
reg    indices_12_blk_n;
wire   [7:0] add_ln94_fu_147_p2;
reg   [7:0] add_ln94_reg_304;
wire   [15:0] add_ln87_fu_192_p2;
wire    ap_CS_fsm_state2;
wire   [0:0] icmp_ln88_fu_198_p2;
reg   [0:0] icmp_ln88_reg_317;
reg   [15:0] ap_phi_mux_empty_phi_fu_114_p4;
reg   [15:0] empty_reg_111;
wire    ap_CS_fsm_state3;
wire   [63:0] zext_ln94_2_fu_226_p1;
wire   [15:0] select_ln97_fu_284_p3;
wire   [1:0] trunc_ln86_fu_164_p1;
reg   [15:0] ap_sig_allocacmp_outputRow_0_load;
reg   [15:0] ap_sig_allocacmp_outputRow_1_load;
reg   [15:0] ap_sig_allocacmp_outputRow_2_load;
reg   [15:0] ap_sig_allocacmp_outputRow_3_load;
reg    ap_block_state1;
wire   [4:0] tmp_1_fu_129_p3;
wire   [7:0] tmp_fu_121_p3;
wire   [7:0] zext_ln94_fu_137_p1;
wire   [7:0] sub_ln94_fu_141_p2;
wire   [5:0] trunc_ln94_fu_212_p1;
wire   [11:0] tmp_3_cast_fu_153_p3;
wire   [11:0] zext_ln94_1_fu_216_p1;
wire   [11:0] add_ln94_1_fu_220_p2;
wire   [15:0] bitcast_ln94_3_fu_255_p1;
wire   [15:0] bitcast_ln94_2_fu_247_p1;
wire   [15:0] bitcast_ln94_1_fu_239_p1;
wire   [15:0] bitcast_ln94_fu_231_p1;
wire   [15:0] add_ln96_fu_272_p2;
wire   [0:0] icmp_ln97_fu_278_p2;
reg   [2:0] ap_NS_fsm;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 3'd1;
#0 outputCount = 16'd0;
#0 outputChanIdx = 16'd0;
#0 outputRow_0 = 16'd0;
#0 outputRow_1 = 16'd0;
#0 outputRow_2 = 16'd0;
#0 outputRow_3 = 16'd0;
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state3)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln88_reg_317 == 1'd1) & (1'b1 == ap_CS_fsm_state3))) begin
        empty_reg_111 <= 16'd0;
    end else if (((icmp_ln88_fu_198_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state2))) begin
        empty_reg_111 <= add_ln87_fu_192_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state1)) begin
        add_ln94_reg_304 <= add_ln94_fu_147_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        icmp_ln88_reg_317 <= icmp_ln88_fu_198_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln88_fu_198_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        outputChanIdx <= select_ln97_fu_284_p3;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state3)) begin
        outputCount <= ap_phi_mux_empty_phi_fu_114_p4;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln86_fu_164_p1 == 2'd0) & (1'b1 == ap_CS_fsm_state2))) begin
        outputRow_0 <= p_read;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln86_fu_164_p1 == 2'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        outputRow_1 <= p_read;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln86_fu_164_p1 == 2'd2) & (1'b1 == ap_CS_fsm_state2))) begin
        outputRow_2 <= p_read;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln86_fu_164_p1 == 2'd3) & (1'b1 == ap_CS_fsm_state2))) begin
        outputRow_3 <= p_read;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state3)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln88_reg_317 == 1'd1) & (1'b1 == ap_CS_fsm_state3))) begin
        ap_phi_mux_empty_phi_fu_114_p4 = 16'd0;
    end else begin
        ap_phi_mux_empty_phi_fu_114_p4 = empty_reg_111;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state3)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((trunc_ln86_fu_164_p1 == 2'd0) & (1'b1 == ap_CS_fsm_state2))) begin
        ap_sig_allocacmp_outputRow_0_load = p_read;
    end else begin
        ap_sig_allocacmp_outputRow_0_load = outputRow_0;
    end
end

always @ (*) begin
    if (((trunc_ln86_fu_164_p1 == 2'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        ap_sig_allocacmp_outputRow_1_load = p_read;
    end else begin
        ap_sig_allocacmp_outputRow_1_load = outputRow_1;
    end
end

always @ (*) begin
    if (((trunc_ln86_fu_164_p1 == 2'd2) & (1'b1 == ap_CS_fsm_state2))) begin
        ap_sig_allocacmp_outputRow_2_load = p_read;
    end else begin
        ap_sig_allocacmp_outputRow_2_load = outputRow_2;
    end
end

always @ (*) begin
    if (((trunc_ln86_fu_164_p1 == 2'd3) & (1'b1 == ap_CS_fsm_state2))) begin
        ap_sig_allocacmp_outputRow_3_load = p_read;
    end else begin
        ap_sig_allocacmp_outputRow_3_load = outputRow_3;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_01_blk_n = indices_01_empty_n;
    end else begin
        indices_01_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_01_read = 1'b1;
    end else begin
        indices_01_read = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_12_blk_n = indices_12_empty_n;
    end else begin
        indices_12_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_start == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indices_12_read = 1'b1;
    end else begin
        indices_12_read = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state2))) begin
        out_data_ce1 = 1'b1;
    end else begin
        out_data_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln88_fu_198_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        out_data_we1 = 1'b1;
    end else begin
        out_data_we1 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_start == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_state2 : begin
            ap_NS_fsm = ap_ST_fsm_state3;
        end
        ap_ST_fsm_state3 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln87_fu_192_p2 = (outputCount + 16'd1);

assign add_ln94_1_fu_220_p2 = (tmp_3_cast_fu_153_p3 + zext_ln94_1_fu_216_p1);

assign add_ln94_fu_147_p2 = (sub_ln94_fu_141_p2 + indices_12_dout);

assign add_ln96_fu_272_p2 = (outputChanIdx + 16'd1);

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (indices_12_empty_n == 1'b0) | (indices_01_empty_n == 1'b0) | (ap_done_reg == 1'b1));
end

assign bitcast_ln94_1_fu_239_p1 = ap_sig_allocacmp_outputRow_1_load;

assign bitcast_ln94_2_fu_247_p1 = ap_sig_allocacmp_outputRow_2_load;

assign bitcast_ln94_3_fu_255_p1 = ap_sig_allocacmp_outputRow_3_load;

assign bitcast_ln94_fu_231_p1 = ap_sig_allocacmp_outputRow_0_load;

assign icmp_ln88_fu_198_p2 = ((add_ln87_fu_192_p2 == 16'd4) ? 1'b1 : 1'b0);

assign icmp_ln97_fu_278_p2 = ((add_ln96_fu_272_p2 == 16'd16) ? 1'b1 : 1'b0);

assign out_data_address1 = zext_ln94_2_fu_226_p1;

assign out_data_d1 = {{{{bitcast_ln94_3_fu_255_p1}, {bitcast_ln94_2_fu_247_p1}}, {bitcast_ln94_1_fu_239_p1}}, {bitcast_ln94_fu_231_p1}};

assign select_ln97_fu_284_p3 = ((icmp_ln97_fu_278_p2[0:0] == 1'b1) ? 16'd0 : add_ln96_fu_272_p2);

assign sub_ln94_fu_141_p2 = (tmp_fu_121_p3 - zext_ln94_fu_137_p1);

assign tmp_1_fu_129_p3 = {{indices_01_dout}, {1'd0}};

assign tmp_3_cast_fu_153_p3 = {{add_ln94_reg_304}, {4'd0}};

assign tmp_fu_121_p3 = {{indices_01_dout}, {4'd0}};

assign trunc_ln86_fu_164_p1 = outputCount[1:0];

assign trunc_ln94_fu_212_p1 = outputChanIdx[5:0];

assign zext_ln94_1_fu_216_p1 = trunc_ln94_fu_212_p1;

assign zext_ln94_2_fu_226_p1 = add_ln94_1_fu_220_p2;

assign zext_ln94_fu_137_p1 = tmp_1_fu_129_p3;

endmodule //td_fused_top_tdf9_writeOutputs_unaligned
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_td_fused_axi_in_p_ram (addr0, ce0, d0, we0, addr1, ce1, q1, addr2, ce2, q2, addr3, ce3, q3, addr4, ce4, q4,  clk);

parameter DWIDTH = 16;
parameter AWIDTH = 2;
parameter MEM_SIZE = 4;

input[AWIDTH-1:0] addr0;
input ce0;
input[DWIDTH-1:0] d0;
input we0;
input[AWIDTH-1:0] addr1;
input ce1;
output reg[DWIDTH-1:0] q1;
input[AWIDTH-1:0] addr2;
input ce2;
output reg[DWIDTH-1:0] q2;
input[AWIDTH-1:0] addr3;
input ce3;
output reg[DWIDTH-1:0] q3;
input[AWIDTH-1:0] addr4;
input ce4;
output reg[DWIDTH-1:0] q4;
input clk;

reg [DWIDTH-1:0] ram0[MEM_SIZE-1:0];
reg [DWIDTH-1:0] ram1[MEM_SIZE-1:0];
reg [DWIDTH-1:0] ram2[MEM_SIZE-1:0];
reg [DWIDTH-1:0] ram3[MEM_SIZE-1:0];



always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram0[addr0] <= d0; 
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        q1 <= ram0[addr1];
    end
end


always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram1[addr0] <= d0; 
    end
end

always @(posedge clk)  
begin 
    if (ce2) begin
        q2 <= ram1[addr2];
    end
end


always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram2[addr0] <= d0; 
    end
end

always @(posedge clk)  
begin 
    if (ce3) begin
        q3 <= ram2[addr3];
    end
end


always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram3[addr0] <= d0; 
    end
end

always @(posedge clk)  
begin 
    if (ce4) begin
        q4 <= ram3[addr4];
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_td_fused_axi_in_p(
    reset,
    clk,
    address0,
    ce0,
    we0,
    d0,
    address1,
    ce1,
    q1,
    address2,
    ce2,
    q2,
    address3,
    ce3,
    q3,
    address4,
    ce4,
    q4);

parameter DataWidth = 32'd16;
parameter AddressRange = 32'd4;
parameter AddressWidth = 32'd2;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
input we0;
input[DataWidth - 1:0] d0;
input[AddressWidth - 1:0] address1;
input ce1;
output[DataWidth - 1:0] q1;
input[AddressWidth - 1:0] address2;
input ce2;
output[DataWidth - 1:0] q2;
input[AddressWidth - 1:0] address3;
input ce3;
output[DataWidth - 1:0] q3;
input[AddressWidth - 1:0] address4;
input ce4;
output[DataWidth - 1:0] q4;



td_fused_top_td_fused_axi_in_p_ram td_fused_top_td_fused_axi_in_p_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .we0( we0 ),
    .d0( d0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .q1( q1 ),
    .addr2( address2 ),
    .ce2( ce2 ),
    .q2( q2 ),
    .addr3( address3 ),
    .ce3( ce3 ),
    .q3( q3 ),
    .addr4( address4 ),
    .ce4( ce4 ),
    .q4( q4 )
);

endmodule

// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_td_fused_axi_in (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        stream_in_TDATA,
        stream_in_TVALID,
        stream_in_TREADY,
        stream_in_TKEEP,
        stream_in_TSTRB,
        stream_in_TLAST,
        fmaps_address1,
        fmaps_ce1,
        fmaps_we1,
        fmaps_d1
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_pp0_stage0 = 3'd2;
parameter    ap_ST_fsm_state6 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
input  [15:0] stream_in_TDATA;
input   stream_in_TVALID;
output   stream_in_TREADY;
input  [1:0] stream_in_TKEEP;
input  [1:0] stream_in_TSTRB;
input  [0:0] stream_in_TLAST;
output  [15:0] fmaps_address1;
output   fmaps_ce1;
output   fmaps_we1;
output  [63:0] fmaps_d1;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg stream_in_TREADY;
reg fmaps_ce1;
reg fmaps_we1;

reg    ap_done_reg;
  reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg   [17:0] indvar_flatten16_reg_185;
reg   [9:0] indvar_flatten_reg_196;
reg   [1:0] ch_reg_207;
reg   [7:0] r_reg_218;
reg   [7:0] c_reg_229;
wire   [17:0] add_ln17_fu_240_p2;
wire    ap_CS_fsm_pp0_stage0;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
wire    ap_block_state4_pp0_stage0_iter2;
wire    ap_block_state5_pp0_stage0_iter3;
wire    ap_block_pp0_stage0_11001;
wire   [0:0] icmp_ln17_fu_246_p2;
reg   [0:0] icmp_ln17_reg_483;
reg   [0:0] icmp_ln17_reg_483_pp0_iter1_reg;
reg   [0:0] icmp_ln17_reg_483_pp0_iter2_reg;
wire   [0:0] icmp_ln18_fu_255_p2;
reg   [0:0] icmp_ln18_reg_487;
reg   [0:0] icmp_ln18_reg_487_pp0_iter1_reg;
wire   [0:0] and_ln22_fu_273_p2;
reg   [0:0] and_ln22_reg_493;
reg   [0:0] and_ln22_reg_493_pp0_iter1_reg;
wire   [0:0] icmp_ln25_fu_319_p2;
reg   [0:0] icmp_ln25_reg_498;
reg   [0:0] icmp_ln25_reg_498_pp0_iter1_reg;
wire   [1:0] add_ln20_fu_330_p2;
wire   [9:0] select_ln18_fu_342_p3;
wire   [15:0] p_q4;
reg   [15:0] p_load_3_reg_512;
reg    ap_enable_reg_pp0_iter1;
wire   [7:0] select_ln22_1_fu_363_p3;
reg   [7:0] select_ln22_1_reg_517;
reg    ap_enable_reg_pp0_iter2;
wire   [7:0] select_ln19_48_fu_402_p3;
reg   [7:0] select_ln19_48_reg_522;
reg    ap_block_state1;
wire    ap_block_pp0_stage0_subdone;
reg    ap_condition_pp0_flush_enable;
reg    ap_condition_pp0_exit_iter2_state4;
reg    ap_enable_reg_pp0_iter3;
wire   [1:0] p_address0;
reg    p_ce0;
reg    p_we0;
wire   [15:0] p_d0;
wire   [1:0] p_address1;
reg    p_ce1;
wire   [15:0] p_q1;
wire   [1:0] p_address2;
reg    p_ce2;
wire   [15:0] p_q2;
wire   [1:0] p_address3;
reg    p_ce3;
wire   [15:0] p_q3;
wire   [1:0] p_address4;
reg    p_ce4;
reg   [7:0] ap_phi_mux_r_phi_fu_222_p4;
wire    ap_block_pp0_stage0;
reg   [7:0] ap_phi_mux_c_phi_fu_233_p4;
wire   [63:0] zext_ln20_fu_293_p1;
wire   [63:0] zext_ln27_2_fu_419_p1;
reg   [15:0] tmp_data_1_fu_88;
wire   [15:0] tmp_data_fu_310_p3;
wire   [0:0] empty_154_nbread_fu_96_p5_0;
wire   [0:0] icmp_ln20_fu_267_p2;
wire   [0:0] xor_ln22_fu_261_p2;
wire   [0:0] or_ln19_fu_279_p2;
wire   [1:0] select_ln19_fu_285_p3;
wire   [15:0] tmp_data_2_fu_306_p1;
wire   [9:0] add_ln18_2_fu_336_p2;
wire   [7:0] r_2_fu_350_p2;
wire   [12:0] tmp_22_fu_378_p3;
wire   [15:0] tmp_fu_370_p3;
wire   [15:0] zext_ln27_fu_386_p1;
wire   [7:0] select_ln22_fu_356_p3;
wire   [7:0] c_2_fu_396_p2;
wire   [15:0] sub_ln27_fu_390_p2;
wire   [15:0] zext_ln27_1_fu_409_p1;
wire   [15:0] add_ln27_fu_413_p2;
wire   [15:0] bitcast_ln27_3_fu_436_p1;
wire   [15:0] bitcast_ln27_2_fu_432_p1;
wire   [15:0] bitcast_ln27_1_fu_428_p1;
wire   [15:0] bitcast_ln27_fu_424_p1;
wire    ap_CS_fsm_state6;
reg   [2:0] ap_NS_fsm;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
end

td_fused_top_td_fused_axi_in_p #(
    .DataWidth( 16 ),
    .AddressRange( 4 ),
    .AddressWidth( 2 ))
p_U(
    .reset(ap_rst),
    .clk(ap_clk),
    .address0(p_address0),
    .ce0(p_ce0),
    .we0(p_we0),
    .d0(p_d0),
    .address1(p_address1),
    .ce1(p_ce1),
    .q1(p_q1),
    .address2(p_address2),
    .ce2(p_ce2),
    .q2(p_q2),
    .address3(p_address3),
    .ce3(p_ce3),
    .q3(p_q3),
    .address4(p_address4),
    .ce4(p_ce4),
    .q4(p_q4)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state6)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if ((1'b1 == ap_condition_pp0_flush_enable)) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end else if ((((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_condition_pp0_exit_iter2_state4) & (ap_enable_reg_pp0_iter1 == 1'b0)) | (~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1)))) begin
            ap_enable_reg_pp0_iter2 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_condition_pp0_exit_iter2_state4))) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter1;
        end else if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter3 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln17_reg_483_pp0_iter2_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter3 == 1'b1))) begin
        c_reg_229 <= select_ln19_48_reg_522;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        c_reg_229 <= 8'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln17_fu_246_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ch_reg_207 <= add_ln20_fu_330_p2;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        ch_reg_207 <= 2'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln17_fu_246_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        indvar_flatten16_reg_185 <= add_ln17_fu_240_p2;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indvar_flatten16_reg_185 <= 18'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln17_fu_246_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        indvar_flatten_reg_196 <= select_ln18_fu_342_p3;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        indvar_flatten_reg_196 <= 10'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln17_reg_483_pp0_iter2_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter3 == 1'b1))) begin
        r_reg_218 <= select_ln22_1_reg_517;
    end else if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
        r_reg_218 <= 8'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln17_fu_246_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        and_ln22_reg_493 <= and_ln22_fu_273_p2;
        icmp_ln18_reg_487 <= icmp_ln18_fu_255_p2;
        icmp_ln25_reg_498 <= icmp_ln25_fu_319_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        and_ln22_reg_493_pp0_iter1_reg <= and_ln22_reg_493;
        icmp_ln17_reg_483 <= icmp_ln17_fu_246_p2;
        icmp_ln17_reg_483_pp0_iter1_reg <= icmp_ln17_reg_483;
        icmp_ln18_reg_487_pp0_iter1_reg <= icmp_ln18_reg_487;
        icmp_ln25_reg_498_pp0_iter1_reg <= icmp_ln25_reg_498;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        icmp_ln17_reg_483_pp0_iter2_reg <= icmp_ln17_reg_483_pp0_iter1_reg;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln25_reg_498 == 1'd1) & (icmp_ln17_reg_483 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        p_load_3_reg_512 <= p_q4;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln17_reg_483_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        select_ln19_48_reg_522 <= select_ln19_48_fu_402_p3;
        select_ln22_1_reg_517 <= select_ln22_1_fu_363_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln17_fu_246_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        tmp_data_1_fu_88 <= tmp_data_fu_310_p3;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
        ap_condition_pp0_exit_iter2_state4 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter2_state4 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln17_fu_246_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_condition_pp0_flush_enable = 1'b1;
    end else begin
        ap_condition_pp0_flush_enable = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state6)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln17_reg_483_pp0_iter2_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter3 == 1'b1))) begin
        ap_phi_mux_c_phi_fu_233_p4 = select_ln19_48_reg_522;
    end else begin
        ap_phi_mux_c_phi_fu_233_p4 = c_reg_229;
    end
end

always @ (*) begin
    if (((icmp_ln17_reg_483_pp0_iter2_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter3 == 1'b1))) begin
        ap_phi_mux_r_phi_fu_222_p4 = select_ln22_1_reg_517;
    end else begin
        ap_phi_mux_r_phi_fu_222_p4 = r_reg_218;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state6)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter3 == 1'b1)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1)))) begin
        fmaps_ce1 = 1'b1;
    end else begin
        fmaps_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln25_reg_498_pp0_iter1_reg == 1'd1) & (icmp_ln17_reg_483_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        fmaps_we1 = 1'b1;
    end else begin
        fmaps_we1 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        p_ce0 = 1'b1;
    end else begin
        p_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        p_ce1 = 1'b1;
    end else begin
        p_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        p_ce2 = 1'b1;
    end else begin
        p_ce2 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
        p_ce3 = 1'b1;
    end else begin
        p_ce3 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        p_ce4 = 1'b1;
    end else begin
        p_ce4 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln17_fu_246_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        p_we0 = 1'b1;
    end else begin
        p_we0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln17_fu_246_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (stream_in_TVALID == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        stream_in_TREADY = 1'b1;
    end else begin
        stream_in_TREADY = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_start == 1'b0) | (ap_done_reg == 1'b1)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if (~((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter2 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter2 == 1'b1) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
                ap_NS_fsm = ap_ST_fsm_state6;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_state6 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln17_fu_240_p2 = (indvar_flatten16_reg_185 + 18'd1);

assign add_ln18_2_fu_336_p2 = (indvar_flatten_reg_196 + 10'd1);

assign add_ln20_fu_330_p2 = (select_ln19_fu_285_p3 + 2'd1);

assign add_ln27_fu_413_p2 = (sub_ln27_fu_390_p2 + zext_ln27_1_fu_409_p1);

assign and_ln22_fu_273_p2 = (xor_ln22_fu_261_p2 & icmp_ln20_fu_267_p2);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state6 = ap_CS_fsm[32'd2];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state1 = ((ap_start == 1'b0) | (ap_done_reg == 1'b1));
end

assign ap_block_state2_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign bitcast_ln27_1_fu_428_p1 = p_q2;

assign bitcast_ln27_2_fu_432_p1 = p_q1;

assign bitcast_ln27_3_fu_436_p1 = p_load_3_reg_512;

assign bitcast_ln27_fu_424_p1 = p_q3;

assign c_2_fu_396_p2 = (select_ln22_fu_356_p3 + 8'd1);

assign empty_154_nbread_fu_96_p5_0 = stream_in_TVALID;

assign fmaps_address1 = zext_ln27_2_fu_419_p1;

assign fmaps_d1 = {{{{bitcast_ln27_3_fu_436_p1}, {bitcast_ln27_2_fu_432_p1}}, {bitcast_ln27_1_fu_428_p1}}, {bitcast_ln27_fu_424_p1}};

assign icmp_ln17_fu_246_p2 = ((indvar_flatten16_reg_185 == 18'd150528) ? 1'b1 : 1'b0);

assign icmp_ln18_fu_255_p2 = ((indvar_flatten_reg_196 == 10'd672) ? 1'b1 : 1'b0);

assign icmp_ln20_fu_267_p2 = ((ch_reg_207 == 2'd3) ? 1'b1 : 1'b0);

assign icmp_ln25_fu_319_p2 = ((select_ln19_fu_285_p3 == 2'd2) ? 1'b1 : 1'b0);

assign or_ln19_fu_279_p2 = (icmp_ln18_fu_255_p2 | and_ln22_fu_273_p2);

assign p_address0 = zext_ln20_fu_293_p1;

assign p_address1 = 64'd2;

assign p_address2 = 64'd1;

assign p_address3 = 64'd0;

assign p_address4 = 64'd3;

assign p_d0 = ((empty_154_nbread_fu_96_p5_0[0:0] == 1'b1) ? tmp_data_2_fu_306_p1 : tmp_data_1_fu_88);

assign r_2_fu_350_p2 = (ap_phi_mux_r_phi_fu_222_p4 + 8'd1);

assign select_ln18_fu_342_p3 = ((icmp_ln18_fu_255_p2[0:0] == 1'b1) ? 10'd1 : add_ln18_2_fu_336_p2);

assign select_ln19_48_fu_402_p3 = ((and_ln22_reg_493_pp0_iter1_reg[0:0] == 1'b1) ? c_2_fu_396_p2 : select_ln22_fu_356_p3);

assign select_ln19_fu_285_p3 = ((or_ln19_fu_279_p2[0:0] == 1'b1) ? 2'd0 : ch_reg_207);

assign select_ln22_1_fu_363_p3 = ((icmp_ln18_reg_487_pp0_iter1_reg[0:0] == 1'b1) ? r_2_fu_350_p2 : ap_phi_mux_r_phi_fu_222_p4);

assign select_ln22_fu_356_p3 = ((icmp_ln18_reg_487_pp0_iter1_reg[0:0] == 1'b1) ? 8'd0 : ap_phi_mux_c_phi_fu_233_p4);

assign sub_ln27_fu_390_p2 = (tmp_fu_370_p3 - zext_ln27_fu_386_p1);

assign tmp_22_fu_378_p3 = {{select_ln22_1_fu_363_p3}, {5'd0}};

assign tmp_data_2_fu_306_p1 = stream_in_TDATA;

assign tmp_data_fu_310_p3 = ((empty_154_nbread_fu_96_p5_0[0:0] == 1'b1) ? tmp_data_2_fu_306_p1 : tmp_data_1_fu_88);

assign tmp_fu_370_p3 = {{select_ln22_1_fu_363_p3}, {8'd0}};

assign xor_ln22_fu_261_p2 = (icmp_ln18_fu_255_p2 ^ 1'd1);

assign zext_ln20_fu_293_p1 = select_ln19_fu_285_p3;

assign zext_ln27_1_fu_409_p1 = select_ln19_48_fu_402_p3;

assign zext_ln27_2_fu_419_p1 = add_ln27_fu_413_p2;

assign zext_ln27_fu_386_p1 = tmp_22_fu_378_p3;

endmodule //td_fused_top_td_fused_axi_in
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_td_fused_axi_out (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        fmaps_address0,
        fmaps_ce0,
        fmaps_q0,
        stream_out_TDATA,
        stream_out_TVALID,
        stream_out_TREADY,
        stream_out_TKEEP,
        stream_out_TSTRB,
        stream_out_TLAST
);

parameter    ap_ST_fsm_state1 = 6'd1;
parameter    ap_ST_fsm_pp0_stage0 = 6'd2;
parameter    ap_ST_fsm_pp0_stage1 = 6'd4;
parameter    ap_ST_fsm_pp0_stage2 = 6'd8;
parameter    ap_ST_fsm_pp0_stage3 = 6'd16;
parameter    ap_ST_fsm_state13 = 6'd32;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
output  [15:0] fmaps_address0;
output   fmaps_ce0;
input  [63:0] fmaps_q0;
output  [15:0] stream_out_TDATA;
output   stream_out_TVALID;
input   stream_out_TREADY;
output  [1:0] stream_out_TKEEP;
output  [1:0] stream_out_TSTRB;
output  [0:0] stream_out_TLAST;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg fmaps_ce0;
reg[15:0] stream_out_TDATA;
reg stream_out_TVALID;

reg    ap_done_reg;
  reg   [5:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    stream_out_TDATA_blk_n;
wire    ap_CS_fsm_pp0_stage3;
reg    ap_enable_reg_pp0_iter1;
wire    ap_block_pp0_stage3;
reg   [0:0] icmp_ln17_reg_400;
reg   [0:0] icmp_ln17_reg_400_pp0_iter1_reg;
wire    ap_CS_fsm_pp0_stage0;
reg    ap_enable_reg_pp0_iter2;
wire    ap_block_pp0_stage0;
wire    ap_CS_fsm_pp0_stage1;
wire    ap_block_pp0_stage1;
reg   [0:0] icmp_ln17_reg_400_pp0_iter2_reg;
wire    ap_CS_fsm_pp0_stage2;
wire    ap_block_pp0_stage2;
reg   [15:0] indvar_flatten13_reg_134;
reg   [3:0] r_reg_145;
reg   [11:0] indvar_flatten_reg_156;
reg   [3:0] c_reg_167;
reg   [9:0] phi_ln25_reg_178;
wire   [15:0] add_ln17_1_fu_189_p2;
reg   [15:0] add_ln17_1_reg_395;
reg    ap_enable_reg_pp0_iter0;
wire    ap_block_state2_pp0_stage0_iter0;
wire    ap_block_state6_pp0_stage0_iter1;
reg    ap_block_state10_pp0_stage0_iter2;
reg    ap_block_state10_io;
reg    ap_block_pp0_stage0_11001;
wire   [0:0] icmp_ln17_fu_195_p2;
wire   [0:0] icmp_ln18_fu_207_p2;
reg   [0:0] icmp_ln18_reg_404;
wire   [3:0] select_ln17_fu_213_p3;
reg   [3:0] select_ln17_reg_411;
wire   [3:0] select_ln17_1_fu_221_p3;
reg   [3:0] select_ln17_1_reg_417;
wire   [11:0] add_ln18_1_fu_229_p2;
reg   [11:0] add_ln18_1_reg_424;
wire   [9:0] select_ln18_fu_294_p3;
reg   [9:0] select_ln18_reg_429;
wire    ap_block_state3_pp0_stage1_iter0;
wire    ap_block_state7_pp0_stage1_iter1;
reg    ap_block_state11_pp0_stage1_iter2;
reg    ap_block_state11_io;
reg    ap_block_pp0_stage1_11001;
wire   [3:0] select_ln18_1_fu_302_p3;
reg   [3:0] select_ln18_1_reg_434;
reg   [7:0] lshr_ln_reg_444;
wire   [11:0] select_ln18_2_fu_333_p3;
reg   [11:0] select_ln18_2_reg_449;
wire    ap_block_state5_pp0_stage3_iter0;
reg    ap_block_state9_pp0_stage3_iter1;
reg    ap_block_state9_io;
reg    ap_block_pp0_stage3_11001;
wire   [9:0] add_ln19_fu_346_p2;
reg   [9:0] add_ln19_reg_464;
reg   [15:0] tmp_s_reg_469;
reg   [15:0] tmp_1_reg_474;
reg   [15:0] tmp_2_reg_479;
reg    ap_block_state1;
reg    ap_block_pp0_stage1_subdone;
reg    ap_condition_pp0_exit_iter0_state3;
reg    ap_block_pp0_stage3_subdone;
wire    ap_block_state4_pp0_stage2_iter0;
wire    ap_block_state8_pp0_stage2_iter1;
reg    ap_block_state12_pp0_stage2_iter2;
reg    ap_block_state12_io;
reg    ap_block_pp0_stage2_subdone;
reg   [15:0] ap_phi_mux_indvar_flatten13_phi_fu_138_p4;
reg   [3:0] ap_phi_mux_r_phi_fu_149_p4;
reg   [11:0] ap_phi_mux_indvar_flatten_phi_fu_160_p4;
reg   [3:0] ap_phi_mux_c_phi_fu_171_p4;
reg   [9:0] ap_phi_mux_phi_ln25_phi_fu_182_p4;
wire   [63:0] zext_ln25_4_fu_342_p1;
wire   [15:0] trunc_ln25_fu_351_p1;
reg    ap_block_pp0_stage3_01001;
reg    ap_block_pp0_stage0_01001;
reg    ap_block_pp0_stage1_01001;
reg    ap_block_pp0_stage2_01001;
reg    ap_block_pp0_stage2_11001;
wire   [3:0] add_ln17_fu_201_p2;
wire   [7:0] tmp_20_fu_235_p3;
wire   [4:0] tmp_21_fu_246_p3;
wire   [8:0] zext_ln25_fu_242_p1;
wire   [8:0] zext_ln25_1_fu_253_p1;
wire   [8:0] sub_ln25_fu_257_p2;
wire   [0:0] icmp_ln19_fu_272_p2;
wire   [0:0] xor_ln17_fu_267_p2;
wire   [0:0] and_ln17_fu_278_p2;
wire   [0:0] or_ln18_fu_289_p2;
wire   [3:0] add_ln18_fu_284_p2;
wire   [9:0] sext_ln18_fu_263_p1;
wire   [9:0] zext_ln25_2_fu_309_p1;
wire   [9:0] add_ln25_fu_313_p2;
wire   [15:0] grp_fu_386_p3;
wire   [8:0] grp_fu_386_p1;
wire   [7:0] grp_fu_386_p2;
reg    grp_fu_386_ce;
wire    ap_CS_fsm_state13;
reg   [5:0] ap_NS_fsm;
reg    ap_block_pp0_stage0_subdone;
reg    ap_idle_pp0;
wire    ap_enable_pp0;
wire   [15:0] grp_fu_386_p20;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 6'd1;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter0 = 1'b0;
end

td_fused_top_mac_muladd_10s_9ns_8ns_16_4_1 #(
    .ID( 1 ),
    .NUM_STAGE( 4 ),
    .din0_WIDTH( 10 ),
    .din1_WIDTH( 9 ),
    .din2_WIDTH( 8 ),
    .dout_WIDTH( 16 ))
mac_muladd_10s_9ns_8ns_16_4_1_U817(
    .clk(ap_clk),
    .reset(ap_rst),
    .ce(grp_fu_386_ce),
    .din0(add_ln25_fu_313_p2),
    .din1(grp_fu_386_p1),
    .din2(grp_fu_386_p2),
    .dout(grp_fu_386_p3)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if ((1'b1 == ap_CS_fsm_state13)) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1) & (1'b1 == ap_condition_pp0_exit_iter0_state3))) begin
            ap_enable_reg_pp0_iter0 <= 1'b0;
        end else if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter0 <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage3_subdone) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
            ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((((1'b0 == ap_block_pp0_stage2_subdone) & (ap_enable_reg_pp0_iter1 == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage2)) | ((1'b0 == ap_block_pp0_stage3_subdone) & (1'b1 == ap_CS_fsm_pp0_stage3)))) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end else if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
            ap_enable_reg_pp0_iter2 <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln17_reg_400 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        c_reg_167 <= select_ln18_1_reg_434;
    end else if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        c_reg_167 <= 4'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln17_reg_400 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        indvar_flatten13_reg_134 <= add_ln17_1_reg_395;
    end else if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indvar_flatten13_reg_134 <= 16'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln17_reg_400 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        indvar_flatten_reg_156 <= select_ln18_2_reg_449;
    end else if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        indvar_flatten_reg_156 <= 12'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln17_reg_400_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
        phi_ln25_reg_178 <= add_ln19_reg_464;
    end else if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        phi_ln25_reg_178 <= 10'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln17_reg_400 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        r_reg_145 <= select_ln17_1_reg_417;
    end else if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        r_reg_145 <= 4'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
        add_ln17_1_reg_395 <= add_ln17_1_fu_189_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (icmp_ln17_fu_195_p2 == 1'd0))) begin
        add_ln18_1_reg_424 <= add_ln18_1_fu_229_p2;
        icmp_ln18_reg_404 <= icmp_ln18_fu_207_p2;
        select_ln17_reg_411 <= select_ln17_fu_213_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln17_reg_400 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        add_ln19_reg_464 <= add_ln19_fu_346_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln17_reg_400 <= icmp_ln17_fu_195_p2;
        icmp_ln17_reg_400_pp0_iter1_reg <= icmp_ln17_reg_400;
        icmp_ln17_reg_400_pp0_iter2_reg <= icmp_ln17_reg_400_pp0_iter1_reg;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln17_reg_400 == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
        lshr_ln_reg_444 <= {{select_ln18_fu_294_p3[9:2]}};
        select_ln18_reg_429 <= select_ln18_fu_294_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (icmp_ln17_fu_195_p2 == 1'd0) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
        select_ln17_1_reg_417 <= select_ln17_1_fu_221_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln17_reg_400 == 1'd0) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
        select_ln18_1_reg_434 <= select_ln18_1_fu_302_p3;
        select_ln18_2_reg_449 <= select_ln18_2_fu_333_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln17_reg_400_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage3_11001) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
        tmp_1_reg_474 <= {{fmaps_q0[47:32]}};
        tmp_2_reg_479 <= {{fmaps_q0[63:48]}};
        tmp_s_reg_469 <= {{fmaps_q0[31:16]}};
    end
end

always @ (*) begin
    if ((icmp_ln17_reg_400 == 1'd1)) begin
        ap_condition_pp0_exit_iter0_state3 = 1'b1;
    end else begin
        ap_condition_pp0_exit_iter0_state3 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state13)) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln17_reg_400 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_phi_mux_c_phi_fu_171_p4 = select_ln18_1_reg_434;
    end else begin
        ap_phi_mux_c_phi_fu_171_p4 = c_reg_167;
    end
end

always @ (*) begin
    if (((icmp_ln17_reg_400 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_phi_mux_indvar_flatten13_phi_fu_138_p4 = add_ln17_1_reg_395;
    end else begin
        ap_phi_mux_indvar_flatten13_phi_fu_138_p4 = indvar_flatten13_reg_134;
    end
end

always @ (*) begin
    if (((icmp_ln17_reg_400 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_phi_mux_indvar_flatten_phi_fu_160_p4 = select_ln18_2_reg_449;
    end else begin
        ap_phi_mux_indvar_flatten_phi_fu_160_p4 = indvar_flatten_reg_156;
    end
end

always @ (*) begin
    if (((icmp_ln17_reg_400_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
        ap_phi_mux_phi_ln25_phi_fu_182_p4 = add_ln19_reg_464;
    end else begin
        ap_phi_mux_phi_ln25_phi_fu_182_p4 = phi_ln25_reg_178;
    end
end

always @ (*) begin
    if (((icmp_ln17_reg_400 == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_phi_mux_r_phi_fu_149_p4 = select_ln17_1_reg_417;
    end else begin
        ap_phi_mux_r_phi_fu_149_p4 = r_reg_145;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state13)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage2_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2)) | ((1'b0 == ap_block_pp0_stage3_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)) | ((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
        fmaps_ce0 = 1'b1;
    end else begin
        fmaps_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage2_11001) & (1'b1 == ap_CS_fsm_pp0_stage2)) | ((1'b0 == ap_block_pp0_stage3_11001) & (1'b1 == ap_CS_fsm_pp0_stage3)) | ((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1)) | ((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
        grp_fu_386_ce = 1'b1;
    end else begin
        grp_fu_386_ce = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln17_reg_400_pp0_iter2_reg == 1'd0) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage2_01001) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
        stream_out_TDATA = tmp_2_reg_479;
    end else if (((icmp_ln17_reg_400_pp0_iter2_reg == 1'd0) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage1_01001) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
        stream_out_TDATA = tmp_1_reg_474;
    end else if (((ap_enable_reg_pp0_iter2 == 1'b1) & (icmp_ln17_reg_400_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_01001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        stream_out_TDATA = tmp_s_reg_469;
    end else if (((icmp_ln17_reg_400_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage3_01001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3))) begin
        stream_out_TDATA = trunc_ln25_fu_351_p1;
    end else begin
        stream_out_TDATA = 'bx;
    end
end

always @ (*) begin
    if ((((icmp_ln17_reg_400_pp0_iter2_reg == 1'd0) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2)) | ((icmp_ln17_reg_400_pp0_iter2_reg == 1'd0) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1)) | ((ap_enable_reg_pp0_iter2 == 1'b1) & (icmp_ln17_reg_400_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((icmp_ln17_reg_400_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage3) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)))) begin
        stream_out_TDATA_blk_n = stream_out_TREADY;
    end else begin
        stream_out_TDATA_blk_n = 1'b1;
    end
end

always @ (*) begin
    if ((((icmp_ln17_reg_400_pp0_iter2_reg == 1'd0) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage2_11001) & (1'b1 == ap_CS_fsm_pp0_stage2)) | ((icmp_ln17_reg_400_pp0_iter2_reg == 1'd0) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1)) | ((ap_enable_reg_pp0_iter2 == 1'b1) & (icmp_ln17_reg_400_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((icmp_ln17_reg_400_pp0_iter1_reg == 1'd0) & (1'b0 == ap_block_pp0_stage3_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage3)))) begin
        stream_out_TVALID = 1'b1;
    end else begin
        stream_out_TVALID = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_pp0_stage0 : begin
            if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_pp0_stage1 : begin
            if ((~((icmp_ln17_reg_400 == 1'd1) & (1'b0 == ap_block_pp0_stage1_subdone) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1)) & (1'b0 == ap_block_pp0_stage1_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage2;
            end else if (((icmp_ln17_reg_400 == 1'd1) & (1'b0 == ap_block_pp0_stage1_subdone) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
                ap_NS_fsm = ap_ST_fsm_state13;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end
        end
        ap_ST_fsm_pp0_stage2 : begin
            if ((~((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage2_subdone) & (ap_enable_reg_pp0_iter1 == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage2)) & (1'b0 == ap_block_pp0_stage2_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage3;
            end else if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage2_subdone) & (ap_enable_reg_pp0_iter1 == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
                ap_NS_fsm = ap_ST_fsm_state13;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage2;
            end
        end
        ap_ST_fsm_pp0_stage3 : begin
            if ((1'b0 == ap_block_pp0_stage3_subdone)) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage3;
            end
        end
        ap_ST_fsm_state13 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln17_1_fu_189_p2 = (ap_phi_mux_indvar_flatten13_phi_fu_138_p4 + 16'd1);

assign add_ln17_fu_201_p2 = (ap_phi_mux_r_phi_fu_149_p4 + 4'd1);

assign add_ln18_1_fu_229_p2 = (ap_phi_mux_indvar_flatten_phi_fu_160_p4 + 12'd1);

assign add_ln18_fu_284_p2 = (select_ln17_reg_411 + 4'd1);

assign add_ln19_fu_346_p2 = (select_ln18_reg_429 + 10'd4);

assign add_ln25_fu_313_p2 = ((sext_ln18_fu_263_p1) + (zext_ln25_2_fu_309_p1));

assign and_ln17_fu_278_p2 = (xor_ln17_fu_267_p2 & icmp_ln19_fu_272_p2);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_pp0_stage1 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_pp0_stage2 = ap_CS_fsm[32'd3];

assign ap_CS_fsm_pp0_stage3 = ap_CS_fsm[32'd4];

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state13 = ap_CS_fsm[32'd5];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_pp0_stage0_01001 = ((ap_enable_reg_pp0_iter2 == 1'b1) & (icmp_ln17_reg_400_pp0_iter1_reg == 1'd0) & (stream_out_TREADY == 1'b0));
end

always @ (*) begin
    ap_block_pp0_stage0_11001 = ((ap_enable_reg_pp0_iter2 == 1'b1) & ((1'b1 == ap_block_state10_io) | ((icmp_ln17_reg_400_pp0_iter1_reg == 1'd0) & (stream_out_TREADY == 1'b0))));
end

always @ (*) begin
    ap_block_pp0_stage0_subdone = ((ap_enable_reg_pp0_iter2 == 1'b1) & ((1'b1 == ap_block_state10_io) | ((icmp_ln17_reg_400_pp0_iter1_reg == 1'd0) & (stream_out_TREADY == 1'b0))));
end

assign ap_block_pp0_stage1 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_pp0_stage1_01001 = ((icmp_ln17_reg_400_pp0_iter2_reg == 1'd0) & (ap_enable_reg_pp0_iter2 == 1'b1) & (stream_out_TREADY == 1'b0));
end

always @ (*) begin
    ap_block_pp0_stage1_11001 = ((ap_enable_reg_pp0_iter2 == 1'b1) & ((1'b1 == ap_block_state11_io) | ((icmp_ln17_reg_400_pp0_iter2_reg == 1'd0) & (stream_out_TREADY == 1'b0))));
end

always @ (*) begin
    ap_block_pp0_stage1_subdone = ((ap_enable_reg_pp0_iter2 == 1'b1) & ((1'b1 == ap_block_state11_io) | ((icmp_ln17_reg_400_pp0_iter2_reg == 1'd0) & (stream_out_TREADY == 1'b0))));
end

assign ap_block_pp0_stage2 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_pp0_stage2_01001 = ((icmp_ln17_reg_400_pp0_iter2_reg == 1'd0) & (ap_enable_reg_pp0_iter2 == 1'b1) & (stream_out_TREADY == 1'b0));
end

always @ (*) begin
    ap_block_pp0_stage2_11001 = ((ap_enable_reg_pp0_iter2 == 1'b1) & ((1'b1 == ap_block_state12_io) | ((icmp_ln17_reg_400_pp0_iter2_reg == 1'd0) & (stream_out_TREADY == 1'b0))));
end

always @ (*) begin
    ap_block_pp0_stage2_subdone = ((ap_enable_reg_pp0_iter2 == 1'b1) & ((1'b1 == ap_block_state12_io) | ((icmp_ln17_reg_400_pp0_iter2_reg == 1'd0) & (stream_out_TREADY == 1'b0))));
end

assign ap_block_pp0_stage3 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_pp0_stage3_01001 = ((icmp_ln17_reg_400_pp0_iter1_reg == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (stream_out_TREADY == 1'b0));
end

always @ (*) begin
    ap_block_pp0_stage3_11001 = ((ap_enable_reg_pp0_iter1 == 1'b1) & ((1'b1 == ap_block_state9_io) | ((icmp_ln17_reg_400_pp0_iter1_reg == 1'd0) & (stream_out_TREADY == 1'b0))));
end

always @ (*) begin
    ap_block_pp0_stage3_subdone = ((ap_enable_reg_pp0_iter1 == 1'b1) & ((1'b1 == ap_block_state9_io) | ((icmp_ln17_reg_400_pp0_iter1_reg == 1'd0) & (stream_out_TREADY == 1'b0))));
end

always @ (*) begin
    ap_block_state1 = ((ap_done_reg == 1'b1) | (ap_start == 1'b0));
end

always @ (*) begin
    ap_block_state10_io = ((icmp_ln17_reg_400_pp0_iter1_reg == 1'd0) & (stream_out_TREADY == 1'b0));
end

always @ (*) begin
    ap_block_state10_pp0_stage0_iter2 = ((icmp_ln17_reg_400_pp0_iter1_reg == 1'd0) & (stream_out_TREADY == 1'b0));
end

always @ (*) begin
    ap_block_state11_io = ((icmp_ln17_reg_400_pp0_iter2_reg == 1'd0) & (stream_out_TREADY == 1'b0));
end

always @ (*) begin
    ap_block_state11_pp0_stage1_iter2 = ((icmp_ln17_reg_400_pp0_iter2_reg == 1'd0) & (stream_out_TREADY == 1'b0));
end

always @ (*) begin
    ap_block_state12_io = ((icmp_ln17_reg_400_pp0_iter2_reg == 1'd0) & (stream_out_TREADY == 1'b0));
end

always @ (*) begin
    ap_block_state12_pp0_stage2_iter2 = ((icmp_ln17_reg_400_pp0_iter2_reg == 1'd0) & (stream_out_TREADY == 1'b0));
end

assign ap_block_state2_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage1_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage2_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage3_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage1_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage2_iter1 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state9_io = ((icmp_ln17_reg_400_pp0_iter1_reg == 1'd0) & (stream_out_TREADY == 1'b0));
end

always @ (*) begin
    ap_block_state9_pp0_stage3_iter1 = ((icmp_ln17_reg_400_pp0_iter1_reg == 1'd0) & (stream_out_TREADY == 1'b0));
end

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign fmaps_address0 = zext_ln25_4_fu_342_p1;

assign grp_fu_386_p1 = 16'd250;

assign grp_fu_386_p2 = grp_fu_386_p20;

assign grp_fu_386_p20 = lshr_ln_reg_444;

assign icmp_ln17_fu_195_p2 = ((ap_phi_mux_indvar_flatten13_phi_fu_138_p4 == 16'd49000) ? 1'b1 : 1'b0);

assign icmp_ln18_fu_207_p2 = ((ap_phi_mux_indvar_flatten_phi_fu_160_p4 == 12'd3500) ? 1'b1 : 1'b0);

assign icmp_ln19_fu_272_p2 = ((ap_phi_mux_phi_ln25_phi_fu_182_p4 == 10'd1000) ? 1'b1 : 1'b0);

assign or_ln18_fu_289_p2 = (icmp_ln18_reg_404 | and_ln17_fu_278_p2);

assign select_ln17_1_fu_221_p3 = ((icmp_ln18_fu_207_p2[0:0] == 1'b1) ? add_ln17_fu_201_p2 : ap_phi_mux_r_phi_fu_149_p4);

assign select_ln17_fu_213_p3 = ((icmp_ln18_fu_207_p2[0:0] == 1'b1) ? 4'd0 : ap_phi_mux_c_phi_fu_171_p4);

assign select_ln18_1_fu_302_p3 = ((and_ln17_fu_278_p2[0:0] == 1'b1) ? add_ln18_fu_284_p2 : select_ln17_reg_411);

assign select_ln18_2_fu_333_p3 = ((icmp_ln18_reg_404[0:0] == 1'b1) ? 12'd1 : add_ln18_1_reg_424);

assign select_ln18_fu_294_p3 = ((or_ln18_fu_289_p2[0:0] == 1'b1) ? 10'd0 : ap_phi_mux_phi_ln25_phi_fu_182_p4);

assign sext_ln18_fu_263_p1 = (sub_ln25_fu_257_p2);

assign stream_out_TKEEP = 2'd0;

assign stream_out_TLAST = 1'd0;

assign stream_out_TSTRB = 2'd0;

assign sub_ln25_fu_257_p2 = (zext_ln25_fu_242_p1 - zext_ln25_1_fu_253_p1);

assign tmp_20_fu_235_p3 = {{select_ln17_1_reg_417}, {4'd0}};

assign tmp_21_fu_246_p3 = {{select_ln17_1_reg_417}, {1'd0}};

assign trunc_ln25_fu_351_p1 = fmaps_q0[15:0];

assign xor_ln17_fu_267_p2 = (icmp_ln18_reg_404 ^ 1'd1);

assign zext_ln25_1_fu_253_p1 = tmp_21_fu_246_p3;

assign zext_ln25_2_fu_309_p1 = select_ln18_1_fu_302_p3;

assign zext_ln25_4_fu_342_p1 = (grp_fu_386_p3);

assign zext_ln25_fu_242_p1 = tmp_20_fu_235_p3;

endmodule //td_fused_top_td_fused_axi_out
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_td_fused_final_fmaps_memcore_ram (addr0, ce0, q0, addr1, ce1, d1, we1,  clk);

parameter DWIDTH = 64;
parameter AWIDTH = 16;
parameter MEM_SIZE = 49000;

input[AWIDTH-1:0] addr0;
input ce0;
output wire[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
input clk;

 reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];
wire [AWIDTH-1:0] addr0_t0; 
reg [AWIDTH-1:0] addr0_t1; 
reg [DWIDTH-1:0] q0_t0;
  reg [DWIDTH-1:0] q0_t1;
wire [AWIDTH-1:0] addr1_t0; 
reg [AWIDTH-1:0] addr1_t1; 
wire [DWIDTH-1:0] d1_t0; 
wire we1_t0; 
reg [DWIDTH-1:0] d1_t1; 
reg we1_t1; 


assign addr0_t0 = addr0;
assign q0 = q0_t1;
assign addr1_t0 = addr1;
assign d1_t0 = d1;
assign we1_t0 = we1;

always @(posedge clk)  
begin
    if (ce0) 
    begin
        addr0_t1 <= addr0_t0; 
        q0_t1 <= q0_t0;
    end
    if (ce1) 
    begin
        addr1_t1 <= addr1_t0; 
        d1_t1 <= d1_t0;
        we1_t1 <= we1_t0;
    end
end


always @(posedge clk)  
begin 
    if (ce0) begin
        q0_t0 <= ram[addr0_t1];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1_t1) 
            ram[addr1_t1] <= d1_t1; 
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_td_fused_final_fmaps_memcore(
    reset,
    clk,
    address0,
    ce0,
    q0,
    address1,
    ce1,
    we1,
    d1);

parameter DataWidth = 32'd64;
parameter AddressRange = 32'd49000;
parameter AddressWidth = 32'd16;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;



td_fused_top_td_fused_final_fmaps_memcore_ram td_fused_top_td_fused_final_fmaps_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_td_fused_final_fmaps
#(parameter
    DataWidth    = 64,
    AddressRange = 32,
    AddressWidth = 16,
    BufferCount  = 2,
    MemLatency   = 3,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire [AddressWidth-1:0] i_address0,
    output wire [DataWidth-1:0]    i_q0,
    input  wire                    i_ce1,
    input  wire                    i_we1,
    input  wire [AddressWidth-1:0] i_address1,
    input  wire [DataWidth-1:0]    i_d1,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire [AddressWidth-1:0] t_address0,
    output wire [DataWidth-1:0]    t_q0,
    input  wire                    t_ce1,
    input  wire                    t_we1,
    input  wire [AddressWidth-1:0] t_address1,
    input  wire [DataWidth-1:0]    t_d1
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth-1:0]   prev_iptr    = 1'b0; // previous initiator index
reg  [IndexWidth-1:0]   prev_tptr    = 1'b0; // previous target index
reg  [DataWidth-1:0]    reg_q0      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid0    = 1'b0; // buffer has valid data
reg  [DataWidth-1:0]    reg_q1      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid1    = 1'b0; // buffer has valid data
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
// buffer signals
wire [BufferCount-1:0] buf_ce0;
wire [AddressWidth-1:0] buf_a0_0, buf_a0_1;
wire [DataWidth-1:0] buf_q0_0, buf_q0_1;
wire [BufferCount-1:0] buf_ce1;
wire [BufferCount-1:0] buf_we1;
wire [AddressWidth-1:0] buf_a1_0, buf_a1_1;
wire [DataWidth-1:0] buf_d1_0, buf_d1_1;
//------------------------Instantiation------------------
//genvar i;
        td_fused_top_td_fused_final_fmaps_memcore td_fused_top_td_fused_final_fmaps_memcore_U_0 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_0 ),
            .ce0      ( buf_ce0[ 0 ] ),
            .q0       ( buf_q0_0 ),
            .address1 ( buf_a1_0 ),
            .ce1      ( buf_ce1[ 0 ] ),
            .we1      ( buf_we1[ 0 ] ),
            .d1       ( buf_d1_0 )
        );
        td_fused_top_td_fused_final_fmaps_memcore td_fused_top_td_fused_final_fmaps_memcore_U_1 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_1 ),
            .ce0      ( buf_ce0[ 1 ] ),
            .q0       ( buf_q0_1 ),
            .address1 ( buf_a1_1 ),
            .ce1      ( buf_ce1[ 1 ] ),
            .we1      ( buf_we1[ 1 ] ),
            .d1       ( buf_d1_1 )
        );

//++++++++++++++++++++++++buffer signals+++++++++++++++++
        assign buf_ce0[ 0 ] = (tptr ==  0  && empty_n) ? t_ce0
                             : (iptr ==  0 ) ? i_ce0 : 1'b0;
        assign buf_a0_0  = (tptr ==  0  && empty_n) ?  t_address0 : i_address0;
        assign buf_ce1[ 0 ] = (tptr ==  0  && empty_n) ? t_ce1
                             : (iptr ==  0 ) ? i_ce1 : 1'b0;
        assign buf_a1_0  = (tptr ==  0  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 0 ] = (tptr ==  0  && empty_n)  ? t_we1
                             : (iptr ==  0 ) ? i_we1 : 1'b0;
        assign buf_d1_0  = (tptr ==  0  && empty_n) ? t_d1       : i_d1;
        assign buf_ce0[ 1 ] = (tptr ==  1  && empty_n) ? t_ce0
                             : (iptr ==  1 ) ? i_ce0 : 1'b0;
        assign buf_a0_1  = (tptr ==  1  && empty_n) ?  t_address0 : i_address0;
        assign buf_ce1[ 1 ] = (tptr ==  1  && empty_n) ? t_ce1
                             : (iptr ==  1 ) ? i_ce1 : 1'b0;
        assign buf_a1_1  = (tptr ==  1  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 1 ] = (tptr ==  1  && empty_n)  ? t_we1
                             : (iptr ==  1 ) ? i_we1 : 1'b0;
        assign buf_d1_1  = (tptr ==  1  && empty_n) ? t_d1       : i_d1;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//------------------------Body---------------------------
assign i_q0      = (prev_iptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign t_q0      = reg_valid0 ? reg_q0 : (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// prev_iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_iptr <= 1'b0;
    else begin
        prev_iptr <= iptr;
    end
end

// prev_tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_tptr <= 1'b0;
    else begin
        prev_tptr <= tptr;
    end
end

// reg_q0 and reg_valid0
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q0     <= 1'b0;
        reg_valid0 <= 1'b0;
    end else if (!t_ce0 && !reg_valid0) begin
        reg_q0     <= (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
        reg_valid0 <= 1'b1;
    end else if (t_ce0) begin
        reg_valid0 <= 1'b0;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_td_fused_tdf10_fmaps_memcore_ram (addr0, ce0, q0, addr1, ce1, d1, we1,  clk);

parameter DWIDTH = 64;
parameter AWIDTH = 12;
parameter MEM_SIZE = 3136;

input[AWIDTH-1:0] addr0;
input ce0;
output wire[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
input clk;

 reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];
wire [AWIDTH-1:0] addr0_t0; 
reg [AWIDTH-1:0] addr0_t1; 
reg [DWIDTH-1:0] q0_t0;
  reg [DWIDTH-1:0] q0_t1;
wire [AWIDTH-1:0] addr1_t0; 
reg [AWIDTH-1:0] addr1_t1; 
wire [DWIDTH-1:0] d1_t0; 
wire we1_t0; 
reg [DWIDTH-1:0] d1_t1; 
reg we1_t1; 


assign addr0_t0 = addr0;
assign q0 = q0_t1;
assign addr1_t0 = addr1;
assign d1_t0 = d1;
assign we1_t0 = we1;

always @(posedge clk)  
begin
    if (ce0) 
    begin
        addr0_t1 <= addr0_t0; 
        q0_t1 <= q0_t0;
    end
    if (ce1) 
    begin
        addr1_t1 <= addr1_t0; 
        d1_t1 <= d1_t0;
        we1_t1 <= we1_t0;
    end
end


always @(posedge clk)  
begin 
    if (ce0) begin
        q0_t0 <= ram[addr0_t1];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1_t1) 
            ram[addr1_t1] <= d1_t1; 
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_td_fused_tdf10_fmaps_memcore(
    reset,
    clk,
    address0,
    ce0,
    q0,
    address1,
    ce1,
    we1,
    d1);

parameter DataWidth = 32'd64;
parameter AddressRange = 32'd3136;
parameter AddressWidth = 32'd12;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;



td_fused_top_td_fused_tdf10_fmaps_memcore_ram td_fused_top_td_fused_tdf10_fmaps_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_td_fused_tdf10_fmaps
#(parameter
    DataWidth    = 64,
    AddressRange = 32,
    AddressWidth = 12,
    BufferCount  = 2,
    MemLatency   = 3,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire [AddressWidth-1:0] i_address0,
    output wire [DataWidth-1:0]    i_q0,
    input  wire                    i_ce1,
    input  wire                    i_we1,
    input  wire [AddressWidth-1:0] i_address1,
    input  wire [DataWidth-1:0]    i_d1,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire [AddressWidth-1:0] t_address0,
    output wire [DataWidth-1:0]    t_q0,
    input  wire                    t_ce1,
    input  wire                    t_we1,
    input  wire [AddressWidth-1:0] t_address1,
    input  wire [DataWidth-1:0]    t_d1
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth-1:0]   prev_iptr    = 1'b0; // previous initiator index
reg  [IndexWidth-1:0]   prev_tptr    = 1'b0; // previous target index
reg  [DataWidth-1:0]    reg_q0      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid0    = 1'b0; // buffer has valid data
reg  [DataWidth-1:0]    reg_q1      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid1    = 1'b0; // buffer has valid data
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
// buffer signals
wire [BufferCount-1:0] buf_ce0;
wire [AddressWidth-1:0] buf_a0_0, buf_a0_1;
wire [DataWidth-1:0] buf_q0_0, buf_q0_1;
wire [BufferCount-1:0] buf_ce1;
wire [BufferCount-1:0] buf_we1;
wire [AddressWidth-1:0] buf_a1_0, buf_a1_1;
wire [DataWidth-1:0] buf_d1_0, buf_d1_1;
//------------------------Instantiation------------------
//genvar i;
        td_fused_top_td_fused_tdf10_fmaps_memcore td_fused_top_td_fused_tdf10_fmaps_memcore_U_0 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_0 ),
            .ce0      ( buf_ce0[ 0 ] ),
            .q0       ( buf_q0_0 ),
            .address1 ( buf_a1_0 ),
            .ce1      ( buf_ce1[ 0 ] ),
            .we1      ( buf_we1[ 0 ] ),
            .d1       ( buf_d1_0 )
        );
        td_fused_top_td_fused_tdf10_fmaps_memcore td_fused_top_td_fused_tdf10_fmaps_memcore_U_1 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_1 ),
            .ce0      ( buf_ce0[ 1 ] ),
            .q0       ( buf_q0_1 ),
            .address1 ( buf_a1_1 ),
            .ce1      ( buf_ce1[ 1 ] ),
            .we1      ( buf_we1[ 1 ] ),
            .d1       ( buf_d1_1 )
        );

//++++++++++++++++++++++++buffer signals+++++++++++++++++
        assign buf_ce0[ 0 ] = (tptr ==  0  && empty_n) ? t_ce0
                             : (iptr ==  0 ) ? i_ce0 : 1'b0;
        assign buf_a0_0  = (tptr ==  0  && empty_n) ?  t_address0 : i_address0;
        assign buf_ce1[ 0 ] = (tptr ==  0  && empty_n) ? t_ce1
                             : (iptr ==  0 ) ? i_ce1 : 1'b0;
        assign buf_a1_0  = (tptr ==  0  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 0 ] = (tptr ==  0  && empty_n)  ? t_we1
                             : (iptr ==  0 ) ? i_we1 : 1'b0;
        assign buf_d1_0  = (tptr ==  0  && empty_n) ? t_d1       : i_d1;
        assign buf_ce0[ 1 ] = (tptr ==  1  && empty_n) ? t_ce0
                             : (iptr ==  1 ) ? i_ce0 : 1'b0;
        assign buf_a0_1  = (tptr ==  1  && empty_n) ?  t_address0 : i_address0;
        assign buf_ce1[ 1 ] = (tptr ==  1  && empty_n) ? t_ce1
                             : (iptr ==  1 ) ? i_ce1 : 1'b0;
        assign buf_a1_1  = (tptr ==  1  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 1 ] = (tptr ==  1  && empty_n)  ? t_we1
                             : (iptr ==  1 ) ? i_we1 : 1'b0;
        assign buf_d1_1  = (tptr ==  1  && empty_n) ? t_d1       : i_d1;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//------------------------Body---------------------------
assign i_q0      = (prev_iptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign t_q0      = reg_valid0 ? reg_q0 : (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// prev_iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_iptr <= 1'b0;
    else begin
        prev_iptr <= iptr;
    end
end

// prev_tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_tptr <= 1'b0;
    else begin
        prev_tptr <= tptr;
    end
end

// reg_q0 and reg_valid0
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q0     <= 1'b0;
        reg_valid0 <= 1'b0;
    end else if (!t_ce0 && !reg_valid0) begin
        reg_q0     <= (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
        reg_valid0 <= 1'b1;
    end else if (t_ce0) begin
        reg_valid0 <= 1'b0;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_td_fused_tdf1_fmaps_memcore_ram (addr0, ce0, q0, addr1, ce1, d1, we1,  clk);

parameter DWIDTH = 64;
parameter AWIDTH = 16;
parameter MEM_SIZE = 50176;

input[AWIDTH-1:0] addr0;
input ce0;
output wire[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
input clk;

 reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];
wire [AWIDTH-1:0] addr0_t0; 
reg [AWIDTH-1:0] addr0_t1; 
reg [DWIDTH-1:0] q0_t0;
  reg [DWIDTH-1:0] q0_t1;
wire [AWIDTH-1:0] addr1_t0; 
reg [AWIDTH-1:0] addr1_t1; 
wire [DWIDTH-1:0] d1_t0; 
wire we1_t0; 
reg [DWIDTH-1:0] d1_t1; 
reg we1_t1; 


assign addr0_t0 = addr0;
assign q0 = q0_t1;
assign addr1_t0 = addr1;
assign d1_t0 = d1;
assign we1_t0 = we1;

always @(posedge clk)  
begin
    if (ce0) 
    begin
        addr0_t1 <= addr0_t0; 
        q0_t1 <= q0_t0;
    end
    if (ce1) 
    begin
        addr1_t1 <= addr1_t0; 
        d1_t1 <= d1_t0;
        we1_t1 <= we1_t0;
    end
end


always @(posedge clk)  
begin 
    if (ce0) begin
        q0_t0 <= ram[addr0_t1];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1_t1) 
            ram[addr1_t1] <= d1_t1; 
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_td_fused_tdf1_fmaps_memcore(
    reset,
    clk,
    address0,
    ce0,
    q0,
    address1,
    ce1,
    we1,
    d1);

parameter DataWidth = 32'd64;
parameter AddressRange = 32'd50176;
parameter AddressWidth = 32'd16;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;



td_fused_top_td_fused_tdf1_fmaps_memcore_ram td_fused_top_td_fused_tdf1_fmaps_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_td_fused_tdf1_fmaps
#(parameter
    DataWidth    = 64,
    AddressRange = 32,
    AddressWidth = 16,
    BufferCount  = 2,
    MemLatency   = 3,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire [AddressWidth-1:0] i_address0,
    output wire [DataWidth-1:0]    i_q0,
    input  wire                    i_ce1,
    input  wire                    i_we1,
    input  wire [AddressWidth-1:0] i_address1,
    input  wire [DataWidth-1:0]    i_d1,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire [AddressWidth-1:0] t_address0,
    output wire [DataWidth-1:0]    t_q0,
    input  wire                    t_ce1,
    input  wire                    t_we1,
    input  wire [AddressWidth-1:0] t_address1,
    input  wire [DataWidth-1:0]    t_d1
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth-1:0]   prev_iptr    = 1'b0; // previous initiator index
reg  [IndexWidth-1:0]   prev_tptr    = 1'b0; // previous target index
reg  [DataWidth-1:0]    reg_q0      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid0    = 1'b0; // buffer has valid data
reg  [DataWidth-1:0]    reg_q1      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid1    = 1'b0; // buffer has valid data
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
// buffer signals
wire [BufferCount-1:0] buf_ce0;
wire [AddressWidth-1:0] buf_a0_0, buf_a0_1;
wire [DataWidth-1:0] buf_q0_0, buf_q0_1;
wire [BufferCount-1:0] buf_ce1;
wire [BufferCount-1:0] buf_we1;
wire [AddressWidth-1:0] buf_a1_0, buf_a1_1;
wire [DataWidth-1:0] buf_d1_0, buf_d1_1;
//------------------------Instantiation------------------
//genvar i;
        td_fused_top_td_fused_tdf1_fmaps_memcore td_fused_top_td_fused_tdf1_fmaps_memcore_U_0 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_0 ),
            .ce0      ( buf_ce0[ 0 ] ),
            .q0       ( buf_q0_0 ),
            .address1 ( buf_a1_0 ),
            .ce1      ( buf_ce1[ 0 ] ),
            .we1      ( buf_we1[ 0 ] ),
            .d1       ( buf_d1_0 )
        );
        td_fused_top_td_fused_tdf1_fmaps_memcore td_fused_top_td_fused_tdf1_fmaps_memcore_U_1 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_1 ),
            .ce0      ( buf_ce0[ 1 ] ),
            .q0       ( buf_q0_1 ),
            .address1 ( buf_a1_1 ),
            .ce1      ( buf_ce1[ 1 ] ),
            .we1      ( buf_we1[ 1 ] ),
            .d1       ( buf_d1_1 )
        );

//++++++++++++++++++++++++buffer signals+++++++++++++++++
        assign buf_ce0[ 0 ] = (tptr ==  0  && empty_n) ? t_ce0
                             : (iptr ==  0 ) ? i_ce0 : 1'b0;
        assign buf_a0_0  = (tptr ==  0  && empty_n) ?  t_address0 : i_address0;
        assign buf_ce1[ 0 ] = (tptr ==  0  && empty_n) ? t_ce1
                             : (iptr ==  0 ) ? i_ce1 : 1'b0;
        assign buf_a1_0  = (tptr ==  0  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 0 ] = (tptr ==  0  && empty_n)  ? t_we1
                             : (iptr ==  0 ) ? i_we1 : 1'b0;
        assign buf_d1_0  = (tptr ==  0  && empty_n) ? t_d1       : i_d1;
        assign buf_ce0[ 1 ] = (tptr ==  1  && empty_n) ? t_ce0
                             : (iptr ==  1 ) ? i_ce0 : 1'b0;
        assign buf_a0_1  = (tptr ==  1  && empty_n) ?  t_address0 : i_address0;
        assign buf_ce1[ 1 ] = (tptr ==  1  && empty_n) ? t_ce1
                             : (iptr ==  1 ) ? i_ce1 : 1'b0;
        assign buf_a1_1  = (tptr ==  1  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 1 ] = (tptr ==  1  && empty_n)  ? t_we1
                             : (iptr ==  1 ) ? i_we1 : 1'b0;
        assign buf_d1_1  = (tptr ==  1  && empty_n) ? t_d1       : i_d1;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//------------------------Body---------------------------
assign i_q0      = (prev_iptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign t_q0      = reg_valid0 ? reg_q0 : (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// prev_iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_iptr <= 1'b0;
    else begin
        prev_iptr <= iptr;
    end
end

// prev_tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_tptr <= 1'b0;
    else begin
        prev_tptr <= tptr;
    end
end

// reg_q0 and reg_valid0
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q0     <= 1'b0;
        reg_valid0 <= 1'b0;
    end else if (!t_ce0 && !reg_valid0) begin
        reg_q0     <= (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
        reg_valid0 <= 1'b1;
    end else if (t_ce0) begin
        reg_valid0 <= 1'b0;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_td_fused_tdf3_fmaps_memcore_ram (addr0, ce0, q0, addr1, ce1, d1, we1,  clk);

parameter DWIDTH = 64;
parameter AWIDTH = 15;
parameter MEM_SIZE = 25088;

input[AWIDTH-1:0] addr0;
input ce0;
output wire[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
input clk;

 reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];
wire [AWIDTH-1:0] addr0_t0; 
reg [AWIDTH-1:0] addr0_t1; 
reg [DWIDTH-1:0] q0_t0;
  reg [DWIDTH-1:0] q0_t1;
wire [AWIDTH-1:0] addr1_t0; 
reg [AWIDTH-1:0] addr1_t1; 
wire [DWIDTH-1:0] d1_t0; 
wire we1_t0; 
reg [DWIDTH-1:0] d1_t1; 
reg we1_t1; 


assign addr0_t0 = addr0;
assign q0 = q0_t1;
assign addr1_t0 = addr1;
assign d1_t0 = d1;
assign we1_t0 = we1;

always @(posedge clk)  
begin
    if (ce0) 
    begin
        addr0_t1 <= addr0_t0; 
        q0_t1 <= q0_t0;
    end
    if (ce1) 
    begin
        addr1_t1 <= addr1_t0; 
        d1_t1 <= d1_t0;
        we1_t1 <= we1_t0;
    end
end


always @(posedge clk)  
begin 
    if (ce0) begin
        q0_t0 <= ram[addr0_t1];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1_t1) 
            ram[addr1_t1] <= d1_t1; 
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_td_fused_tdf3_fmaps_memcore(
    reset,
    clk,
    address0,
    ce0,
    q0,
    address1,
    ce1,
    we1,
    d1);

parameter DataWidth = 32'd64;
parameter AddressRange = 32'd25088;
parameter AddressWidth = 32'd15;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;



td_fused_top_td_fused_tdf3_fmaps_memcore_ram td_fused_top_td_fused_tdf3_fmaps_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_td_fused_tdf3_fmaps
#(parameter
    DataWidth    = 64,
    AddressRange = 32,
    AddressWidth = 15,
    BufferCount  = 2,
    MemLatency   = 3,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire [AddressWidth-1:0] i_address0,
    output wire [DataWidth-1:0]    i_q0,
    input  wire                    i_ce1,
    input  wire                    i_we1,
    input  wire [AddressWidth-1:0] i_address1,
    input  wire [DataWidth-1:0]    i_d1,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire [AddressWidth-1:0] t_address0,
    output wire [DataWidth-1:0]    t_q0,
    input  wire                    t_ce1,
    input  wire                    t_we1,
    input  wire [AddressWidth-1:0] t_address1,
    input  wire [DataWidth-1:0]    t_d1
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth-1:0]   prev_iptr    = 1'b0; // previous initiator index
reg  [IndexWidth-1:0]   prev_tptr    = 1'b0; // previous target index
reg  [DataWidth-1:0]    reg_q0      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid0    = 1'b0; // buffer has valid data
reg  [DataWidth-1:0]    reg_q1      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid1    = 1'b0; // buffer has valid data
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
// buffer signals
wire [BufferCount-1:0] buf_ce0;
wire [AddressWidth-1:0] buf_a0_0, buf_a0_1;
wire [DataWidth-1:0] buf_q0_0, buf_q0_1;
wire [BufferCount-1:0] buf_ce1;
wire [BufferCount-1:0] buf_we1;
wire [AddressWidth-1:0] buf_a1_0, buf_a1_1;
wire [DataWidth-1:0] buf_d1_0, buf_d1_1;
//------------------------Instantiation------------------
//genvar i;
        td_fused_top_td_fused_tdf3_fmaps_memcore td_fused_top_td_fused_tdf3_fmaps_memcore_U_0 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_0 ),
            .ce0      ( buf_ce0[ 0 ] ),
            .q0       ( buf_q0_0 ),
            .address1 ( buf_a1_0 ),
            .ce1      ( buf_ce1[ 0 ] ),
            .we1      ( buf_we1[ 0 ] ),
            .d1       ( buf_d1_0 )
        );
        td_fused_top_td_fused_tdf3_fmaps_memcore td_fused_top_td_fused_tdf3_fmaps_memcore_U_1 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_1 ),
            .ce0      ( buf_ce0[ 1 ] ),
            .q0       ( buf_q0_1 ),
            .address1 ( buf_a1_1 ),
            .ce1      ( buf_ce1[ 1 ] ),
            .we1      ( buf_we1[ 1 ] ),
            .d1       ( buf_d1_1 )
        );

//++++++++++++++++++++++++buffer signals+++++++++++++++++
        assign buf_ce0[ 0 ] = (tptr ==  0  && empty_n) ? t_ce0
                             : (iptr ==  0 ) ? i_ce0 : 1'b0;
        assign buf_a0_0  = (tptr ==  0  && empty_n) ?  t_address0 : i_address0;
        assign buf_ce1[ 0 ] = (tptr ==  0  && empty_n) ? t_ce1
                             : (iptr ==  0 ) ? i_ce1 : 1'b0;
        assign buf_a1_0  = (tptr ==  0  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 0 ] = (tptr ==  0  && empty_n)  ? t_we1
                             : (iptr ==  0 ) ? i_we1 : 1'b0;
        assign buf_d1_0  = (tptr ==  0  && empty_n) ? t_d1       : i_d1;
        assign buf_ce0[ 1 ] = (tptr ==  1  && empty_n) ? t_ce0
                             : (iptr ==  1 ) ? i_ce0 : 1'b0;
        assign buf_a0_1  = (tptr ==  1  && empty_n) ?  t_address0 : i_address0;
        assign buf_ce1[ 1 ] = (tptr ==  1  && empty_n) ? t_ce1
                             : (iptr ==  1 ) ? i_ce1 : 1'b0;
        assign buf_a1_1  = (tptr ==  1  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 1 ] = (tptr ==  1  && empty_n)  ? t_we1
                             : (iptr ==  1 ) ? i_we1 : 1'b0;
        assign buf_d1_1  = (tptr ==  1  && empty_n) ? t_d1       : i_d1;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//------------------------Body---------------------------
assign i_q0      = (prev_iptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign t_q0      = reg_valid0 ? reg_q0 : (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// prev_iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_iptr <= 1'b0;
    else begin
        prev_iptr <= iptr;
    end
end

// prev_tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_tptr <= 1'b0;
    else begin
        prev_tptr <= tptr;
    end
end

// reg_q0 and reg_valid0
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q0     <= 1'b0;
        reg_valid0 <= 1'b0;
    end else if (!t_ce0 && !reg_valid0) begin
        reg_q0     <= (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
        reg_valid0 <= 1'b1;
    end else if (t_ce0) begin
        reg_valid0 <= 1'b0;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_td_fused_tdf4_fmaps_memcore_ram (addr0, ce0, q0, addr1, ce1, d1, we1,  clk);

parameter DWIDTH = 64;
parameter AWIDTH = 14;
parameter MEM_SIZE = 12544;

input[AWIDTH-1:0] addr0;
input ce0;
output wire[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
input clk;

 reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];
wire [AWIDTH-1:0] addr0_t0; 
reg [AWIDTH-1:0] addr0_t1; 
reg [DWIDTH-1:0] q0_t0;
  reg [DWIDTH-1:0] q0_t1;
wire [AWIDTH-1:0] addr1_t0; 
reg [AWIDTH-1:0] addr1_t1; 
wire [DWIDTH-1:0] d1_t0; 
wire we1_t0; 
reg [DWIDTH-1:0] d1_t1; 
reg we1_t1; 


assign addr0_t0 = addr0;
assign q0 = q0_t1;
assign addr1_t0 = addr1;
assign d1_t0 = d1;
assign we1_t0 = we1;

always @(posedge clk)  
begin
    if (ce0) 
    begin
        addr0_t1 <= addr0_t0; 
        q0_t1 <= q0_t0;
    end
    if (ce1) 
    begin
        addr1_t1 <= addr1_t0; 
        d1_t1 <= d1_t0;
        we1_t1 <= we1_t0;
    end
end


always @(posedge clk)  
begin 
    if (ce0) begin
        q0_t0 <= ram[addr0_t1];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1_t1) 
            ram[addr1_t1] <= d1_t1; 
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_td_fused_tdf4_fmaps_memcore(
    reset,
    clk,
    address0,
    ce0,
    q0,
    address1,
    ce1,
    we1,
    d1);

parameter DataWidth = 32'd64;
parameter AddressRange = 32'd12544;
parameter AddressWidth = 32'd14;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;



td_fused_top_td_fused_tdf4_fmaps_memcore_ram td_fused_top_td_fused_tdf4_fmaps_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_td_fused_tdf4_fmaps
#(parameter
    DataWidth    = 64,
    AddressRange = 32,
    AddressWidth = 14,
    BufferCount  = 2,
    MemLatency   = 3,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire [AddressWidth-1:0] i_address0,
    output wire [DataWidth-1:0]    i_q0,
    input  wire                    i_ce1,
    input  wire                    i_we1,
    input  wire [AddressWidth-1:0] i_address1,
    input  wire [DataWidth-1:0]    i_d1,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire [AddressWidth-1:0] t_address0,
    output wire [DataWidth-1:0]    t_q0,
    input  wire                    t_ce1,
    input  wire                    t_we1,
    input  wire [AddressWidth-1:0] t_address1,
    input  wire [DataWidth-1:0]    t_d1
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth-1:0]   prev_iptr    = 1'b0; // previous initiator index
reg  [IndexWidth-1:0]   prev_tptr    = 1'b0; // previous target index
reg  [DataWidth-1:0]    reg_q0      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid0    = 1'b0; // buffer has valid data
reg  [DataWidth-1:0]    reg_q1      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid1    = 1'b0; // buffer has valid data
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
// buffer signals
wire [BufferCount-1:0] buf_ce0;
wire [AddressWidth-1:0] buf_a0_0, buf_a0_1;
wire [DataWidth-1:0] buf_q0_0, buf_q0_1;
wire [BufferCount-1:0] buf_ce1;
wire [BufferCount-1:0] buf_we1;
wire [AddressWidth-1:0] buf_a1_0, buf_a1_1;
wire [DataWidth-1:0] buf_d1_0, buf_d1_1;
//------------------------Instantiation------------------
//genvar i;
        td_fused_top_td_fused_tdf4_fmaps_memcore td_fused_top_td_fused_tdf4_fmaps_memcore_U_0 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_0 ),
            .ce0      ( buf_ce0[ 0 ] ),
            .q0       ( buf_q0_0 ),
            .address1 ( buf_a1_0 ),
            .ce1      ( buf_ce1[ 0 ] ),
            .we1      ( buf_we1[ 0 ] ),
            .d1       ( buf_d1_0 )
        );
        td_fused_top_td_fused_tdf4_fmaps_memcore td_fused_top_td_fused_tdf4_fmaps_memcore_U_1 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_1 ),
            .ce0      ( buf_ce0[ 1 ] ),
            .q0       ( buf_q0_1 ),
            .address1 ( buf_a1_1 ),
            .ce1      ( buf_ce1[ 1 ] ),
            .we1      ( buf_we1[ 1 ] ),
            .d1       ( buf_d1_1 )
        );

//++++++++++++++++++++++++buffer signals+++++++++++++++++
        assign buf_ce0[ 0 ] = (tptr ==  0  && empty_n) ? t_ce0
                             : (iptr ==  0 ) ? i_ce0 : 1'b0;
        assign buf_a0_0  = (tptr ==  0  && empty_n) ?  t_address0 : i_address0;
        assign buf_ce1[ 0 ] = (tptr ==  0  && empty_n) ? t_ce1
                             : (iptr ==  0 ) ? i_ce1 : 1'b0;
        assign buf_a1_0  = (tptr ==  0  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 0 ] = (tptr ==  0  && empty_n)  ? t_we1
                             : (iptr ==  0 ) ? i_we1 : 1'b0;
        assign buf_d1_0  = (tptr ==  0  && empty_n) ? t_d1       : i_d1;
        assign buf_ce0[ 1 ] = (tptr ==  1  && empty_n) ? t_ce0
                             : (iptr ==  1 ) ? i_ce0 : 1'b0;
        assign buf_a0_1  = (tptr ==  1  && empty_n) ?  t_address0 : i_address0;
        assign buf_ce1[ 1 ] = (tptr ==  1  && empty_n) ? t_ce1
                             : (iptr ==  1 ) ? i_ce1 : 1'b0;
        assign buf_a1_1  = (tptr ==  1  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 1 ] = (tptr ==  1  && empty_n)  ? t_we1
                             : (iptr ==  1 ) ? i_we1 : 1'b0;
        assign buf_d1_1  = (tptr ==  1  && empty_n) ? t_d1       : i_d1;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//------------------------Body---------------------------
assign i_q0      = (prev_iptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign t_q0      = reg_valid0 ? reg_q0 : (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// prev_iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_iptr <= 1'b0;
    else begin
        prev_iptr <= iptr;
    end
end

// prev_tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_tptr <= 1'b0;
    else begin
        prev_tptr <= tptr;
    end
end

// reg_q0 and reg_valid0
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q0     <= 1'b0;
        reg_valid0 <= 1'b0;
    end else if (!t_ce0 && !reg_valid0) begin
        reg_q0     <= (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
        reg_valid0 <= 1'b1;
    end else if (t_ce0) begin
        reg_valid0 <= 1'b0;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module td_fused_top_td_fused_tdf7_fmaps_memcore_ram (addr0, ce0, q0, addr1, ce1, d1, we1,  clk);

parameter DWIDTH = 64;
parameter AWIDTH = 13;
parameter MEM_SIZE = 6272;

input[AWIDTH-1:0] addr0;
input ce0;
output wire[DWIDTH-1:0] q0;
input[AWIDTH-1:0] addr1;
input ce1;
input[DWIDTH-1:0] d1;
input we1;
input clk;

 reg [DWIDTH-1:0] ram[MEM_SIZE-1:0];
wire [AWIDTH-1:0] addr0_t0; 
reg [AWIDTH-1:0] addr0_t1; 
reg [DWIDTH-1:0] q0_t0;
  reg [DWIDTH-1:0] q0_t1;
wire [AWIDTH-1:0] addr1_t0; 
reg [AWIDTH-1:0] addr1_t1; 
wire [DWIDTH-1:0] d1_t0; 
wire we1_t0; 
reg [DWIDTH-1:0] d1_t1; 
reg we1_t1; 


assign addr0_t0 = addr0;
assign q0 = q0_t1;
assign addr1_t0 = addr1;
assign d1_t0 = d1;
assign we1_t0 = we1;

always @(posedge clk)  
begin
    if (ce0) 
    begin
        addr0_t1 <= addr0_t0; 
        q0_t1 <= q0_t0;
    end
    if (ce1) 
    begin
        addr1_t1 <= addr1_t0; 
        d1_t1 <= d1_t0;
        we1_t1 <= we1_t0;
    end
end


always @(posedge clk)  
begin 
    if (ce0) begin
        q0_t0 <= ram[addr0_t1];
    end
end


always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1_t1) 
            ram[addr1_t1] <= d1_t1; 
    end
end


endmodule

`timescale 1 ns / 1 ps
module td_fused_top_td_fused_tdf7_fmaps_memcore(
    reset,
    clk,
    address0,
    ce0,
    q0,
    address1,
    ce1,
    we1,
    d1);

parameter DataWidth = 32'd64;
parameter AddressRange = 32'd6272;
parameter AddressWidth = 32'd13;
input reset;
input clk;
input[AddressWidth - 1:0] address0;
input ce0;
output[DataWidth - 1:0] q0;
input[AddressWidth - 1:0] address1;
input ce1;
input we1;
input[DataWidth - 1:0] d1;



td_fused_top_td_fused_tdf7_fmaps_memcore_ram td_fused_top_td_fused_tdf7_fmaps_memcore_ram_U(
    .clk( clk ),
    .addr0( address0 ),
    .ce0( ce0 ),
    .q0( q0 ),
    .addr1( address1 ),
    .ce1( ce1 ),
    .we1( we1 ),
    .d1( d1 )
);

endmodule

// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1ns/1ps

module td_fused_top_td_fused_tdf7_fmaps
#(parameter
    DataWidth    = 64,
    AddressRange = 32,
    AddressWidth = 13,
    BufferCount  = 2,
    MemLatency   = 3,
    IndexWidth   = 1
) (
    // system signals
    input  wire                    clk,
    input  wire                    reset,
    // initiator
    input  wire                    i_ce,
    input  wire                    i_write,
    output wire                    i_full_n,
    input  wire                    i_ce0,
    input  wire [AddressWidth-1:0] i_address0,
    output wire [DataWidth-1:0]    i_q0,
    input  wire                    i_ce1,
    input  wire                    i_we1,
    input  wire [AddressWidth-1:0] i_address1,
    input  wire [DataWidth-1:0]    i_d1,
    // target
    input  wire                    t_ce,
    input  wire                    t_read,
    output wire                    t_empty_n,
    input  wire                    t_ce0,
    input  wire [AddressWidth-1:0] t_address0,
    output wire [DataWidth-1:0]    t_q0,
    input  wire                    t_ce1,
    input  wire                    t_we1,
    input  wire [AddressWidth-1:0] t_address1,
    input  wire [DataWidth-1:0]    t_d1
);
//------------------------Local signal-------------------
// control/status
reg  [IndexWidth-1:0]   iptr    = 1'b0; // initiator index
reg  [IndexWidth-1:0]   tptr    = 1'b0; // target index
reg  [IndexWidth-1:0]   prev_iptr    = 1'b0; // previous initiator index
reg  [IndexWidth-1:0]   prev_tptr    = 1'b0; // previous target index
reg  [DataWidth-1:0]    reg_q0      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid0    = 1'b0; // buffer has valid data
reg  [DataWidth-1:0]    reg_q1      = 1'b0; // buffer used if reader is stalled
reg                     reg_valid1    = 1'b0; // buffer has valid data
reg  [IndexWidth:0]     count   = 1'b0; // count of written buffers
reg                     full_n  = 1'b1; // whether all buffers are written
reg                     empty_n = 1'b0; // whether none of the buffers is written
wire                    push_buf;       // finish writing a buffer
wire                    write_buf;      // write a buffer
wire                    pop_buf;        // finish reading a buffer
// buffer signals
wire [BufferCount-1:0] buf_ce0;
wire [AddressWidth-1:0] buf_a0_0, buf_a0_1;
wire [DataWidth-1:0] buf_q0_0, buf_q0_1;
wire [BufferCount-1:0] buf_ce1;
wire [BufferCount-1:0] buf_we1;
wire [AddressWidth-1:0] buf_a1_0, buf_a1_1;
wire [DataWidth-1:0] buf_d1_0, buf_d1_1;
//------------------------Instantiation------------------
//genvar i;
        td_fused_top_td_fused_tdf7_fmaps_memcore td_fused_top_td_fused_tdf7_fmaps_memcore_U_0 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_0 ),
            .ce0      ( buf_ce0[ 0 ] ),
            .q0       ( buf_q0_0 ),
            .address1 ( buf_a1_0 ),
            .ce1      ( buf_ce1[ 0 ] ),
            .we1      ( buf_we1[ 0 ] ),
            .d1       ( buf_d1_0 )
        );
        td_fused_top_td_fused_tdf7_fmaps_memcore td_fused_top_td_fused_tdf7_fmaps_memcore_U_1 (
            .reset    ( reset ),
            .clk      ( clk ),
            .address0 ( buf_a0_1 ),
            .ce0      ( buf_ce0[ 1 ] ),
            .q0       ( buf_q0_1 ),
            .address1 ( buf_a1_1 ),
            .ce1      ( buf_ce1[ 1 ] ),
            .we1      ( buf_we1[ 1 ] ),
            .d1       ( buf_d1_1 )
        );

//++++++++++++++++++++++++buffer signals+++++++++++++++++
        assign buf_ce0[ 0 ] = (tptr ==  0  && empty_n) ? t_ce0
                             : (iptr ==  0 ) ? i_ce0 : 1'b0;
        assign buf_a0_0  = (tptr ==  0  && empty_n) ?  t_address0 : i_address0;
        assign buf_ce1[ 0 ] = (tptr ==  0  && empty_n) ? t_ce1
                             : (iptr ==  0 ) ? i_ce1 : 1'b0;
        assign buf_a1_0  = (tptr ==  0  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 0 ] = (tptr ==  0  && empty_n)  ? t_we1
                             : (iptr ==  0 ) ? i_we1 : 1'b0;
        assign buf_d1_0  = (tptr ==  0  && empty_n) ? t_d1       : i_d1;
        assign buf_ce0[ 1 ] = (tptr ==  1  && empty_n) ? t_ce0
                             : (iptr ==  1 ) ? i_ce0 : 1'b0;
        assign buf_a0_1  = (tptr ==  1  && empty_n) ?  t_address0 : i_address0;
        assign buf_ce1[ 1 ] = (tptr ==  1  && empty_n) ? t_ce1
                             : (iptr ==  1 ) ? i_ce1 : 1'b0;
        assign buf_a1_1  = (tptr ==  1  && empty_n) ?  t_address1 : i_address1;
        assign buf_we1[ 1 ] = (tptr ==  1  && empty_n)  ? t_we1
                             : (iptr ==  1 ) ? i_we1 : 1'b0;
        assign buf_d1_1  = (tptr ==  1  && empty_n) ? t_d1       : i_d1;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//------------------------Body---------------------------
assign i_q0      = (prev_iptr == 1'b1 ? buf_q0_1 : buf_q0_0);
assign t_q0      = reg_valid0 ? reg_q0 : (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);

//++++++++++++++++++++++++output+++++++++++++++++++++++++
assign i_full_n  = full_n;
assign t_empty_n = empty_n;
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

//++++++++++++++++++++++++control/status+++++++++++++++++
assign push_buf = i_ce & i_write & full_n;
assign write_buf = i_ce & i_write;
assign pop_buf  = t_ce & t_read & empty_n;

// iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        iptr <= 1'b0;
    else if (push_buf) begin
        if (iptr == BufferCount - 1'b1)
            iptr <= 1'b0;
        else
            iptr <= iptr + 1'b1;
    end
end

// tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        tptr <= 1'b0;
    else if (pop_buf) begin
        if (tptr == BufferCount - 1'b1)
            tptr <= 1'b0;
        else
            tptr <= tptr + 1'b1;
    end
end

// prev_iptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_iptr <= 1'b0;
    else begin
        prev_iptr <= iptr;
    end
end

// prev_tptr
always @(posedge clk) begin
    if (reset == 1'b1)
        prev_tptr <= 1'b0;
    else begin
        prev_tptr <= tptr;
    end
end

// reg_q0 and reg_valid0
always @(posedge clk) begin
    if (reset == 1'b1) begin
        reg_q0     <= 1'b0;
        reg_valid0 <= 1'b0;
    end else if (!t_ce0 && !reg_valid0) begin
        reg_q0     <= (prev_tptr == 1'b1 ? buf_q0_1 : buf_q0_0);
        reg_valid0 <= 1'b1;
    end else if (t_ce0) begin
        reg_valid0 <= 1'b0;
    end
end

// count
always @(posedge clk) begin
    if (reset == 1'b1)
        count <= 1'b0;
    else if (push_buf && !pop_buf)
        count <= count + 1'b1;
    else if (!push_buf && pop_buf)
        count <= count - 1'b1;
end

// full_n
always @(posedge clk) begin
    if (reset == 1'b1)
        full_n <= 1'b1;
    else if (push_buf && !pop_buf && count == BufferCount - 2'd2)
        full_n <= 1'b0;
    else if (!push_buf && pop_buf)
        full_n <= 1'b1;
end

// empty_n
always @(posedge clk) begin
    if (reset == 1'b1)
        empty_n <= 1'b0;
    else if ((!write_buf && pop_buf && count == 1'b1)
             || (pop_buf && count == 1'b0))
        empty_n <= 1'b0;
    else if (write_buf && !pop_buf)
        empty_n <= 1'b1;
end
//+++++++++++++++++++++++++++++++++++++++++++++++++++++++

endmodule

// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module td_fused_top_td_fused (
        ap_clk,
        ap_rst,
        tdf1_filters_address0,
        tdf1_filters_ce0,
        tdf1_filters_d0,
        tdf1_filters_q0,
        tdf1_filters_we0,
        tdf1_filters_address1,
        tdf1_filters_ce1,
        tdf1_filters_d1,
        tdf1_filters_q1,
        tdf1_filters_we1,
        tdf2_filters_address0,
        tdf2_filters_ce0,
        tdf2_filters_d0,
        tdf2_filters_q0,
        tdf2_filters_we0,
        tdf2_filters_address1,
        tdf2_filters_ce1,
        tdf2_filters_d1,
        tdf2_filters_q1,
        tdf2_filters_we1,
        tdf3_filters_address0,
        tdf3_filters_ce0,
        tdf3_filters_d0,
        tdf3_filters_q0,
        tdf3_filters_we0,
        tdf3_filters_address1,
        tdf3_filters_ce1,
        tdf3_filters_d1,
        tdf3_filters_q1,
        tdf3_filters_we1,
        tdf4_filters_address0,
        tdf4_filters_ce0,
        tdf4_filters_d0,
        tdf4_filters_q0,
        tdf4_filters_we0,
        tdf4_filters_address1,
        tdf4_filters_ce1,
        tdf4_filters_d1,
        tdf4_filters_q1,
        tdf4_filters_we1,
        tdf4_l2_filters_address0,
        tdf4_l2_filters_ce0,
        tdf4_l2_filters_d0,
        tdf4_l2_filters_q0,
        tdf4_l2_filters_we0,
        tdf4_l2_filters_address1,
        tdf4_l2_filters_ce1,
        tdf4_l2_filters_d1,
        tdf4_l2_filters_q1,
        tdf4_l2_filters_we1,
        tdf5_filters_address0,
        tdf5_filters_ce0,
        tdf5_filters_d0,
        tdf5_filters_q0,
        tdf5_filters_we0,
        tdf5_filters_address1,
        tdf5_filters_ce1,
        tdf5_filters_d1,
        tdf5_filters_q1,
        tdf5_filters_we1,
        tdf6_filters_address0,
        tdf6_filters_ce0,
        tdf6_filters_d0,
        tdf6_filters_q0,
        tdf6_filters_we0,
        tdf6_filters_address1,
        tdf6_filters_ce1,
        tdf6_filters_d1,
        tdf6_filters_q1,
        tdf6_filters_we1,
        tdf7_filters_address0,
        tdf7_filters_ce0,
        tdf7_filters_d0,
        tdf7_filters_q0,
        tdf7_filters_we0,
        tdf7_filters_address1,
        tdf7_filters_ce1,
        tdf7_filters_d1,
        tdf7_filters_q1,
        tdf7_filters_we1,
        tdf7_l2_filters_address0,
        tdf7_l2_filters_ce0,
        tdf7_l2_filters_d0,
        tdf7_l2_filters_q0,
        tdf7_l2_filters_we0,
        tdf7_l2_filters_address1,
        tdf7_l2_filters_ce1,
        tdf7_l2_filters_d1,
        tdf7_l2_filters_q1,
        tdf7_l2_filters_we1,
        tdf8_filters_address0,
        tdf8_filters_ce0,
        tdf8_filters_d0,
        tdf8_filters_q0,
        tdf8_filters_we0,
        tdf8_filters_address1,
        tdf8_filters_ce1,
        tdf8_filters_d1,
        tdf8_filters_q1,
        tdf8_filters_we1,
        tdf9_filters_address0,
        tdf9_filters_ce0,
        tdf9_filters_d0,
        tdf9_filters_q0,
        tdf9_filters_we0,
        tdf9_filters_address1,
        tdf9_filters_ce1,
        tdf9_filters_d1,
        tdf9_filters_q1,
        tdf9_filters_we1,
        tdf10_filters_address0,
        tdf10_filters_ce0,
        tdf10_filters_d0,
        tdf10_filters_q0,
        tdf10_filters_we0,
        tdf10_filters_address1,
        tdf10_filters_ce1,
        tdf10_filters_d1,
        tdf10_filters_q1,
        tdf10_filters_we1,
        tdf10_l2_filters_address0,
        tdf10_l2_filters_ce0,
        tdf10_l2_filters_d0,
        tdf10_l2_filters_q0,
        tdf10_l2_filters_we0,
        tdf10_l2_filters_address1,
        tdf10_l2_filters_ce1,
        tdf10_l2_filters_d1,
        tdf10_l2_filters_q1,
        tdf10_l2_filters_we1,
        tdf11_filters_address0,
        tdf11_filters_ce0,
        tdf11_filters_d0,
        tdf11_filters_q0,
        tdf11_filters_we0,
        tdf11_filters_address1,
        tdf11_filters_ce1,
        tdf11_filters_d1,
        tdf11_filters_q1,
        tdf11_filters_we1,
        tdf11_l2_filters_address0,
        tdf11_l2_filters_ce0,
        tdf11_l2_filters_d0,
        tdf11_l2_filters_q0,
        tdf11_l2_filters_we0,
        tdf11_l2_filters_address1,
        tdf11_l2_filters_ce1,
        tdf11_l2_filters_d1,
        tdf11_l2_filters_q1,
        tdf11_l2_filters_we1,
        tdf12_filters_address0,
        tdf12_filters_ce0,
        tdf12_filters_d0,
        tdf12_filters_q0,
        tdf12_filters_we0,
        tdf12_filters_address1,
        tdf12_filters_ce1,
        tdf12_filters_d1,
        tdf12_filters_q1,
        tdf12_filters_we1,
        tdf1_adjustments_address0,
        tdf1_adjustments_ce0,
        tdf1_adjustments_d0,
        tdf1_adjustments_q0,
        tdf1_adjustments_we0,
        tdf1_adjustments_address1,
        tdf1_adjustments_ce1,
        tdf1_adjustments_d1,
        tdf1_adjustments_q1,
        tdf1_adjustments_we1,
        tdf2_adjustments_address0,
        tdf2_adjustments_ce0,
        tdf2_adjustments_d0,
        tdf2_adjustments_q0,
        tdf2_adjustments_we0,
        tdf2_adjustments_address1,
        tdf2_adjustments_ce1,
        tdf2_adjustments_d1,
        tdf2_adjustments_q1,
        tdf2_adjustments_we1,
        tdf3_adjustments_address0,
        tdf3_adjustments_ce0,
        tdf3_adjustments_d0,
        tdf3_adjustments_q0,
        tdf3_adjustments_we0,
        tdf3_adjustments_address1,
        tdf3_adjustments_ce1,
        tdf3_adjustments_d1,
        tdf3_adjustments_q1,
        tdf3_adjustments_we1,
        tdf4_adjustments_address0,
        tdf4_adjustments_ce0,
        tdf4_adjustments_d0,
        tdf4_adjustments_q0,
        tdf4_adjustments_we0,
        tdf4_adjustments_address1,
        tdf4_adjustments_ce1,
        tdf4_adjustments_d1,
        tdf4_adjustments_q1,
        tdf4_adjustments_we1,
        tdf4_l2_adjustments_address0,
        tdf4_l2_adjustments_ce0,
        tdf4_l2_adjustments_d0,
        tdf4_l2_adjustments_q0,
        tdf4_l2_adjustments_we0,
        tdf4_l2_adjustments_address1,
        tdf4_l2_adjustments_ce1,
        tdf4_l2_adjustments_d1,
        tdf4_l2_adjustments_q1,
        tdf4_l2_adjustments_we1,
        tdf5_adjustments_address0,
        tdf5_adjustments_ce0,
        tdf5_adjustments_d0,
        tdf5_adjustments_q0,
        tdf5_adjustments_we0,
        tdf5_adjustments_address1,
        tdf5_adjustments_ce1,
        tdf5_adjustments_d1,
        tdf5_adjustments_q1,
        tdf5_adjustments_we1,
        tdf6_adjustments_address0,
        tdf6_adjustments_ce0,
        tdf6_adjustments_d0,
        tdf6_adjustments_q0,
        tdf6_adjustments_we0,
        tdf6_adjustments_address1,
        tdf6_adjustments_ce1,
        tdf6_adjustments_d1,
        tdf6_adjustments_q1,
        tdf6_adjustments_we1,
        tdf7_adjustments_address0,
        tdf7_adjustments_ce0,
        tdf7_adjustments_d0,
        tdf7_adjustments_q0,
        tdf7_adjustments_we0,
        tdf7_adjustments_address1,
        tdf7_adjustments_ce1,
        tdf7_adjustments_d1,
        tdf7_adjustments_q1,
        tdf7_adjustments_we1,
        tdf7_l2_adjustments_address0,
        tdf7_l2_adjustments_ce0,
        tdf7_l2_adjustments_d0,
        tdf7_l2_adjustments_q0,
        tdf7_l2_adjustments_we0,
        tdf7_l2_adjustments_address1,
        tdf7_l2_adjustments_ce1,
        tdf7_l2_adjustments_d1,
        tdf7_l2_adjustments_q1,
        tdf7_l2_adjustments_we1,
        tdf8_adjustments_address0,
        tdf8_adjustments_ce0,
        tdf8_adjustments_d0,
        tdf8_adjustments_q0,
        tdf8_adjustments_we0,
        tdf8_adjustments_address1,
        tdf8_adjustments_ce1,
        tdf8_adjustments_d1,
        tdf8_adjustments_q1,
        tdf8_adjustments_we1,
        tdf9_adjustments_address0,
        tdf9_adjustments_ce0,
        tdf9_adjustments_d0,
        tdf9_adjustments_q0,
        tdf9_adjustments_we0,
        tdf9_adjustments_address1,
        tdf9_adjustments_ce1,
        tdf9_adjustments_d1,
        tdf9_adjustments_q1,
        tdf9_adjustments_we1,
        tdf10_adjustments_address0,
        tdf10_adjustments_ce0,
        tdf10_adjustments_d0,
        tdf10_adjustments_q0,
        tdf10_adjustments_we0,
        tdf10_adjustments_address1,
        tdf10_adjustments_ce1,
        tdf10_adjustments_d1,
        tdf10_adjustments_q1,
        tdf10_adjustments_we1,
        tdf10_l2_adjustments_address0,
        tdf10_l2_adjustments_ce0,
        tdf10_l2_adjustments_d0,
        tdf10_l2_adjustments_q0,
        tdf10_l2_adjustments_we0,
        tdf10_l2_adjustments_address1,
        tdf10_l2_adjustments_ce1,
        tdf10_l2_adjustments_d1,
        tdf10_l2_adjustments_q1,
        tdf10_l2_adjustments_we1,
        tdf11_adjustments_address0,
        tdf11_adjustments_ce0,
        tdf11_adjustments_d0,
        tdf11_adjustments_q0,
        tdf11_adjustments_we0,
        tdf11_adjustments_address1,
        tdf11_adjustments_ce1,
        tdf11_adjustments_d1,
        tdf11_adjustments_q1,
        tdf11_adjustments_we1,
        tdf11_l2_adjustments_address0,
        tdf11_l2_adjustments_ce0,
        tdf11_l2_adjustments_d0,
        tdf11_l2_adjustments_q0,
        tdf11_l2_adjustments_we0,
        tdf11_l2_adjustments_address1,
        tdf11_l2_adjustments_ce1,
        tdf11_l2_adjustments_d1,
        tdf11_l2_adjustments_q1,
        tdf11_l2_adjustments_we1,
        tdf12_adjustments_address0,
        tdf12_adjustments_ce0,
        tdf12_adjustments_d0,
        tdf12_adjustments_q0,
        tdf12_adjustments_we0,
        tdf12_adjustments_address1,
        tdf12_adjustments_ce1,
        tdf12_adjustments_d1,
        tdf12_adjustments_q1,
        tdf12_adjustments_we1,
        stream_in_TDATA,
        stream_in_TKEEP,
        stream_in_TSTRB,
        stream_in_TLAST,
        stream_out_TDATA,
        stream_out_TKEEP,
        stream_out_TSTRB,
        stream_out_TLAST,
        stream_in_TVALID,
        stream_in_TREADY,
        ap_start,
        stream_out_TVALID,
        stream_out_TREADY,
        ap_done,
        ap_ready,
        ap_idle,
        ap_continue
);


input   ap_clk;
input   ap_rst;
output  [8:0] tdf1_filters_address0;
output   tdf1_filters_ce0;
output  [15:0] tdf1_filters_d0;
input  [15:0] tdf1_filters_q0;
output   tdf1_filters_we0;
output  [8:0] tdf1_filters_address1;
output   tdf1_filters_ce1;
output  [15:0] tdf1_filters_d1;
input  [15:0] tdf1_filters_q1;
output   tdf1_filters_we1;
output  [12:0] tdf2_filters_address0;
output   tdf2_filters_ce0;
output  [15:0] tdf2_filters_d0;
input  [15:0] tdf2_filters_q0;
output   tdf2_filters_we0;
output  [12:0] tdf2_filters_address1;
output   tdf2_filters_ce1;
output  [15:0] tdf2_filters_d1;
input  [15:0] tdf2_filters_q1;
output   tdf2_filters_we1;
output  [8:0] tdf3_filters_address0;
output   tdf3_filters_ce0;
output  [15:0] tdf3_filters_d0;
input  [15:0] tdf3_filters_q0;
output   tdf3_filters_we0;
output  [8:0] tdf3_filters_address1;
output   tdf3_filters_ce1;
output  [15:0] tdf3_filters_d1;
input  [15:0] tdf3_filters_q1;
output   tdf3_filters_we1;
output  [14:0] tdf4_filters_address0;
output   tdf4_filters_ce0;
output  [15:0] tdf4_filters_d0;
input  [15:0] tdf4_filters_q0;
output   tdf4_filters_we0;
output  [14:0] tdf4_filters_address1;
output   tdf4_filters_ce1;
output  [15:0] tdf4_filters_d1;
input  [15:0] tdf4_filters_q1;
output   tdf4_filters_we1;
output  [10:0] tdf4_l2_filters_address0;
output   tdf4_l2_filters_ce0;
output  [15:0] tdf4_l2_filters_d0;
input  [15:0] tdf4_l2_filters_q0;
output   tdf4_l2_filters_we0;
output  [10:0] tdf4_l2_filters_address1;
output   tdf4_l2_filters_ce1;
output  [15:0] tdf4_l2_filters_d1;
input  [15:0] tdf4_l2_filters_q1;
output   tdf4_l2_filters_we1;
output  [14:0] tdf5_filters_address0;
output   tdf5_filters_ce0;
output  [15:0] tdf5_filters_d0;
input  [15:0] tdf5_filters_q0;
output   tdf5_filters_we0;
output  [14:0] tdf5_filters_address1;
output   tdf5_filters_ce1;
output  [15:0] tdf5_filters_d1;
input  [15:0] tdf5_filters_q1;
output   tdf5_filters_we1;
output  [11:0] tdf6_filters_address0;
output   tdf6_filters_ce0;
output  [15:0] tdf6_filters_d0;
input  [15:0] tdf6_filters_q0;
output   tdf6_filters_we0;
output  [11:0] tdf6_filters_address1;
output   tdf6_filters_ce1;
output  [15:0] tdf6_filters_d1;
input  [15:0] tdf6_filters_q1;
output   tdf6_filters_we1;
output  [16:0] tdf7_filters_address0;
output   tdf7_filters_ce0;
output  [15:0] tdf7_filters_d0;
input  [15:0] tdf7_filters_q0;
output   tdf7_filters_we0;
output  [16:0] tdf7_filters_address1;
output   tdf7_filters_ce1;
output  [15:0] tdf7_filters_d1;
input  [15:0] tdf7_filters_q1;
output   tdf7_filters_we1;
output  [12:0] tdf7_l2_filters_address0;
output   tdf7_l2_filters_ce0;
output  [15:0] tdf7_l2_filters_d0;
input  [15:0] tdf7_l2_filters_q0;
output   tdf7_l2_filters_we0;
output  [12:0] tdf7_l2_filters_address1;
output   tdf7_l2_filters_ce1;
output  [15:0] tdf7_l2_filters_d1;
input  [15:0] tdf7_l2_filters_q1;
output   tdf7_l2_filters_we1;
output  [16:0] tdf8_filters_address0;
output   tdf8_filters_ce0;
output  [15:0] tdf8_filters_d0;
input  [15:0] tdf8_filters_q0;
output   tdf8_filters_we0;
output  [16:0] tdf8_filters_address1;
output   tdf8_filters_ce1;
output  [15:0] tdf8_filters_d1;
input  [15:0] tdf8_filters_q1;
output   tdf8_filters_we1;
output  [13:0] tdf9_filters_address0;
output   tdf9_filters_ce0;
output  [15:0] tdf9_filters_d0;
input  [15:0] tdf9_filters_q0;
output   tdf9_filters_we0;
output  [13:0] tdf9_filters_address1;
output   tdf9_filters_ce1;
output  [15:0] tdf9_filters_d1;
input  [15:0] tdf9_filters_q1;
output   tdf9_filters_we1;
output  [16:0] tdf10_filters_address0;
output   tdf10_filters_ce0;
output  [63:0] tdf10_filters_d0;
input  [63:0] tdf10_filters_q0;
output   tdf10_filters_we0;
output  [16:0] tdf10_filters_address1;
output   tdf10_filters_ce1;
output  [63:0] tdf10_filters_d1;
input  [63:0] tdf10_filters_q1;
output   tdf10_filters_we1;
output  [14:0] tdf10_l2_filters_address0;
output   tdf10_l2_filters_ce0;
output  [15:0] tdf10_l2_filters_d0;
input  [15:0] tdf10_l2_filters_q0;
output   tdf10_l2_filters_we0;
output  [14:0] tdf10_l2_filters_address1;
output   tdf10_l2_filters_ce1;
output  [15:0] tdf10_l2_filters_d1;
input  [15:0] tdf10_l2_filters_q1;
output   tdf10_l2_filters_we1;
output  [16:0] tdf11_filters_address0;
output   tdf11_filters_ce0;
output  [63:0] tdf11_filters_d0;
input  [63:0] tdf11_filters_q0;
output   tdf11_filters_we0;
output  [16:0] tdf11_filters_address1;
output   tdf11_filters_ce1;
output  [63:0] tdf11_filters_d1;
input  [63:0] tdf11_filters_q1;
output   tdf11_filters_we1;
output  [15:0] tdf11_l2_filters_address0;
output   tdf11_l2_filters_ce0;
output  [15:0] tdf11_l2_filters_d0;
input  [15:0] tdf11_l2_filters_q0;
output   tdf11_l2_filters_we0;
output  [15:0] tdf11_l2_filters_address1;
output   tdf11_l2_filters_ce1;
output  [15:0] tdf11_l2_filters_d1;
input  [15:0] tdf11_l2_filters_q1;
output   tdf11_l2_filters_we1;
output  [16:0] tdf12_filters_address0;
output   tdf12_filters_ce0;
output  [15:0] tdf12_filters_d0;
input  [15:0] tdf12_filters_q0;
output   tdf12_filters_we0;
output  [16:0] tdf12_filters_address1;
output   tdf12_filters_ce1;
output  [15:0] tdf12_filters_d1;
input  [15:0] tdf12_filters_q1;
output   tdf12_filters_we1;
output  [3:0] tdf1_adjustments_address0;
output   tdf1_adjustments_ce0;
output  [47:0] tdf1_adjustments_d0;
input  [47:0] tdf1_adjustments_q0;
output   tdf1_adjustments_we0;
output  [3:0] tdf1_adjustments_address1;
output   tdf1_adjustments_ce1;
output  [47:0] tdf1_adjustments_d1;
input  [47:0] tdf1_adjustments_q1;
output   tdf1_adjustments_we1;
output  [4:0] tdf2_adjustments_address0;
output   tdf2_adjustments_ce0;
output  [47:0] tdf2_adjustments_d0;
input  [47:0] tdf2_adjustments_q0;
output   tdf2_adjustments_we0;
output  [4:0] tdf2_adjustments_address1;
output   tdf2_adjustments_ce1;
output  [47:0] tdf2_adjustments_d1;
input  [47:0] tdf2_adjustments_q1;
output   tdf2_adjustments_we1;
output  [3:0] tdf3_adjustments_address0;
output   tdf3_adjustments_ce0;
output  [47:0] tdf3_adjustments_d0;
input  [47:0] tdf3_adjustments_q0;
output   tdf3_adjustments_we0;
output  [3:0] tdf3_adjustments_address1;
output   tdf3_adjustments_ce1;
output  [47:0] tdf3_adjustments_d1;
input  [47:0] tdf3_adjustments_q1;
output   tdf3_adjustments_we1;
output  [6:0] tdf4_adjustments_address0;
output   tdf4_adjustments_ce0;
output  [47:0] tdf4_adjustments_d0;
input  [47:0] tdf4_adjustments_q0;
output   tdf4_adjustments_we0;
output  [6:0] tdf4_adjustments_address1;
output   tdf4_adjustments_ce1;
output  [47:0] tdf4_adjustments_d1;
input  [47:0] tdf4_adjustments_q1;
output   tdf4_adjustments_we1;
output  [3:0] tdf4_l2_adjustments_address0;
output   tdf4_l2_adjustments_ce0;
output  [47:0] tdf4_l2_adjustments_d0;
input  [47:0] tdf4_l2_adjustments_q0;
output   tdf4_l2_adjustments_we0;
output  [3:0] tdf4_l2_adjustments_address1;
output   tdf4_l2_adjustments_ce1;
output  [47:0] tdf4_l2_adjustments_d1;
input  [47:0] tdf4_l2_adjustments_q1;
output   tdf4_l2_adjustments_we1;
output  [6:0] tdf5_adjustments_address0;
output   tdf5_adjustments_ce0;
output  [47:0] tdf5_adjustments_d0;
input  [47:0] tdf5_adjustments_q0;
output   tdf5_adjustments_we0;
output  [6:0] tdf5_adjustments_address1;
output   tdf5_adjustments_ce1;
output  [47:0] tdf5_adjustments_d1;
input  [47:0] tdf5_adjustments_q1;
output   tdf5_adjustments_we1;
output  [4:0] tdf6_adjustments_address0;
output   tdf6_adjustments_ce0;
output  [47:0] tdf6_adjustments_d0;
input  [47:0] tdf6_adjustments_q0;
output   tdf6_adjustments_we0;
output  [4:0] tdf6_adjustments_address1;
output   tdf6_adjustments_ce1;
output  [47:0] tdf6_adjustments_d1;
input  [47:0] tdf6_adjustments_q1;
output   tdf6_adjustments_we1;
output  [7:0] tdf7_adjustments_address0;
output   tdf7_adjustments_ce0;
output  [47:0] tdf7_adjustments_d0;
input  [47:0] tdf7_adjustments_q0;
output   tdf7_adjustments_we0;
output  [7:0] tdf7_adjustments_address1;
output   tdf7_adjustments_ce1;
output  [47:0] tdf7_adjustments_d1;
input  [47:0] tdf7_adjustments_q1;
output   tdf7_adjustments_we1;
output  [4:0] tdf7_l2_adjustments_address0;
output   tdf7_l2_adjustments_ce0;
output  [47:0] tdf7_l2_adjustments_d0;
input  [47:0] tdf7_l2_adjustments_q0;
output   tdf7_l2_adjustments_we0;
output  [4:0] tdf7_l2_adjustments_address1;
output   tdf7_l2_adjustments_ce1;
output  [47:0] tdf7_l2_adjustments_d1;
input  [47:0] tdf7_l2_adjustments_q1;
output   tdf7_l2_adjustments_we1;
output  [7:0] tdf8_adjustments_address0;
output   tdf8_adjustments_ce0;
output  [47:0] tdf8_adjustments_d0;
input  [47:0] tdf8_adjustments_q0;
output   tdf8_adjustments_we0;
output  [7:0] tdf8_adjustments_address1;
output   tdf8_adjustments_ce1;
output  [47:0] tdf8_adjustments_d1;
input  [47:0] tdf8_adjustments_q1;
output   tdf8_adjustments_we1;
output  [5:0] tdf9_adjustments_address0;
output   tdf9_adjustments_ce0;
output  [47:0] tdf9_adjustments_d0;
input  [47:0] tdf9_adjustments_q0;
output   tdf9_adjustments_we0;
output  [5:0] tdf9_adjustments_address1;
output   tdf9_adjustments_ce1;
output  [47:0] tdf9_adjustments_d1;
input  [47:0] tdf9_adjustments_q1;
output   tdf9_adjustments_we1;
output  [8:0] tdf10_adjustments_address0;
output   tdf10_adjustments_ce0;
output  [47:0] tdf10_adjustments_d0;
input  [47:0] tdf10_adjustments_q0;
output   tdf10_adjustments_we0;
output  [8:0] tdf10_adjustments_address1;
output   tdf10_adjustments_ce1;
output  [47:0] tdf10_adjustments_d1;
input  [47:0] tdf10_adjustments_q1;
output   tdf10_adjustments_we1;
output  [5:0] tdf10_l2_adjustments_address0;
output   tdf10_l2_adjustments_ce0;
output  [47:0] tdf10_l2_adjustments_d0;
input  [47:0] tdf10_l2_adjustments_q0;
output   tdf10_l2_adjustments_we0;
output  [5:0] tdf10_l2_adjustments_address1;
output   tdf10_l2_adjustments_ce1;
output  [47:0] tdf10_l2_adjustments_d1;
input  [47:0] tdf10_l2_adjustments_q1;
output   tdf10_l2_adjustments_we1;
output  [8:0] tdf11_adjustments_address0;
output   tdf11_adjustments_ce0;
output  [47:0] tdf11_adjustments_d0;
input  [47:0] tdf11_adjustments_q0;
output   tdf11_adjustments_we0;
output  [8:0] tdf11_adjustments_address1;
output   tdf11_adjustments_ce1;
output  [47:0] tdf11_adjustments_d1;
input  [47:0] tdf11_adjustments_q1;
output   tdf11_adjustments_we1;
output  [6:0] tdf11_l2_adjustments_address0;
output   tdf11_l2_adjustments_ce0;
output  [47:0] tdf11_l2_adjustments_d0;
input  [47:0] tdf11_l2_adjustments_q0;
output   tdf11_l2_adjustments_we0;
output  [6:0] tdf11_l2_adjustments_address1;
output   tdf11_l2_adjustments_ce1;
output  [47:0] tdf11_l2_adjustments_d1;
input  [47:0] tdf11_l2_adjustments_q1;
output   tdf11_l2_adjustments_we1;
output  [9:0] tdf12_adjustments_address0;
output   tdf12_adjustments_ce0;
output  [47:0] tdf12_adjustments_d0;
input  [47:0] tdf12_adjustments_q0;
output   tdf12_adjustments_we0;
output  [9:0] tdf12_adjustments_address1;
output   tdf12_adjustments_ce1;
output  [47:0] tdf12_adjustments_d1;
input  [47:0] tdf12_adjustments_q1;
output   tdf12_adjustments_we1;
input  [15:0] stream_in_TDATA;
input  [1:0] stream_in_TKEEP;
input  [1:0] stream_in_TSTRB;
input  [0:0] stream_in_TLAST;
output  [15:0] stream_out_TDATA;
output  [1:0] stream_out_TKEEP;
output  [1:0] stream_out_TSTRB;
output  [0:0] stream_out_TLAST;
input   stream_in_TVALID;
output   stream_in_TREADY;
input   ap_start;
output   stream_out_TVALID;
input   stream_out_TREADY;
output   ap_done;
output   ap_ready;
output   ap_idle;
input   ap_continue;

wire   [63:0] tdf1_fmaps_i_q0;
wire   [63:0] tdf1_fmaps_t_q0;
wire   [63:0] tdf2_fmaps_i_q0;
wire   [63:0] tdf2_fmaps_t_q0;
wire   [63:0] tdf3_fmaps_i_q0;
wire   [63:0] tdf3_fmaps_t_q0;
wire   [63:0] tdf4_fmaps_i_q0;
wire   [63:0] tdf4_fmaps_t_q0;
wire   [63:0] tdf5_fmaps_i_q0;
wire   [63:0] tdf5_fmaps_t_q0;
wire   [63:0] tdf6_fmaps_i_q0;
wire   [63:0] tdf6_fmaps_t_q0;
wire   [63:0] tdf7_fmaps_i_q0;
wire   [63:0] tdf7_fmaps_t_q0;
wire   [63:0] tdf8_fmaps_i_q0;
wire   [63:0] tdf8_fmaps_t_q0;
wire   [63:0] tdf9_fmaps_i_q0;
wire   [63:0] tdf9_fmaps_t_q0;
wire   [63:0] tdf10_fmaps_i_q0;
wire   [63:0] tdf10_fmaps_t_q0;
wire   [63:0] tdf11_fmaps_i_q0;
wire   [63:0] tdf11_fmaps_t_q0;
wire   [63:0] tdf12_fmaps_i_q0;
wire   [63:0] tdf12_fmaps_t_q0;
wire   [63:0] final_fmaps_i_q0;
wire   [63:0] final_fmaps_t_q0;
wire    td_fused_axi_in_U0_ap_start;
wire    td_fused_axi_in_U0_ap_done;
wire    td_fused_axi_in_U0_ap_continue;
wire    td_fused_axi_in_U0_ap_idle;
wire    td_fused_axi_in_U0_ap_ready;
wire    td_fused_axi_in_U0_stream_in_TREADY;
wire   [15:0] td_fused_axi_in_U0_fmaps_address1;
wire    td_fused_axi_in_U0_fmaps_ce1;
wire    td_fused_axi_in_U0_fmaps_we1;
wire   [63:0] td_fused_axi_in_U0_fmaps_d1;
wire    ap_channel_done_tdf1_fmaps;
wire    td_fused_axi_in_U0_fmaps_full_n;
wire   [15:0] tdf1_114_U0_in_data_address0;
wire    tdf1_114_U0_in_data_ce0;
wire   [63:0] tdf1_114_U0_in_data_d0;
wire    tdf1_114_U0_in_data_we0;
wire   [15:0] tdf1_114_U0_in_data_address1;
wire    tdf1_114_U0_in_data_ce1;
wire   [63:0] tdf1_114_U0_in_data_d1;
wire    tdf1_114_U0_in_data_we1;
wire   [15:0] tdf1_114_U0_out_data_address0;
wire    tdf1_114_U0_out_data_ce0;
wire   [63:0] tdf1_114_U0_out_data_d0;
wire    tdf1_114_U0_out_data_we0;
wire   [15:0] tdf1_114_U0_out_data_address1;
wire    tdf1_114_U0_out_data_ce1;
wire   [63:0] tdf1_114_U0_out_data_d1;
wire    tdf1_114_U0_out_data_we1;
wire   [8:0] tdf1_114_U0_filter_data_address0;
wire    tdf1_114_U0_filter_data_ce0;
wire   [15:0] tdf1_114_U0_filter_data_d0;
wire    tdf1_114_U0_filter_data_we0;
wire   [8:0] tdf1_114_U0_filter_data_address1;
wire    tdf1_114_U0_filter_data_ce1;
wire   [15:0] tdf1_114_U0_filter_data_d1;
wire    tdf1_114_U0_filter_data_we1;
wire   [3:0] tdf1_114_U0_adjustments_address0;
wire    tdf1_114_U0_adjustments_ce0;
wire   [47:0] tdf1_114_U0_adjustments_d0;
wire    tdf1_114_U0_adjustments_we0;
wire   [3:0] tdf1_114_U0_adjustments_address1;
wire    tdf1_114_U0_adjustments_ce1;
wire   [47:0] tdf1_114_U0_adjustments_d1;
wire    tdf1_114_U0_adjustments_we1;
wire    tdf1_114_U0_in_data_read;
wire    tdf1_114_U0_out_data_full_n;
wire    tdf1_114_U0_out_data_write;
wire    tdf1_114_U0_ap_start;
wire    tdf1_114_U0_ap_done;
wire    tdf1_114_U0_ap_ready;
wire    tdf1_114_U0_ap_idle;
wire    tdf1_114_U0_ap_continue;
wire    ap_channel_done_tdf2_fmaps;
wire   [15:0] tdf2_113_U0_in_data_address0;
wire    tdf2_113_U0_in_data_ce0;
wire   [63:0] tdf2_113_U0_in_data_d0;
wire    tdf2_113_U0_in_data_we0;
wire   [15:0] tdf2_113_U0_in_data_address1;
wire    tdf2_113_U0_in_data_ce1;
wire   [63:0] tdf2_113_U0_in_data_d1;
wire    tdf2_113_U0_in_data_we1;
wire   [14:0] tdf2_113_U0_out_data_address0;
wire    tdf2_113_U0_out_data_ce0;
wire   [63:0] tdf2_113_U0_out_data_d0;
wire    tdf2_113_U0_out_data_we0;
wire   [14:0] tdf2_113_U0_out_data_address1;
wire    tdf2_113_U0_out_data_ce1;
wire   [63:0] tdf2_113_U0_out_data_d1;
wire    tdf2_113_U0_out_data_we1;
wire   [12:0] tdf2_113_U0_filter_data_address0;
wire    tdf2_113_U0_filter_data_ce0;
wire   [15:0] tdf2_113_U0_filter_data_d0;
wire    tdf2_113_U0_filter_data_we0;
wire   [12:0] tdf2_113_U0_filter_data_address1;
wire    tdf2_113_U0_filter_data_ce1;
wire   [15:0] tdf2_113_U0_filter_data_d1;
wire    tdf2_113_U0_filter_data_we1;
wire   [4:0] tdf2_113_U0_adjustments_address0;
wire    tdf2_113_U0_adjustments_ce0;
wire   [47:0] tdf2_113_U0_adjustments_d0;
wire    tdf2_113_U0_adjustments_we0;
wire   [4:0] tdf2_113_U0_adjustments_address1;
wire    tdf2_113_U0_adjustments_ce1;
wire   [47:0] tdf2_113_U0_adjustments_d1;
wire    tdf2_113_U0_adjustments_we1;
wire    tdf2_113_U0_in_data_read;
wire    tdf2_113_U0_out_data_full_n;
wire    tdf2_113_U0_out_data_write;
wire    tdf2_113_U0_ap_start;
wire    tdf2_113_U0_ap_done;
wire    tdf2_113_U0_ap_ready;
wire    tdf2_113_U0_ap_idle;
wire    tdf2_113_U0_ap_continue;
wire    ap_channel_done_tdf3_fmaps;
wire   [14:0] tdf3_112_U0_in_data_address0;
wire    tdf3_112_U0_in_data_ce0;
wire   [63:0] tdf3_112_U0_in_data_d0;
wire    tdf3_112_U0_in_data_we0;
wire   [14:0] tdf3_112_U0_in_data_address1;
wire    tdf3_112_U0_in_data_ce1;
wire   [63:0] tdf3_112_U0_in_data_d1;
wire    tdf3_112_U0_in_data_we1;
wire   [13:0] tdf3_112_U0_out_data_address0;
wire    tdf3_112_U0_out_data_ce0;
wire   [63:0] tdf3_112_U0_out_data_d0;
wire    tdf3_112_U0_out_data_we0;
wire   [13:0] tdf3_112_U0_out_data_address1;
wire    tdf3_112_U0_out_data_ce1;
wire   [63:0] tdf3_112_U0_out_data_d1;
wire    tdf3_112_U0_out_data_we1;
wire   [8:0] tdf3_112_U0_filter_data_address0;
wire    tdf3_112_U0_filter_data_ce0;
wire   [15:0] tdf3_112_U0_filter_data_d0;
wire    tdf3_112_U0_filter_data_we0;
wire   [8:0] tdf3_112_U0_filter_data_address1;
wire    tdf3_112_U0_filter_data_ce1;
wire   [15:0] tdf3_112_U0_filter_data_d1;
wire    tdf3_112_U0_filter_data_we1;
wire   [3:0] tdf3_112_U0_adjustments_address0;
wire    tdf3_112_U0_adjustments_ce0;
wire   [47:0] tdf3_112_U0_adjustments_d0;
wire    tdf3_112_U0_adjustments_we0;
wire   [3:0] tdf3_112_U0_adjustments_address1;
wire    tdf3_112_U0_adjustments_ce1;
wire   [47:0] tdf3_112_U0_adjustments_d1;
wire    tdf3_112_U0_adjustments_we1;
wire    tdf3_112_U0_in_data_read;
wire    tdf3_112_U0_out_data_full_n;
wire    tdf3_112_U0_out_data_write;
wire    tdf3_112_U0_ap_start;
wire    tdf3_112_U0_ap_done;
wire    tdf3_112_U0_ap_ready;
wire    tdf3_112_U0_ap_idle;
wire    tdf3_112_U0_ap_continue;
wire    ap_channel_done_tdf4_fmaps;
wire   [13:0] tdf4_111_U0_in_data_address0;
wire    tdf4_111_U0_in_data_ce0;
wire   [63:0] tdf4_111_U0_in_data_d0;
wire    tdf4_111_U0_in_data_we0;
wire   [13:0] tdf4_111_U0_in_data_address1;
wire    tdf4_111_U0_in_data_ce1;
wire   [63:0] tdf4_111_U0_in_data_d1;
wire    tdf4_111_U0_in_data_we1;
wire   [13:0] tdf4_111_U0_out_data_address0;
wire    tdf4_111_U0_out_data_ce0;
wire   [63:0] tdf4_111_U0_out_data_d0;
wire    tdf4_111_U0_out_data_we0;
wire   [13:0] tdf4_111_U0_out_data_address1;
wire    tdf4_111_U0_out_data_ce1;
wire   [63:0] tdf4_111_U0_out_data_d1;
wire    tdf4_111_U0_out_data_we1;
wire   [14:0] tdf4_111_U0_l1_filter_data_address0;
wire    tdf4_111_U0_l1_filter_data_ce0;
wire   [15:0] tdf4_111_U0_l1_filter_data_d0;
wire    tdf4_111_U0_l1_filter_data_we0;
wire   [14:0] tdf4_111_U0_l1_filter_data_address1;
wire    tdf4_111_U0_l1_filter_data_ce1;
wire   [15:0] tdf4_111_U0_l1_filter_data_d1;
wire    tdf4_111_U0_l1_filter_data_we1;
wire   [10:0] tdf4_111_U0_l2_filter_data_address0;
wire    tdf4_111_U0_l2_filter_data_ce0;
wire   [15:0] tdf4_111_U0_l2_filter_data_d0;
wire    tdf4_111_U0_l2_filter_data_we0;
wire   [10:0] tdf4_111_U0_l2_filter_data_address1;
wire    tdf4_111_U0_l2_filter_data_ce1;
wire   [15:0] tdf4_111_U0_l2_filter_data_d1;
wire    tdf4_111_U0_l2_filter_data_we1;
wire   [6:0] tdf4_111_U0_l1_adjustments_address0;
wire    tdf4_111_U0_l1_adjustments_ce0;
wire   [47:0] tdf4_111_U0_l1_adjustments_d0;
wire    tdf4_111_U0_l1_adjustments_we0;
wire   [6:0] tdf4_111_U0_l1_adjustments_address1;
wire    tdf4_111_U0_l1_adjustments_ce1;
wire   [47:0] tdf4_111_U0_l1_adjustments_d1;
wire    tdf4_111_U0_l1_adjustments_we1;
wire   [3:0] tdf4_111_U0_l2_adjustments_address0;
wire    tdf4_111_U0_l2_adjustments_ce0;
wire   [47:0] tdf4_111_U0_l2_adjustments_d0;
wire    tdf4_111_U0_l2_adjustments_we0;
wire   [3:0] tdf4_111_U0_l2_adjustments_address1;
wire    tdf4_111_U0_l2_adjustments_ce1;
wire   [47:0] tdf4_111_U0_l2_adjustments_d1;
wire    tdf4_111_U0_l2_adjustments_we1;
wire    tdf4_111_U0_in_data_read;
wire    tdf4_111_U0_out_data_full_n;
wire    tdf4_111_U0_out_data_write;
wire    tdf4_111_U0_ap_start;
wire    tdf4_111_U0_ap_done;
wire    tdf4_111_U0_ap_ready;
wire    tdf4_111_U0_ap_idle;
wire    tdf4_111_U0_ap_continue;
wire    ap_channel_done_tdf5_fmaps;
wire   [13:0] tdf5_110_U0_in_data_address0;
wire    tdf5_110_U0_in_data_ce0;
wire   [63:0] tdf5_110_U0_in_data_d0;
wire    tdf5_110_U0_in_data_we0;
wire   [13:0] tdf5_110_U0_in_data_address1;
wire    tdf5_110_U0_in_data_ce1;
wire   [63:0] tdf5_110_U0_in_data_d1;
wire    tdf5_110_U0_in_data_we1;
wire   [14:0] tdf5_110_U0_out_data_address0;
wire    tdf5_110_U0_out_data_ce0;
wire   [63:0] tdf5_110_U0_out_data_d0;
wire    tdf5_110_U0_out_data_we0;
wire   [14:0] tdf5_110_U0_out_data_address1;
wire    tdf5_110_U0_out_data_ce1;
wire   [63:0] tdf5_110_U0_out_data_d1;
wire    tdf5_110_U0_out_data_we1;
wire   [14:0] tdf5_110_U0_filter_data_address0;
wire    tdf5_110_U0_filter_data_ce0;
wire   [15:0] tdf5_110_U0_filter_data_d0;
wire    tdf5_110_U0_filter_data_we0;
wire   [14:0] tdf5_110_U0_filter_data_address1;
wire    tdf5_110_U0_filter_data_ce1;
wire   [15:0] tdf5_110_U0_filter_data_d1;
wire    tdf5_110_U0_filter_data_we1;
wire   [6:0] tdf5_110_U0_adjustments_address0;
wire    tdf5_110_U0_adjustments_ce0;
wire   [47:0] tdf5_110_U0_adjustments_d0;
wire    tdf5_110_U0_adjustments_we0;
wire   [6:0] tdf5_110_U0_adjustments_address1;
wire    tdf5_110_U0_adjustments_ce1;
wire   [47:0] tdf5_110_U0_adjustments_d1;
wire    tdf5_110_U0_adjustments_we1;
wire    tdf5_110_U0_in_data_read;
wire    tdf5_110_U0_out_data_full_n;
wire    tdf5_110_U0_out_data_write;
wire    tdf5_110_U0_ap_start;
wire    tdf5_110_U0_ap_done;
wire    tdf5_110_U0_ap_ready;
wire    tdf5_110_U0_ap_idle;
wire    tdf5_110_U0_ap_continue;
wire    ap_channel_done_tdf6_fmaps;
wire   [14:0] tdf6_19_U0_in_data_address0;
wire    tdf6_19_U0_in_data_ce0;
wire   [63:0] tdf6_19_U0_in_data_d0;
wire    tdf6_19_U0_in_data_we0;
wire   [14:0] tdf6_19_U0_in_data_address1;
wire    tdf6_19_U0_in_data_ce1;
wire   [63:0] tdf6_19_U0_in_data_d1;
wire    tdf6_19_U0_in_data_we1;
wire   [12:0] tdf6_19_U0_out_data_address0;
wire    tdf6_19_U0_out_data_ce0;
wire   [63:0] tdf6_19_U0_out_data_d0;
wire    tdf6_19_U0_out_data_we0;
wire   [12:0] tdf6_19_U0_out_data_address1;
wire    tdf6_19_U0_out_data_ce1;
wire   [63:0] tdf6_19_U0_out_data_d1;
wire    tdf6_19_U0_out_data_we1;
wire   [11:0] tdf6_19_U0_filter_data_address0;
wire    tdf6_19_U0_filter_data_ce0;
wire   [15:0] tdf6_19_U0_filter_data_d0;
wire    tdf6_19_U0_filter_data_we0;
wire   [11:0] tdf6_19_U0_filter_data_address1;
wire    tdf6_19_U0_filter_data_ce1;
wire   [15:0] tdf6_19_U0_filter_data_d1;
wire    tdf6_19_U0_filter_data_we1;
wire   [4:0] tdf6_19_U0_adjustments_address0;
wire    tdf6_19_U0_adjustments_ce0;
wire   [47:0] tdf6_19_U0_adjustments_d0;
wire    tdf6_19_U0_adjustments_we0;
wire   [4:0] tdf6_19_U0_adjustments_address1;
wire    tdf6_19_U0_adjustments_ce1;
wire   [47:0] tdf6_19_U0_adjustments_d1;
wire    tdf6_19_U0_adjustments_we1;
wire    tdf6_19_U0_in_data_read;
wire    tdf6_19_U0_out_data_full_n;
wire    tdf6_19_U0_out_data_write;
wire    tdf6_19_U0_ap_start;
wire    tdf6_19_U0_ap_done;
wire    tdf6_19_U0_ap_ready;
wire    tdf6_19_U0_ap_idle;
wire    tdf6_19_U0_ap_continue;
wire    ap_channel_done_tdf7_fmaps;
wire   [12:0] tdf7_18_U0_in_data_address0;
wire    tdf7_18_U0_in_data_ce0;
wire   [63:0] tdf7_18_U0_in_data_d0;
wire    tdf7_18_U0_in_data_we0;
wire   [12:0] tdf7_18_U0_in_data_address1;
wire    tdf7_18_U0_in_data_ce1;
wire   [63:0] tdf7_18_U0_in_data_d1;
wire    tdf7_18_U0_in_data_we1;
wire   [12:0] tdf7_18_U0_out_data_address0;
wire    tdf7_18_U0_out_data_ce0;
wire   [63:0] tdf7_18_U0_out_data_d0;
wire    tdf7_18_U0_out_data_we0;
wire   [12:0] tdf7_18_U0_out_data_address1;
wire    tdf7_18_U0_out_data_ce1;
wire   [63:0] tdf7_18_U0_out_data_d1;
wire    tdf7_18_U0_out_data_we1;
wire   [16:0] tdf7_18_U0_l1_filter_data_address0;
wire    tdf7_18_U0_l1_filter_data_ce0;
wire   [15:0] tdf7_18_U0_l1_filter_data_d0;
wire    tdf7_18_U0_l1_filter_data_we0;
wire   [16:0] tdf7_18_U0_l1_filter_data_address1;
wire    tdf7_18_U0_l1_filter_data_ce1;
wire   [15:0] tdf7_18_U0_l1_filter_data_d1;
wire    tdf7_18_U0_l1_filter_data_we1;
wire   [12:0] tdf7_18_U0_l2_filter_data_address0;
wire    tdf7_18_U0_l2_filter_data_ce0;
wire   [15:0] tdf7_18_U0_l2_filter_data_d0;
wire    tdf7_18_U0_l2_filter_data_we0;
wire   [12:0] tdf7_18_U0_l2_filter_data_address1;
wire    tdf7_18_U0_l2_filter_data_ce1;
wire   [15:0] tdf7_18_U0_l2_filter_data_d1;
wire    tdf7_18_U0_l2_filter_data_we1;
wire   [7:0] tdf7_18_U0_l1_adjustments_address0;
wire    tdf7_18_U0_l1_adjustments_ce0;
wire   [47:0] tdf7_18_U0_l1_adjustments_d0;
wire    tdf7_18_U0_l1_adjustments_we0;
wire   [7:0] tdf7_18_U0_l1_adjustments_address1;
wire    tdf7_18_U0_l1_adjustments_ce1;
wire   [47:0] tdf7_18_U0_l1_adjustments_d1;
wire    tdf7_18_U0_l1_adjustments_we1;
wire   [4:0] tdf7_18_U0_l2_adjustments_address0;
wire    tdf7_18_U0_l2_adjustments_ce0;
wire   [47:0] tdf7_18_U0_l2_adjustments_d0;
wire    tdf7_18_U0_l2_adjustments_we0;
wire   [4:0] tdf7_18_U0_l2_adjustments_address1;
wire    tdf7_18_U0_l2_adjustments_ce1;
wire   [47:0] tdf7_18_U0_l2_adjustments_d1;
wire    tdf7_18_U0_l2_adjustments_we1;
wire    tdf7_18_U0_in_data_read;
wire    tdf7_18_U0_out_data_full_n;
wire    tdf7_18_U0_out_data_write;
wire    tdf7_18_U0_ap_start;
wire    tdf7_18_U0_ap_done;
wire    tdf7_18_U0_ap_ready;
wire    tdf7_18_U0_ap_idle;
wire    tdf7_18_U0_ap_continue;
wire    ap_channel_done_tdf8_fmaps;
wire   [12:0] tdf8_17_U0_in_data_address0;
wire    tdf8_17_U0_in_data_ce0;
wire   [63:0] tdf8_17_U0_in_data_d0;
wire    tdf8_17_U0_in_data_we0;
wire   [12:0] tdf8_17_U0_in_data_address1;
wire    tdf8_17_U0_in_data_ce1;
wire   [63:0] tdf8_17_U0_in_data_d1;
wire    tdf8_17_U0_in_data_we1;
wire   [13:0] tdf8_17_U0_out_data_address0;
wire    tdf8_17_U0_out_data_ce0;
wire   [63:0] tdf8_17_U0_out_data_d0;
wire    tdf8_17_U0_out_data_we0;
wire   [13:0] tdf8_17_U0_out_data_address1;
wire    tdf8_17_U0_out_data_ce1;
wire   [63:0] tdf8_17_U0_out_data_d1;
wire    tdf8_17_U0_out_data_we1;
wire   [16:0] tdf8_17_U0_filter_data_address0;
wire    tdf8_17_U0_filter_data_ce0;
wire   [15:0] tdf8_17_U0_filter_data_d0;
wire    tdf8_17_U0_filter_data_we0;
wire   [16:0] tdf8_17_U0_filter_data_address1;
wire    tdf8_17_U0_filter_data_ce1;
wire   [15:0] tdf8_17_U0_filter_data_d1;
wire    tdf8_17_U0_filter_data_we1;
wire   [7:0] tdf8_17_U0_adjustments_address0;
wire    tdf8_17_U0_adjustments_ce0;
wire   [47:0] tdf8_17_U0_adjustments_d0;
wire    tdf8_17_U0_adjustments_we0;
wire   [7:0] tdf8_17_U0_adjustments_address1;
wire    tdf8_17_U0_adjustments_ce1;
wire   [47:0] tdf8_17_U0_adjustments_d1;
wire    tdf8_17_U0_adjustments_we1;
wire    tdf8_17_U0_in_data_read;
wire    tdf8_17_U0_out_data_full_n;
wire    tdf8_17_U0_out_data_write;
wire    tdf8_17_U0_ap_start;
wire    tdf8_17_U0_ap_done;
wire    tdf8_17_U0_ap_ready;
wire    tdf8_17_U0_ap_idle;
wire    tdf8_17_U0_ap_continue;
wire    ap_channel_done_tdf9_fmaps;
wire   [13:0] tdf9_16_U0_in_data_address0;
wire    tdf9_16_U0_in_data_ce0;
wire   [63:0] tdf9_16_U0_in_data_d0;
wire    tdf9_16_U0_in_data_we0;
wire   [13:0] tdf9_16_U0_in_data_address1;
wire    tdf9_16_U0_in_data_ce1;
wire   [63:0] tdf9_16_U0_in_data_d1;
wire    tdf9_16_U0_in_data_we1;
wire   [11:0] tdf9_16_U0_out_data_address0;
wire    tdf9_16_U0_out_data_ce0;
wire   [63:0] tdf9_16_U0_out_data_d0;
wire    tdf9_16_U0_out_data_we0;
wire   [11:0] tdf9_16_U0_out_data_address1;
wire    tdf9_16_U0_out_data_ce1;
wire   [63:0] tdf9_16_U0_out_data_d1;
wire    tdf9_16_U0_out_data_we1;
wire   [13:0] tdf9_16_U0_filter_data_address0;
wire    tdf9_16_U0_filter_data_ce0;
wire   [15:0] tdf9_16_U0_filter_data_d0;
wire    tdf9_16_U0_filter_data_we0;
wire   [13:0] tdf9_16_U0_filter_data_address1;
wire    tdf9_16_U0_filter_data_ce1;
wire   [15:0] tdf9_16_U0_filter_data_d1;
wire    tdf9_16_U0_filter_data_we1;
wire   [5:0] tdf9_16_U0_adjustments_address0;
wire    tdf9_16_U0_adjustments_ce0;
wire   [47:0] tdf9_16_U0_adjustments_d0;
wire    tdf9_16_U0_adjustments_we0;
wire   [5:0] tdf9_16_U0_adjustments_address1;
wire    tdf9_16_U0_adjustments_ce1;
wire   [47:0] tdf9_16_U0_adjustments_d1;
wire    tdf9_16_U0_adjustments_we1;
wire    tdf9_16_U0_in_data_read;
wire    tdf9_16_U0_out_data_full_n;
wire    tdf9_16_U0_out_data_write;
wire    tdf9_16_U0_ap_start;
wire    tdf9_16_U0_ap_done;
wire    tdf9_16_U0_ap_ready;
wire    tdf9_16_U0_ap_idle;
wire    tdf9_16_U0_ap_continue;
wire    ap_channel_done_tdf10_fmaps;
wire   [11:0] tdf10_15_U0_in_data_address0;
wire    tdf10_15_U0_in_data_ce0;
wire   [63:0] tdf10_15_U0_in_data_d0;
wire    tdf10_15_U0_in_data_we0;
wire   [11:0] tdf10_15_U0_in_data_address1;
wire    tdf10_15_U0_in_data_ce1;
wire   [63:0] tdf10_15_U0_in_data_d1;
wire    tdf10_15_U0_in_data_we1;
wire   [11:0] tdf10_15_U0_out_data_address0;
wire    tdf10_15_U0_out_data_ce0;
wire   [63:0] tdf10_15_U0_out_data_d0;
wire    tdf10_15_U0_out_data_we0;
wire   [11:0] tdf10_15_U0_out_data_address1;
wire    tdf10_15_U0_out_data_ce1;
wire   [63:0] tdf10_15_U0_out_data_d1;
wire    tdf10_15_U0_out_data_we1;
wire   [16:0] tdf10_15_U0_l1_filter_data_address0;
wire    tdf10_15_U0_l1_filter_data_ce0;
wire   [63:0] tdf10_15_U0_l1_filter_data_d0;
wire    tdf10_15_U0_l1_filter_data_we0;
wire   [16:0] tdf10_15_U0_l1_filter_data_address1;
wire    tdf10_15_U0_l1_filter_data_ce1;
wire   [63:0] tdf10_15_U0_l1_filter_data_d1;
wire    tdf10_15_U0_l1_filter_data_we1;
wire   [14:0] tdf10_15_U0_l2_filter_data_address0;
wire    tdf10_15_U0_l2_filter_data_ce0;
wire   [15:0] tdf10_15_U0_l2_filter_data_d0;
wire    tdf10_15_U0_l2_filter_data_we0;
wire   [14:0] tdf10_15_U0_l2_filter_data_address1;
wire    tdf10_15_U0_l2_filter_data_ce1;
wire   [15:0] tdf10_15_U0_l2_filter_data_d1;
wire    tdf10_15_U0_l2_filter_data_we1;
wire   [8:0] tdf10_15_U0_l1_adjustments_address0;
wire    tdf10_15_U0_l1_adjustments_ce0;
wire   [47:0] tdf10_15_U0_l1_adjustments_d0;
wire    tdf10_15_U0_l1_adjustments_we0;
wire   [8:0] tdf10_15_U0_l1_adjustments_address1;
wire    tdf10_15_U0_l1_adjustments_ce1;
wire   [47:0] tdf10_15_U0_l1_adjustments_d1;
wire    tdf10_15_U0_l1_adjustments_we1;
wire   [5:0] tdf10_15_U0_l2_adjustments_address0;
wire    tdf10_15_U0_l2_adjustments_ce0;
wire   [47:0] tdf10_15_U0_l2_adjustments_d0;
wire    tdf10_15_U0_l2_adjustments_we0;
wire   [5:0] tdf10_15_U0_l2_adjustments_address1;
wire    tdf10_15_U0_l2_adjustments_ce1;
wire   [47:0] tdf10_15_U0_l2_adjustments_d1;
wire    tdf10_15_U0_l2_adjustments_we1;
wire    tdf10_15_U0_in_data_read;
wire    tdf10_15_U0_out_data_full_n;
wire    tdf10_15_U0_out_data_write;
wire    tdf10_15_U0_ap_start;
wire    tdf10_15_U0_ap_done;
wire    tdf10_15_U0_ap_ready;
wire    tdf10_15_U0_ap_idle;
wire    tdf10_15_U0_ap_continue;
wire    ap_channel_done_tdf11_fmaps;
wire   [11:0] tdf11_14_U0_in_data_address0;
wire    tdf11_14_U0_in_data_ce0;
wire   [63:0] tdf11_14_U0_in_data_d0;
wire    tdf11_14_U0_in_data_we0;
wire   [11:0] tdf11_14_U0_in_data_address1;
wire    tdf11_14_U0_in_data_ce1;
wire   [63:0] tdf11_14_U0_in_data_d1;
wire    tdf11_14_U0_in_data_we1;
wire   [12:0] tdf11_14_U0_out_data_address0;
wire    tdf11_14_U0_out_data_ce0;
wire   [63:0] tdf11_14_U0_out_data_d0;
wire    tdf11_14_U0_out_data_we0;
wire   [12:0] tdf11_14_U0_out_data_address1;
wire    tdf11_14_U0_out_data_ce1;
wire   [63:0] tdf11_14_U0_out_data_d1;
wire    tdf11_14_U0_out_data_we1;
wire   [16:0] tdf11_14_U0_l1_filter_data_address0;
wire    tdf11_14_U0_l1_filter_data_ce0;
wire   [63:0] tdf11_14_U0_l1_filter_data_d0;
wire    tdf11_14_U0_l1_filter_data_we0;
wire   [16:0] tdf11_14_U0_l1_filter_data_address1;
wire    tdf11_14_U0_l1_filter_data_ce1;
wire   [63:0] tdf11_14_U0_l1_filter_data_d1;
wire    tdf11_14_U0_l1_filter_data_we1;
wire   [15:0] tdf11_14_U0_l2_filter_data_address0;
wire    tdf11_14_U0_l2_filter_data_ce0;
wire   [15:0] tdf11_14_U0_l2_filter_data_d0;
wire    tdf11_14_U0_l2_filter_data_we0;
wire   [15:0] tdf11_14_U0_l2_filter_data_address1;
wire    tdf11_14_U0_l2_filter_data_ce1;
wire   [15:0] tdf11_14_U0_l2_filter_data_d1;
wire    tdf11_14_U0_l2_filter_data_we1;
wire   [8:0] tdf11_14_U0_l1_adjustments_address0;
wire    tdf11_14_U0_l1_adjustments_ce0;
wire   [47:0] tdf11_14_U0_l1_adjustments_d0;
wire    tdf11_14_U0_l1_adjustments_we0;
wire   [8:0] tdf11_14_U0_l1_adjustments_address1;
wire    tdf11_14_U0_l1_adjustments_ce1;
wire   [47:0] tdf11_14_U0_l1_adjustments_d1;
wire    tdf11_14_U0_l1_adjustments_we1;
wire   [6:0] tdf11_14_U0_l2_adjustments_address0;
wire    tdf11_14_U0_l2_adjustments_ce0;
wire   [47:0] tdf11_14_U0_l2_adjustments_d0;
wire    tdf11_14_U0_l2_adjustments_we0;
wire   [6:0] tdf11_14_U0_l2_adjustments_address1;
wire    tdf11_14_U0_l2_adjustments_ce1;
wire   [47:0] tdf11_14_U0_l2_adjustments_d1;
wire    tdf11_14_U0_l2_adjustments_we1;
wire    tdf11_14_U0_in_data_read;
wire    tdf11_14_U0_out_data_full_n;
wire    tdf11_14_U0_out_data_write;
wire    tdf11_14_U0_ap_start;
wire    tdf11_14_U0_ap_done;
wire    tdf11_14_U0_ap_ready;
wire    tdf11_14_U0_ap_idle;
wire    tdf11_14_U0_ap_continue;
wire    ap_channel_done_tdf12_fmaps;
wire   [12:0] tdf12_13_U0_in_data_address0;
wire    tdf12_13_U0_in_data_ce0;
wire   [63:0] tdf12_13_U0_in_data_d0;
wire    tdf12_13_U0_in_data_we0;
wire   [12:0] tdf12_13_U0_in_data_address1;
wire    tdf12_13_U0_in_data_ce1;
wire   [63:0] tdf12_13_U0_in_data_d1;
wire    tdf12_13_U0_in_data_we1;
wire   [15:0] tdf12_13_U0_out_data_address0;
wire    tdf12_13_U0_out_data_ce0;
wire   [63:0] tdf12_13_U0_out_data_d0;
wire    tdf12_13_U0_out_data_we0;
wire   [15:0] tdf12_13_U0_out_data_address1;
wire    tdf12_13_U0_out_data_ce1;
wire   [63:0] tdf12_13_U0_out_data_d1;
wire    tdf12_13_U0_out_data_we1;
wire   [16:0] tdf12_13_U0_filter_data_address0;
wire    tdf12_13_U0_filter_data_ce0;
wire   [15:0] tdf12_13_U0_filter_data_d0;
wire    tdf12_13_U0_filter_data_we0;
wire   [16:0] tdf12_13_U0_filter_data_address1;
wire    tdf12_13_U0_filter_data_ce1;
wire   [15:0] tdf12_13_U0_filter_data_d1;
wire    tdf12_13_U0_filter_data_we1;
wire   [9:0] tdf12_13_U0_adjustments_address0;
wire    tdf12_13_U0_adjustments_ce0;
wire   [47:0] tdf12_13_U0_adjustments_d0;
wire    tdf12_13_U0_adjustments_we0;
wire   [9:0] tdf12_13_U0_adjustments_address1;
wire    tdf12_13_U0_adjustments_ce1;
wire   [47:0] tdf12_13_U0_adjustments_d1;
wire    tdf12_13_U0_adjustments_we1;
wire    tdf12_13_U0_in_data_read;
wire    tdf12_13_U0_out_data_full_n;
wire    tdf12_13_U0_out_data_write;
wire    tdf12_13_U0_ap_start;
wire    tdf12_13_U0_ap_done;
wire    tdf12_13_U0_ap_ready;
wire    tdf12_13_U0_ap_idle;
wire    tdf12_13_U0_ap_continue;
wire    ap_channel_done_final_fmaps;
wire    td_fused_axi_out_U0_ap_start;
wire    td_fused_axi_out_U0_ap_done;
wire    td_fused_axi_out_U0_ap_continue;
wire    td_fused_axi_out_U0_ap_idle;
wire    td_fused_axi_out_U0_ap_ready;
wire   [15:0] td_fused_axi_out_U0_fmaps_address0;
wire    td_fused_axi_out_U0_fmaps_ce0;
wire   [15:0] td_fused_axi_out_U0_stream_out_TDATA;
wire    td_fused_axi_out_U0_stream_out_TVALID;
wire   [1:0] td_fused_axi_out_U0_stream_out_TKEEP;
wire   [1:0] td_fused_axi_out_U0_stream_out_TSTRB;
wire   [0:0] td_fused_axi_out_U0_stream_out_TLAST;
wire    ap_sync_continue;
wire    tdf1_fmaps_i_full_n;
wire    tdf1_fmaps_t_empty_n;
wire   [63:0] tdf1_fmaps_t_d0;
wire    tdf1_fmaps_t_we0;
wire    tdf2_fmaps_i_full_n;
wire    tdf2_fmaps_t_empty_n;
wire   [63:0] tdf2_fmaps_t_d0;
wire    tdf2_fmaps_t_we0;
wire    tdf3_fmaps_i_full_n;
wire    tdf3_fmaps_t_empty_n;
wire   [63:0] tdf3_fmaps_t_d0;
wire    tdf3_fmaps_t_we0;
wire    tdf4_fmaps_i_full_n;
wire    tdf4_fmaps_t_empty_n;
wire   [63:0] tdf4_fmaps_t_d0;
wire    tdf4_fmaps_t_we0;
wire    tdf5_fmaps_i_full_n;
wire    tdf5_fmaps_t_empty_n;
wire   [63:0] tdf5_fmaps_t_d0;
wire    tdf5_fmaps_t_we0;
wire    tdf6_fmaps_i_full_n;
wire    tdf6_fmaps_t_empty_n;
wire   [63:0] tdf6_fmaps_t_d0;
wire    tdf6_fmaps_t_we0;
wire    tdf7_fmaps_i_full_n;
wire    tdf7_fmaps_t_empty_n;
wire   [63:0] tdf7_fmaps_t_d0;
wire    tdf7_fmaps_t_we0;
wire    tdf8_fmaps_i_full_n;
wire    tdf8_fmaps_t_empty_n;
wire   [63:0] tdf8_fmaps_t_d0;
wire    tdf8_fmaps_t_we0;
wire    tdf9_fmaps_i_full_n;
wire    tdf9_fmaps_t_empty_n;
wire   [63:0] tdf9_fmaps_t_d0;
wire    tdf9_fmaps_t_we0;
wire    tdf10_fmaps_i_full_n;
wire    tdf10_fmaps_t_empty_n;
wire   [63:0] tdf10_fmaps_t_d0;
wire    tdf10_fmaps_t_we0;
wire    tdf11_fmaps_i_full_n;
wire    tdf11_fmaps_t_empty_n;
wire   [63:0] tdf11_fmaps_t_d0;
wire    tdf11_fmaps_t_we0;
wire    tdf12_fmaps_i_full_n;
wire    tdf12_fmaps_t_empty_n;
wire   [63:0] tdf12_fmaps_t_d0;
wire    tdf12_fmaps_t_we0;
wire    final_fmaps_i_full_n;
wire    final_fmaps_t_empty_n;
wire   [63:0] final_fmaps_t_d0;
wire    final_fmaps_t_we0;
wire    ap_sync_done;
wire    ap_sync_ready;
wire    td_fused_axi_in_U0_start_full_n;
wire    td_fused_axi_in_U0_start_write;
wire    tdf1_114_U0_start_full_n;
wire    tdf1_114_U0_start_write;
wire    tdf2_113_U0_start_full_n;
wire    tdf2_113_U0_start_write;
wire    tdf3_112_U0_start_full_n;
wire    tdf3_112_U0_start_write;
wire    tdf4_111_U0_start_full_n;
wire    tdf4_111_U0_start_write;
wire    tdf5_110_U0_start_full_n;
wire    tdf5_110_U0_start_write;
wire    tdf6_19_U0_start_full_n;
wire    tdf6_19_U0_start_write;
wire    tdf7_18_U0_start_full_n;
wire    tdf7_18_U0_start_write;
wire    tdf8_17_U0_start_full_n;
wire    tdf8_17_U0_start_write;
wire    tdf9_16_U0_start_full_n;
wire    tdf9_16_U0_start_write;
wire    tdf10_15_U0_start_full_n;
wire    tdf10_15_U0_start_write;
wire    tdf11_14_U0_start_full_n;
wire    tdf11_14_U0_start_write;
wire    tdf12_13_U0_start_full_n;
wire    tdf12_13_U0_start_write;
wire    td_fused_axi_out_U0_start_full_n;
wire    td_fused_axi_out_U0_start_write;

td_fused_top_td_fused_tdf1_fmaps #(
    .DataWidth( 64 ),
    .AddressRange( 50176 ),
    .AddressWidth( 16 ))
tdf1_fmaps_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(td_fused_axi_in_U0_ap_done),
    .i_full_n(tdf1_fmaps_i_full_n),
    .i_ce0(1'b0),
    .i_address0(16'd0),
    .i_q0(tdf1_fmaps_i_q0),
    .i_ce1(td_fused_axi_in_U0_fmaps_ce1),
    .i_we1(td_fused_axi_in_U0_fmaps_we1),
    .i_address1(td_fused_axi_in_U0_fmaps_address1),
    .i_d1(td_fused_axi_in_U0_fmaps_d1),
    .t_ce(1'b1),
    .t_read(tdf1_114_U0_ap_ready),
    .t_empty_n(tdf1_fmaps_t_empty_n),
    .t_ce0(tdf1_114_U0_in_data_ce0),
    .t_address0(tdf1_114_U0_in_data_address0),
    .t_q0(tdf1_fmaps_t_q0),
    .t_ce1(1'b0),
    .t_we1(1'b0),
    .t_address1(16'd0),
    .t_d1(64'd0)
);

td_fused_top_td_fused_tdf1_fmaps #(
    .DataWidth( 64 ),
    .AddressRange( 50176 ),
    .AddressWidth( 16 ))
tdf2_fmaps_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf1_114_U0_ap_done),
    .i_full_n(tdf2_fmaps_i_full_n),
    .i_ce0(1'b0),
    .i_address0(16'd0),
    .i_q0(tdf2_fmaps_i_q0),
    .i_ce1(tdf1_114_U0_out_data_ce1),
    .i_we1(tdf1_114_U0_out_data_we1),
    .i_address1(tdf1_114_U0_out_data_address1),
    .i_d1(tdf1_114_U0_out_data_d1),
    .t_ce(1'b1),
    .t_read(tdf2_113_U0_ap_ready),
    .t_empty_n(tdf2_fmaps_t_empty_n),
    .t_ce0(tdf2_113_U0_in_data_ce0),
    .t_address0(tdf2_113_U0_in_data_address0),
    .t_q0(tdf2_fmaps_t_q0),
    .t_ce1(1'b0),
    .t_we1(1'b0),
    .t_address1(16'd0),
    .t_d1(64'd0)
);

td_fused_top_td_fused_tdf3_fmaps #(
    .DataWidth( 64 ),
    .AddressRange( 25088 ),
    .AddressWidth( 15 ))
tdf3_fmaps_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf2_113_U0_ap_done),
    .i_full_n(tdf3_fmaps_i_full_n),
    .i_ce0(1'b0),
    .i_address0(15'd0),
    .i_q0(tdf3_fmaps_i_q0),
    .i_ce1(tdf2_113_U0_out_data_ce1),
    .i_we1(tdf2_113_U0_out_data_we1),
    .i_address1(tdf2_113_U0_out_data_address1),
    .i_d1(tdf2_113_U0_out_data_d1),
    .t_ce(1'b1),
    .t_read(tdf3_112_U0_ap_ready),
    .t_empty_n(tdf3_fmaps_t_empty_n),
    .t_ce0(tdf3_112_U0_in_data_ce0),
    .t_address0(tdf3_112_U0_in_data_address0),
    .t_q0(tdf3_fmaps_t_q0),
    .t_ce1(1'b0),
    .t_we1(1'b0),
    .t_address1(15'd0),
    .t_d1(64'd0)
);

td_fused_top_td_fused_tdf4_fmaps #(
    .DataWidth( 64 ),
    .AddressRange( 12544 ),
    .AddressWidth( 14 ))
tdf4_fmaps_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf3_112_U0_ap_done),
    .i_full_n(tdf4_fmaps_i_full_n),
    .i_ce0(1'b0),
    .i_address0(14'd0),
    .i_q0(tdf4_fmaps_i_q0),
    .i_ce1(tdf3_112_U0_out_data_ce1),
    .i_we1(tdf3_112_U0_out_data_we1),
    .i_address1(tdf3_112_U0_out_data_address1),
    .i_d1(tdf3_112_U0_out_data_d1),
    .t_ce(1'b1),
    .t_read(tdf4_111_U0_ap_ready),
    .t_empty_n(tdf4_fmaps_t_empty_n),
    .t_ce0(tdf4_111_U0_in_data_ce0),
    .t_address0(tdf4_111_U0_in_data_address0),
    .t_q0(tdf4_fmaps_t_q0),
    .t_ce1(1'b0),
    .t_we1(1'b0),
    .t_address1(14'd0),
    .t_d1(64'd0)
);

td_fused_top_td_fused_tdf4_fmaps #(
    .DataWidth( 64 ),
    .AddressRange( 12544 ),
    .AddressWidth( 14 ))
tdf5_fmaps_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf4_111_U0_ap_done),
    .i_full_n(tdf5_fmaps_i_full_n),
    .i_ce0(1'b0),
    .i_address0(14'd0),
    .i_q0(tdf5_fmaps_i_q0),
    .i_ce1(tdf4_111_U0_out_data_ce1),
    .i_we1(tdf4_111_U0_out_data_we1),
    .i_address1(tdf4_111_U0_out_data_address1),
    .i_d1(tdf4_111_U0_out_data_d1),
    .t_ce(1'b1),
    .t_read(tdf5_110_U0_ap_ready),
    .t_empty_n(tdf5_fmaps_t_empty_n),
    .t_ce0(tdf5_110_U0_in_data_ce0),
    .t_address0(tdf5_110_U0_in_data_address0),
    .t_q0(tdf5_fmaps_t_q0),
    .t_ce1(1'b0),
    .t_we1(1'b0),
    .t_address1(14'd0),
    .t_d1(64'd0)
);

td_fused_top_td_fused_tdf3_fmaps #(
    .DataWidth( 64 ),
    .AddressRange( 25088 ),
    .AddressWidth( 15 ))
tdf6_fmaps_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf5_110_U0_ap_done),
    .i_full_n(tdf6_fmaps_i_full_n),
    .i_ce0(1'b0),
    .i_address0(15'd0),
    .i_q0(tdf6_fmaps_i_q0),
    .i_ce1(tdf5_110_U0_out_data_ce1),
    .i_we1(tdf5_110_U0_out_data_we1),
    .i_address1(tdf5_110_U0_out_data_address1),
    .i_d1(tdf5_110_U0_out_data_d1),
    .t_ce(1'b1),
    .t_read(tdf6_19_U0_ap_ready),
    .t_empty_n(tdf6_fmaps_t_empty_n),
    .t_ce0(tdf6_19_U0_in_data_ce0),
    .t_address0(tdf6_19_U0_in_data_address0),
    .t_q0(tdf6_fmaps_t_q0),
    .t_ce1(1'b0),
    .t_we1(1'b0),
    .t_address1(15'd0),
    .t_d1(64'd0)
);

td_fused_top_td_fused_tdf7_fmaps #(
    .DataWidth( 64 ),
    .AddressRange( 6272 ),
    .AddressWidth( 13 ))
tdf7_fmaps_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf6_19_U0_ap_done),
    .i_full_n(tdf7_fmaps_i_full_n),
    .i_ce0(1'b0),
    .i_address0(13'd0),
    .i_q0(tdf7_fmaps_i_q0),
    .i_ce1(tdf6_19_U0_out_data_ce1),
    .i_we1(tdf6_19_U0_out_data_we1),
    .i_address1(tdf6_19_U0_out_data_address1),
    .i_d1(tdf6_19_U0_out_data_d1),
    .t_ce(1'b1),
    .t_read(tdf7_18_U0_ap_ready),
    .t_empty_n(tdf7_fmaps_t_empty_n),
    .t_ce0(tdf7_18_U0_in_data_ce0),
    .t_address0(tdf7_18_U0_in_data_address0),
    .t_q0(tdf7_fmaps_t_q0),
    .t_ce1(1'b0),
    .t_we1(1'b0),
    .t_address1(13'd0),
    .t_d1(64'd0)
);

td_fused_top_td_fused_tdf7_fmaps #(
    .DataWidth( 64 ),
    .AddressRange( 6272 ),
    .AddressWidth( 13 ))
tdf8_fmaps_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf7_18_U0_ap_done),
    .i_full_n(tdf8_fmaps_i_full_n),
    .i_ce0(1'b0),
    .i_address0(13'd0),
    .i_q0(tdf8_fmaps_i_q0),
    .i_ce1(tdf7_18_U0_out_data_ce1),
    .i_we1(tdf7_18_U0_out_data_we1),
    .i_address1(tdf7_18_U0_out_data_address1),
    .i_d1(tdf7_18_U0_out_data_d1),
    .t_ce(1'b1),
    .t_read(tdf8_17_U0_ap_ready),
    .t_empty_n(tdf8_fmaps_t_empty_n),
    .t_ce0(tdf8_17_U0_in_data_ce0),
    .t_address0(tdf8_17_U0_in_data_address0),
    .t_q0(tdf8_fmaps_t_q0),
    .t_ce1(1'b0),
    .t_we1(1'b0),
    .t_address1(13'd0),
    .t_d1(64'd0)
);

td_fused_top_td_fused_tdf4_fmaps #(
    .DataWidth( 64 ),
    .AddressRange( 12544 ),
    .AddressWidth( 14 ))
tdf9_fmaps_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf8_17_U0_ap_done),
    .i_full_n(tdf9_fmaps_i_full_n),
    .i_ce0(1'b0),
    .i_address0(14'd0),
    .i_q0(tdf9_fmaps_i_q0),
    .i_ce1(tdf8_17_U0_out_data_ce1),
    .i_we1(tdf8_17_U0_out_data_we1),
    .i_address1(tdf8_17_U0_out_data_address1),
    .i_d1(tdf8_17_U0_out_data_d1),
    .t_ce(1'b1),
    .t_read(tdf9_16_U0_ap_ready),
    .t_empty_n(tdf9_fmaps_t_empty_n),
    .t_ce0(tdf9_16_U0_in_data_ce0),
    .t_address0(tdf9_16_U0_in_data_address0),
    .t_q0(tdf9_fmaps_t_q0),
    .t_ce1(1'b0),
    .t_we1(1'b0),
    .t_address1(14'd0),
    .t_d1(64'd0)
);

td_fused_top_td_fused_tdf10_fmaps #(
    .DataWidth( 64 ),
    .AddressRange( 3136 ),
    .AddressWidth( 12 ))
tdf10_fmaps_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf9_16_U0_ap_done),
    .i_full_n(tdf10_fmaps_i_full_n),
    .i_ce0(1'b0),
    .i_address0(12'd0),
    .i_q0(tdf10_fmaps_i_q0),
    .i_ce1(tdf9_16_U0_out_data_ce1),
    .i_we1(tdf9_16_U0_out_data_we1),
    .i_address1(tdf9_16_U0_out_data_address1),
    .i_d1(tdf9_16_U0_out_data_d1),
    .t_ce(1'b1),
    .t_read(tdf10_15_U0_ap_ready),
    .t_empty_n(tdf10_fmaps_t_empty_n),
    .t_ce0(tdf10_15_U0_in_data_ce0),
    .t_address0(tdf10_15_U0_in_data_address0),
    .t_q0(tdf10_fmaps_t_q0),
    .t_ce1(1'b0),
    .t_we1(1'b0),
    .t_address1(12'd0),
    .t_d1(64'd0)
);

td_fused_top_td_fused_tdf10_fmaps #(
    .DataWidth( 64 ),
    .AddressRange( 3136 ),
    .AddressWidth( 12 ))
tdf11_fmaps_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf10_15_U0_ap_done),
    .i_full_n(tdf11_fmaps_i_full_n),
    .i_ce0(1'b0),
    .i_address0(12'd0),
    .i_q0(tdf11_fmaps_i_q0),
    .i_ce1(tdf10_15_U0_out_data_ce1),
    .i_we1(tdf10_15_U0_out_data_we1),
    .i_address1(tdf10_15_U0_out_data_address1),
    .i_d1(tdf10_15_U0_out_data_d1),
    .t_ce(1'b1),
    .t_read(tdf11_14_U0_ap_ready),
    .t_empty_n(tdf11_fmaps_t_empty_n),
    .t_ce0(tdf11_14_U0_in_data_ce0),
    .t_address0(tdf11_14_U0_in_data_address0),
    .t_q0(tdf11_fmaps_t_q0),
    .t_ce1(1'b0),
    .t_we1(1'b0),
    .t_address1(12'd0),
    .t_d1(64'd0)
);

td_fused_top_td_fused_tdf7_fmaps #(
    .DataWidth( 64 ),
    .AddressRange( 6272 ),
    .AddressWidth( 13 ))
tdf12_fmaps_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf11_14_U0_ap_done),
    .i_full_n(tdf12_fmaps_i_full_n),
    .i_ce0(1'b0),
    .i_address0(13'd0),
    .i_q0(tdf12_fmaps_i_q0),
    .i_ce1(tdf11_14_U0_out_data_ce1),
    .i_we1(tdf11_14_U0_out_data_we1),
    .i_address1(tdf11_14_U0_out_data_address1),
    .i_d1(tdf11_14_U0_out_data_d1),
    .t_ce(1'b1),
    .t_read(tdf12_13_U0_ap_ready),
    .t_empty_n(tdf12_fmaps_t_empty_n),
    .t_ce0(tdf12_13_U0_in_data_ce0),
    .t_address0(tdf12_13_U0_in_data_address0),
    .t_q0(tdf12_fmaps_t_q0),
    .t_ce1(1'b0),
    .t_we1(1'b0),
    .t_address1(13'd0),
    .t_d1(64'd0)
);

td_fused_top_td_fused_final_fmaps #(
    .DataWidth( 64 ),
    .AddressRange( 49000 ),
    .AddressWidth( 16 ))
final_fmaps_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .i_ce(1'b1),
    .i_write(tdf12_13_U0_ap_done),
    .i_full_n(final_fmaps_i_full_n),
    .i_ce0(1'b0),
    .i_address0(16'd0),
    .i_q0(final_fmaps_i_q0),
    .i_ce1(tdf12_13_U0_out_data_ce1),
    .i_we1(tdf12_13_U0_out_data_we1),
    .i_address1(tdf12_13_U0_out_data_address1),
    .i_d1(tdf12_13_U0_out_data_d1),
    .t_ce(1'b1),
    .t_read(td_fused_axi_out_U0_ap_ready),
    .t_empty_n(final_fmaps_t_empty_n),
    .t_ce0(td_fused_axi_out_U0_fmaps_ce0),
    .t_address0(td_fused_axi_out_U0_fmaps_address0),
    .t_q0(final_fmaps_t_q0),
    .t_ce1(1'b0),
    .t_we1(1'b0),
    .t_address1(16'd0),
    .t_d1(64'd0)
);

td_fused_top_td_fused_axi_in td_fused_axi_in_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(td_fused_axi_in_U0_ap_start),
    .ap_done(td_fused_axi_in_U0_ap_done),
    .ap_continue(td_fused_axi_in_U0_ap_continue),
    .ap_idle(td_fused_axi_in_U0_ap_idle),
    .ap_ready(td_fused_axi_in_U0_ap_ready),
    .stream_in_TDATA(stream_in_TDATA),
    .stream_in_TVALID(stream_in_TVALID),
    .stream_in_TREADY(td_fused_axi_in_U0_stream_in_TREADY),
    .stream_in_TKEEP(stream_in_TKEEP),
    .stream_in_TSTRB(stream_in_TSTRB),
    .stream_in_TLAST(stream_in_TLAST),
    .fmaps_address1(td_fused_axi_in_U0_fmaps_address1),
    .fmaps_ce1(td_fused_axi_in_U0_fmaps_ce1),
    .fmaps_we1(td_fused_axi_in_U0_fmaps_we1),
    .fmaps_d1(td_fused_axi_in_U0_fmaps_d1)
);

td_fused_top_tdf1_114 tdf1_114_U0(
    .in_data_address0(tdf1_114_U0_in_data_address0),
    .in_data_ce0(tdf1_114_U0_in_data_ce0),
    .in_data_d0(tdf1_114_U0_in_data_d0),
    .in_data_q0(tdf1_fmaps_t_q0),
    .in_data_we0(tdf1_114_U0_in_data_we0),
    .in_data_address1(tdf1_114_U0_in_data_address1),
    .in_data_ce1(tdf1_114_U0_in_data_ce1),
    .in_data_d1(tdf1_114_U0_in_data_d1),
    .in_data_q1(64'd0),
    .in_data_we1(tdf1_114_U0_in_data_we1),
    .out_data_address0(tdf1_114_U0_out_data_address0),
    .out_data_ce0(tdf1_114_U0_out_data_ce0),
    .out_data_d0(tdf1_114_U0_out_data_d0),
    .out_data_q0(64'd0),
    .out_data_we0(tdf1_114_U0_out_data_we0),
    .out_data_address1(tdf1_114_U0_out_data_address1),
    .out_data_ce1(tdf1_114_U0_out_data_ce1),
    .out_data_d1(tdf1_114_U0_out_data_d1),
    .out_data_q1(64'd0),
    .out_data_we1(tdf1_114_U0_out_data_we1),
    .filter_data_address0(tdf1_114_U0_filter_data_address0),
    .filter_data_ce0(tdf1_114_U0_filter_data_ce0),
    .filter_data_d0(tdf1_114_U0_filter_data_d0),
    .filter_data_q0(tdf1_filters_q0),
    .filter_data_we0(tdf1_114_U0_filter_data_we0),
    .filter_data_address1(tdf1_114_U0_filter_data_address1),
    .filter_data_ce1(tdf1_114_U0_filter_data_ce1),
    .filter_data_d1(tdf1_114_U0_filter_data_d1),
    .filter_data_q1(16'd0),
    .filter_data_we1(tdf1_114_U0_filter_data_we1),
    .adjustments_address0(tdf1_114_U0_adjustments_address0),
    .adjustments_ce0(tdf1_114_U0_adjustments_ce0),
    .adjustments_d0(tdf1_114_U0_adjustments_d0),
    .adjustments_q0(tdf1_adjustments_q0),
    .adjustments_we0(tdf1_114_U0_adjustments_we0),
    .adjustments_address1(tdf1_114_U0_adjustments_address1),
    .adjustments_ce1(tdf1_114_U0_adjustments_ce1),
    .adjustments_d1(tdf1_114_U0_adjustments_d1),
    .adjustments_q1(48'd0),
    .adjustments_we1(tdf1_114_U0_adjustments_we1),
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .in_data_empty_n(1'b0),
    .in_data_read(tdf1_114_U0_in_data_read),
    .out_data_full_n(tdf2_fmaps_i_full_n),
    .out_data_write(tdf1_114_U0_out_data_write),
    .ap_start(tdf1_114_U0_ap_start),
    .ap_done(tdf1_114_U0_ap_done),
    .ap_ready(tdf1_114_U0_ap_ready),
    .ap_idle(tdf1_114_U0_ap_idle),
    .ap_continue(tdf1_114_U0_ap_continue)
);

td_fused_top_tdf2_113 tdf2_113_U0(
    .in_data_address0(tdf2_113_U0_in_data_address0),
    .in_data_ce0(tdf2_113_U0_in_data_ce0),
    .in_data_d0(tdf2_113_U0_in_data_d0),
    .in_data_q0(tdf2_fmaps_t_q0),
    .in_data_we0(tdf2_113_U0_in_data_we0),
    .in_data_address1(tdf2_113_U0_in_data_address1),
    .in_data_ce1(tdf2_113_U0_in_data_ce1),
    .in_data_d1(tdf2_113_U0_in_data_d1),
    .in_data_q1(64'd0),
    .in_data_we1(tdf2_113_U0_in_data_we1),
    .out_data_address0(tdf2_113_U0_out_data_address0),
    .out_data_ce0(tdf2_113_U0_out_data_ce0),
    .out_data_d0(tdf2_113_U0_out_data_d0),
    .out_data_q0(64'd0),
    .out_data_we0(tdf2_113_U0_out_data_we0),
    .out_data_address1(tdf2_113_U0_out_data_address1),
    .out_data_ce1(tdf2_113_U0_out_data_ce1),
    .out_data_d1(tdf2_113_U0_out_data_d1),
    .out_data_q1(64'd0),
    .out_data_we1(tdf2_113_U0_out_data_we1),
    .filter_data_address0(tdf2_113_U0_filter_data_address0),
    .filter_data_ce0(tdf2_113_U0_filter_data_ce0),
    .filter_data_d0(tdf2_113_U0_filter_data_d0),
    .filter_data_q0(tdf2_filters_q0),
    .filter_data_we0(tdf2_113_U0_filter_data_we0),
    .filter_data_address1(tdf2_113_U0_filter_data_address1),
    .filter_data_ce1(tdf2_113_U0_filter_data_ce1),
    .filter_data_d1(tdf2_113_U0_filter_data_d1),
    .filter_data_q1(16'd0),
    .filter_data_we1(tdf2_113_U0_filter_data_we1),
    .adjustments_address0(tdf2_113_U0_adjustments_address0),
    .adjustments_ce0(tdf2_113_U0_adjustments_ce0),
    .adjustments_d0(tdf2_113_U0_adjustments_d0),
    .adjustments_q0(tdf2_adjustments_q0),
    .adjustments_we0(tdf2_113_U0_adjustments_we0),
    .adjustments_address1(tdf2_113_U0_adjustments_address1),
    .adjustments_ce1(tdf2_113_U0_adjustments_ce1),
    .adjustments_d1(tdf2_113_U0_adjustments_d1),
    .adjustments_q1(48'd0),
    .adjustments_we1(tdf2_113_U0_adjustments_we1),
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .in_data_empty_n(1'b0),
    .in_data_read(tdf2_113_U0_in_data_read),
    .out_data_full_n(tdf3_fmaps_i_full_n),
    .out_data_write(tdf2_113_U0_out_data_write),
    .ap_start(tdf2_113_U0_ap_start),
    .ap_done(tdf2_113_U0_ap_done),
    .ap_ready(tdf2_113_U0_ap_ready),
    .ap_idle(tdf2_113_U0_ap_idle),
    .ap_continue(tdf2_113_U0_ap_continue)
);

td_fused_top_tdf3_112 tdf3_112_U0(
    .in_data_address0(tdf3_112_U0_in_data_address0),
    .in_data_ce0(tdf3_112_U0_in_data_ce0),
    .in_data_d0(tdf3_112_U0_in_data_d0),
    .in_data_q0(tdf3_fmaps_t_q0),
    .in_data_we0(tdf3_112_U0_in_data_we0),
    .in_data_address1(tdf3_112_U0_in_data_address1),
    .in_data_ce1(tdf3_112_U0_in_data_ce1),
    .in_data_d1(tdf3_112_U0_in_data_d1),
    .in_data_q1(64'd0),
    .in_data_we1(tdf3_112_U0_in_data_we1),
    .out_data_address0(tdf3_112_U0_out_data_address0),
    .out_data_ce0(tdf3_112_U0_out_data_ce0),
    .out_data_d0(tdf3_112_U0_out_data_d0),
    .out_data_q0(64'd0),
    .out_data_we0(tdf3_112_U0_out_data_we0),
    .out_data_address1(tdf3_112_U0_out_data_address1),
    .out_data_ce1(tdf3_112_U0_out_data_ce1),
    .out_data_d1(tdf3_112_U0_out_data_d1),
    .out_data_q1(64'd0),
    .out_data_we1(tdf3_112_U0_out_data_we1),
    .filter_data_address0(tdf3_112_U0_filter_data_address0),
    .filter_data_ce0(tdf3_112_U0_filter_data_ce0),
    .filter_data_d0(tdf3_112_U0_filter_data_d0),
    .filter_data_q0(tdf3_filters_q0),
    .filter_data_we0(tdf3_112_U0_filter_data_we0),
    .filter_data_address1(tdf3_112_U0_filter_data_address1),
    .filter_data_ce1(tdf3_112_U0_filter_data_ce1),
    .filter_data_d1(tdf3_112_U0_filter_data_d1),
    .filter_data_q1(16'd0),
    .filter_data_we1(tdf3_112_U0_filter_data_we1),
    .adjustments_address0(tdf3_112_U0_adjustments_address0),
    .adjustments_ce0(tdf3_112_U0_adjustments_ce0),
    .adjustments_d0(tdf3_112_U0_adjustments_d0),
    .adjustments_q0(tdf3_adjustments_q0),
    .adjustments_we0(tdf3_112_U0_adjustments_we0),
    .adjustments_address1(tdf3_112_U0_adjustments_address1),
    .adjustments_ce1(tdf3_112_U0_adjustments_ce1),
    .adjustments_d1(tdf3_112_U0_adjustments_d1),
    .adjustments_q1(48'd0),
    .adjustments_we1(tdf3_112_U0_adjustments_we1),
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .in_data_empty_n(1'b0),
    .in_data_read(tdf3_112_U0_in_data_read),
    .out_data_full_n(tdf4_fmaps_i_full_n),
    .out_data_write(tdf3_112_U0_out_data_write),
    .ap_start(tdf3_112_U0_ap_start),
    .ap_done(tdf3_112_U0_ap_done),
    .ap_ready(tdf3_112_U0_ap_ready),
    .ap_idle(tdf3_112_U0_ap_idle),
    .ap_continue(tdf3_112_U0_ap_continue)
);

td_fused_top_tdf4_111 tdf4_111_U0(
    .in_data_address0(tdf4_111_U0_in_data_address0),
    .in_data_ce0(tdf4_111_U0_in_data_ce0),
    .in_data_d0(tdf4_111_U0_in_data_d0),
    .in_data_q0(tdf4_fmaps_t_q0),
    .in_data_we0(tdf4_111_U0_in_data_we0),
    .in_data_address1(tdf4_111_U0_in_data_address1),
    .in_data_ce1(tdf4_111_U0_in_data_ce1),
    .in_data_d1(tdf4_111_U0_in_data_d1),
    .in_data_q1(64'd0),
    .in_data_we1(tdf4_111_U0_in_data_we1),
    .out_data_address0(tdf4_111_U0_out_data_address0),
    .out_data_ce0(tdf4_111_U0_out_data_ce0),
    .out_data_d0(tdf4_111_U0_out_data_d0),
    .out_data_q0(64'd0),
    .out_data_we0(tdf4_111_U0_out_data_we0),
    .out_data_address1(tdf4_111_U0_out_data_address1),
    .out_data_ce1(tdf4_111_U0_out_data_ce1),
    .out_data_d1(tdf4_111_U0_out_data_d1),
    .out_data_q1(64'd0),
    .out_data_we1(tdf4_111_U0_out_data_we1),
    .l1_filter_data_address0(tdf4_111_U0_l1_filter_data_address0),
    .l1_filter_data_ce0(tdf4_111_U0_l1_filter_data_ce0),
    .l1_filter_data_d0(tdf4_111_U0_l1_filter_data_d0),
    .l1_filter_data_q0(tdf4_filters_q0),
    .l1_filter_data_we0(tdf4_111_U0_l1_filter_data_we0),
    .l1_filter_data_address1(tdf4_111_U0_l1_filter_data_address1),
    .l1_filter_data_ce1(tdf4_111_U0_l1_filter_data_ce1),
    .l1_filter_data_d1(tdf4_111_U0_l1_filter_data_d1),
    .l1_filter_data_q1(16'd0),
    .l1_filter_data_we1(tdf4_111_U0_l1_filter_data_we1),
    .l2_filter_data_address0(tdf4_111_U0_l2_filter_data_address0),
    .l2_filter_data_ce0(tdf4_111_U0_l2_filter_data_ce0),
    .l2_filter_data_d0(tdf4_111_U0_l2_filter_data_d0),
    .l2_filter_data_q0(tdf4_l2_filters_q0),
    .l2_filter_data_we0(tdf4_111_U0_l2_filter_data_we0),
    .l2_filter_data_address1(tdf4_111_U0_l2_filter_data_address1),
    .l2_filter_data_ce1(tdf4_111_U0_l2_filter_data_ce1),
    .l2_filter_data_d1(tdf4_111_U0_l2_filter_data_d1),
    .l2_filter_data_q1(16'd0),
    .l2_filter_data_we1(tdf4_111_U0_l2_filter_data_we1),
    .l1_adjustments_address0(tdf4_111_U0_l1_adjustments_address0),
    .l1_adjustments_ce0(tdf4_111_U0_l1_adjustments_ce0),
    .l1_adjustments_d0(tdf4_111_U0_l1_adjustments_d0),
    .l1_adjustments_q0(tdf4_adjustments_q0),
    .l1_adjustments_we0(tdf4_111_U0_l1_adjustments_we0),
    .l1_adjustments_address1(tdf4_111_U0_l1_adjustments_address1),
    .l1_adjustments_ce1(tdf4_111_U0_l1_adjustments_ce1),
    .l1_adjustments_d1(tdf4_111_U0_l1_adjustments_d1),
    .l1_adjustments_q1(48'd0),
    .l1_adjustments_we1(tdf4_111_U0_l1_adjustments_we1),
    .l2_adjustments_address0(tdf4_111_U0_l2_adjustments_address0),
    .l2_adjustments_ce0(tdf4_111_U0_l2_adjustments_ce0),
    .l2_adjustments_d0(tdf4_111_U0_l2_adjustments_d0),
    .l2_adjustments_q0(tdf4_l2_adjustments_q0),
    .l2_adjustments_we0(tdf4_111_U0_l2_adjustments_we0),
    .l2_adjustments_address1(tdf4_111_U0_l2_adjustments_address1),
    .l2_adjustments_ce1(tdf4_111_U0_l2_adjustments_ce1),
    .l2_adjustments_d1(tdf4_111_U0_l2_adjustments_d1),
    .l2_adjustments_q1(48'd0),
    .l2_adjustments_we1(tdf4_111_U0_l2_adjustments_we1),
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .in_data_empty_n(1'b0),
    .in_data_read(tdf4_111_U0_in_data_read),
    .out_data_full_n(tdf5_fmaps_i_full_n),
    .out_data_write(tdf4_111_U0_out_data_write),
    .ap_start(tdf4_111_U0_ap_start),
    .ap_done(tdf4_111_U0_ap_done),
    .ap_ready(tdf4_111_U0_ap_ready),
    .ap_idle(tdf4_111_U0_ap_idle),
    .ap_continue(tdf4_111_U0_ap_continue)
);

td_fused_top_tdf5_110 tdf5_110_U0(
    .in_data_address0(tdf5_110_U0_in_data_address0),
    .in_data_ce0(tdf5_110_U0_in_data_ce0),
    .in_data_d0(tdf5_110_U0_in_data_d0),
    .in_data_q0(tdf5_fmaps_t_q0),
    .in_data_we0(tdf5_110_U0_in_data_we0),
    .in_data_address1(tdf5_110_U0_in_data_address1),
    .in_data_ce1(tdf5_110_U0_in_data_ce1),
    .in_data_d1(tdf5_110_U0_in_data_d1),
    .in_data_q1(64'd0),
    .in_data_we1(tdf5_110_U0_in_data_we1),
    .out_data_address0(tdf5_110_U0_out_data_address0),
    .out_data_ce0(tdf5_110_U0_out_data_ce0),
    .out_data_d0(tdf5_110_U0_out_data_d0),
    .out_data_q0(64'd0),
    .out_data_we0(tdf5_110_U0_out_data_we0),
    .out_data_address1(tdf5_110_U0_out_data_address1),
    .out_data_ce1(tdf5_110_U0_out_data_ce1),
    .out_data_d1(tdf5_110_U0_out_data_d1),
    .out_data_q1(64'd0),
    .out_data_we1(tdf5_110_U0_out_data_we1),
    .filter_data_address0(tdf5_110_U0_filter_data_address0),
    .filter_data_ce0(tdf5_110_U0_filter_data_ce0),
    .filter_data_d0(tdf5_110_U0_filter_data_d0),
    .filter_data_q0(tdf5_filters_q0),
    .filter_data_we0(tdf5_110_U0_filter_data_we0),
    .filter_data_address1(tdf5_110_U0_filter_data_address1),
    .filter_data_ce1(tdf5_110_U0_filter_data_ce1),
    .filter_data_d1(tdf5_110_U0_filter_data_d1),
    .filter_data_q1(16'd0),
    .filter_data_we1(tdf5_110_U0_filter_data_we1),
    .adjustments_address0(tdf5_110_U0_adjustments_address0),
    .adjustments_ce0(tdf5_110_U0_adjustments_ce0),
    .adjustments_d0(tdf5_110_U0_adjustments_d0),
    .adjustments_q0(tdf5_adjustments_q0),
    .adjustments_we0(tdf5_110_U0_adjustments_we0),
    .adjustments_address1(tdf5_110_U0_adjustments_address1),
    .adjustments_ce1(tdf5_110_U0_adjustments_ce1),
    .adjustments_d1(tdf5_110_U0_adjustments_d1),
    .adjustments_q1(48'd0),
    .adjustments_we1(tdf5_110_U0_adjustments_we1),
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .in_data_empty_n(1'b0),
    .in_data_read(tdf5_110_U0_in_data_read),
    .out_data_full_n(tdf6_fmaps_i_full_n),
    .out_data_write(tdf5_110_U0_out_data_write),
    .ap_start(tdf5_110_U0_ap_start),
    .ap_done(tdf5_110_U0_ap_done),
    .ap_ready(tdf5_110_U0_ap_ready),
    .ap_idle(tdf5_110_U0_ap_idle),
    .ap_continue(tdf5_110_U0_ap_continue)
);

td_fused_top_tdf6_19 tdf6_19_U0(
    .in_data_address0(tdf6_19_U0_in_data_address0),
    .in_data_ce0(tdf6_19_U0_in_data_ce0),
    .in_data_d0(tdf6_19_U0_in_data_d0),
    .in_data_q0(tdf6_fmaps_t_q0),
    .in_data_we0(tdf6_19_U0_in_data_we0),
    .in_data_address1(tdf6_19_U0_in_data_address1),
    .in_data_ce1(tdf6_19_U0_in_data_ce1),
    .in_data_d1(tdf6_19_U0_in_data_d1),
    .in_data_q1(64'd0),
    .in_data_we1(tdf6_19_U0_in_data_we1),
    .out_data_address0(tdf6_19_U0_out_data_address0),
    .out_data_ce0(tdf6_19_U0_out_data_ce0),
    .out_data_d0(tdf6_19_U0_out_data_d0),
    .out_data_q0(64'd0),
    .out_data_we0(tdf6_19_U0_out_data_we0),
    .out_data_address1(tdf6_19_U0_out_data_address1),
    .out_data_ce1(tdf6_19_U0_out_data_ce1),
    .out_data_d1(tdf6_19_U0_out_data_d1),
    .out_data_q1(64'd0),
    .out_data_we1(tdf6_19_U0_out_data_we1),
    .filter_data_address0(tdf6_19_U0_filter_data_address0),
    .filter_data_ce0(tdf6_19_U0_filter_data_ce0),
    .filter_data_d0(tdf6_19_U0_filter_data_d0),
    .filter_data_q0(tdf6_filters_q0),
    .filter_data_we0(tdf6_19_U0_filter_data_we0),
    .filter_data_address1(tdf6_19_U0_filter_data_address1),
    .filter_data_ce1(tdf6_19_U0_filter_data_ce1),
    .filter_data_d1(tdf6_19_U0_filter_data_d1),
    .filter_data_q1(16'd0),
    .filter_data_we1(tdf6_19_U0_filter_data_we1),
    .adjustments_address0(tdf6_19_U0_adjustments_address0),
    .adjustments_ce0(tdf6_19_U0_adjustments_ce0),
    .adjustments_d0(tdf6_19_U0_adjustments_d0),
    .adjustments_q0(tdf6_adjustments_q0),
    .adjustments_we0(tdf6_19_U0_adjustments_we0),
    .adjustments_address1(tdf6_19_U0_adjustments_address1),
    .adjustments_ce1(tdf6_19_U0_adjustments_ce1),
    .adjustments_d1(tdf6_19_U0_adjustments_d1),
    .adjustments_q1(48'd0),
    .adjustments_we1(tdf6_19_U0_adjustments_we1),
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .in_data_empty_n(1'b0),
    .in_data_read(tdf6_19_U0_in_data_read),
    .out_data_full_n(tdf7_fmaps_i_full_n),
    .out_data_write(tdf6_19_U0_out_data_write),
    .ap_start(tdf6_19_U0_ap_start),
    .ap_done(tdf6_19_U0_ap_done),
    .ap_ready(tdf6_19_U0_ap_ready),
    .ap_idle(tdf6_19_U0_ap_idle),
    .ap_continue(tdf6_19_U0_ap_continue)
);

td_fused_top_tdf7_18 tdf7_18_U0(
    .in_data_address0(tdf7_18_U0_in_data_address0),
    .in_data_ce0(tdf7_18_U0_in_data_ce0),
    .in_data_d0(tdf7_18_U0_in_data_d0),
    .in_data_q0(tdf7_fmaps_t_q0),
    .in_data_we0(tdf7_18_U0_in_data_we0),
    .in_data_address1(tdf7_18_U0_in_data_address1),
    .in_data_ce1(tdf7_18_U0_in_data_ce1),
    .in_data_d1(tdf7_18_U0_in_data_d1),
    .in_data_q1(64'd0),
    .in_data_we1(tdf7_18_U0_in_data_we1),
    .out_data_address0(tdf7_18_U0_out_data_address0),
    .out_data_ce0(tdf7_18_U0_out_data_ce0),
    .out_data_d0(tdf7_18_U0_out_data_d0),
    .out_data_q0(64'd0),
    .out_data_we0(tdf7_18_U0_out_data_we0),
    .out_data_address1(tdf7_18_U0_out_data_address1),
    .out_data_ce1(tdf7_18_U0_out_data_ce1),
    .out_data_d1(tdf7_18_U0_out_data_d1),
    .out_data_q1(64'd0),
    .out_data_we1(tdf7_18_U0_out_data_we1),
    .l1_filter_data_address0(tdf7_18_U0_l1_filter_data_address0),
    .l1_filter_data_ce0(tdf7_18_U0_l1_filter_data_ce0),
    .l1_filter_data_d0(tdf7_18_U0_l1_filter_data_d0),
    .l1_filter_data_q0(tdf7_filters_q0),
    .l1_filter_data_we0(tdf7_18_U0_l1_filter_data_we0),
    .l1_filter_data_address1(tdf7_18_U0_l1_filter_data_address1),
    .l1_filter_data_ce1(tdf7_18_U0_l1_filter_data_ce1),
    .l1_filter_data_d1(tdf7_18_U0_l1_filter_data_d1),
    .l1_filter_data_q1(16'd0),
    .l1_filter_data_we1(tdf7_18_U0_l1_filter_data_we1),
    .l2_filter_data_address0(tdf7_18_U0_l2_filter_data_address0),
    .l2_filter_data_ce0(tdf7_18_U0_l2_filter_data_ce0),
    .l2_filter_data_d0(tdf7_18_U0_l2_filter_data_d0),
    .l2_filter_data_q0(tdf7_l2_filters_q0),
    .l2_filter_data_we0(tdf7_18_U0_l2_filter_data_we0),
    .l2_filter_data_address1(tdf7_18_U0_l2_filter_data_address1),
    .l2_filter_data_ce1(tdf7_18_U0_l2_filter_data_ce1),
    .l2_filter_data_d1(tdf7_18_U0_l2_filter_data_d1),
    .l2_filter_data_q1(16'd0),
    .l2_filter_data_we1(tdf7_18_U0_l2_filter_data_we1),
    .l1_adjustments_address0(tdf7_18_U0_l1_adjustments_address0),
    .l1_adjustments_ce0(tdf7_18_U0_l1_adjustments_ce0),
    .l1_adjustments_d0(tdf7_18_U0_l1_adjustments_d0),
    .l1_adjustments_q0(tdf7_adjustments_q0),
    .l1_adjustments_we0(tdf7_18_U0_l1_adjustments_we0),
    .l1_adjustments_address1(tdf7_18_U0_l1_adjustments_address1),
    .l1_adjustments_ce1(tdf7_18_U0_l1_adjustments_ce1),
    .l1_adjustments_d1(tdf7_18_U0_l1_adjustments_d1),
    .l1_adjustments_q1(48'd0),
    .l1_adjustments_we1(tdf7_18_U0_l1_adjustments_we1),
    .l2_adjustments_address0(tdf7_18_U0_l2_adjustments_address0),
    .l2_adjustments_ce0(tdf7_18_U0_l2_adjustments_ce0),
    .l2_adjustments_d0(tdf7_18_U0_l2_adjustments_d0),
    .l2_adjustments_q0(tdf7_l2_adjustments_q0),
    .l2_adjustments_we0(tdf7_18_U0_l2_adjustments_we0),
    .l2_adjustments_address1(tdf7_18_U0_l2_adjustments_address1),
    .l2_adjustments_ce1(tdf7_18_U0_l2_adjustments_ce1),
    .l2_adjustments_d1(tdf7_18_U0_l2_adjustments_d1),
    .l2_adjustments_q1(48'd0),
    .l2_adjustments_we1(tdf7_18_U0_l2_adjustments_we1),
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .in_data_empty_n(1'b0),
    .in_data_read(tdf7_18_U0_in_data_read),
    .out_data_full_n(tdf8_fmaps_i_full_n),
    .out_data_write(tdf7_18_U0_out_data_write),
    .ap_start(tdf7_18_U0_ap_start),
    .ap_done(tdf7_18_U0_ap_done),
    .ap_ready(tdf7_18_U0_ap_ready),
    .ap_idle(tdf7_18_U0_ap_idle),
    .ap_continue(tdf7_18_U0_ap_continue)
);

td_fused_top_tdf8_17 tdf8_17_U0(
    .in_data_address0(tdf8_17_U0_in_data_address0),
    .in_data_ce0(tdf8_17_U0_in_data_ce0),
    .in_data_d0(tdf8_17_U0_in_data_d0),
    .in_data_q0(tdf8_fmaps_t_q0),
    .in_data_we0(tdf8_17_U0_in_data_we0),
    .in_data_address1(tdf8_17_U0_in_data_address1),
    .in_data_ce1(tdf8_17_U0_in_data_ce1),
    .in_data_d1(tdf8_17_U0_in_data_d1),
    .in_data_q1(64'd0),
    .in_data_we1(tdf8_17_U0_in_data_we1),
    .out_data_address0(tdf8_17_U0_out_data_address0),
    .out_data_ce0(tdf8_17_U0_out_data_ce0),
    .out_data_d0(tdf8_17_U0_out_data_d0),
    .out_data_q0(64'd0),
    .out_data_we0(tdf8_17_U0_out_data_we0),
    .out_data_address1(tdf8_17_U0_out_data_address1),
    .out_data_ce1(tdf8_17_U0_out_data_ce1),
    .out_data_d1(tdf8_17_U0_out_data_d1),
    .out_data_q1(64'd0),
    .out_data_we1(tdf8_17_U0_out_data_we1),
    .filter_data_address0(tdf8_17_U0_filter_data_address0),
    .filter_data_ce0(tdf8_17_U0_filter_data_ce0),
    .filter_data_d0(tdf8_17_U0_filter_data_d0),
    .filter_data_q0(tdf8_filters_q0),
    .filter_data_we0(tdf8_17_U0_filter_data_we0),
    .filter_data_address1(tdf8_17_U0_filter_data_address1),
    .filter_data_ce1(tdf8_17_U0_filter_data_ce1),
    .filter_data_d1(tdf8_17_U0_filter_data_d1),
    .filter_data_q1(16'd0),
    .filter_data_we1(tdf8_17_U0_filter_data_we1),
    .adjustments_address0(tdf8_17_U0_adjustments_address0),
    .adjustments_ce0(tdf8_17_U0_adjustments_ce0),
    .adjustments_d0(tdf8_17_U0_adjustments_d0),
    .adjustments_q0(tdf8_adjustments_q0),
    .adjustments_we0(tdf8_17_U0_adjustments_we0),
    .adjustments_address1(tdf8_17_U0_adjustments_address1),
    .adjustments_ce1(tdf8_17_U0_adjustments_ce1),
    .adjustments_d1(tdf8_17_U0_adjustments_d1),
    .adjustments_q1(48'd0),
    .adjustments_we1(tdf8_17_U0_adjustments_we1),
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .in_data_empty_n(1'b0),
    .in_data_read(tdf8_17_U0_in_data_read),
    .out_data_full_n(tdf9_fmaps_i_full_n),
    .out_data_write(tdf8_17_U0_out_data_write),
    .ap_start(tdf8_17_U0_ap_start),
    .ap_done(tdf8_17_U0_ap_done),
    .ap_ready(tdf8_17_U0_ap_ready),
    .ap_idle(tdf8_17_U0_ap_idle),
    .ap_continue(tdf8_17_U0_ap_continue)
);

td_fused_top_tdf9_16 tdf9_16_U0(
    .in_data_address0(tdf9_16_U0_in_data_address0),
    .in_data_ce0(tdf9_16_U0_in_data_ce0),
    .in_data_d0(tdf9_16_U0_in_data_d0),
    .in_data_q0(tdf9_fmaps_t_q0),
    .in_data_we0(tdf9_16_U0_in_data_we0),
    .in_data_address1(tdf9_16_U0_in_data_address1),
    .in_data_ce1(tdf9_16_U0_in_data_ce1),
    .in_data_d1(tdf9_16_U0_in_data_d1),
    .in_data_q1(64'd0),
    .in_data_we1(tdf9_16_U0_in_data_we1),
    .out_data_address0(tdf9_16_U0_out_data_address0),
    .out_data_ce0(tdf9_16_U0_out_data_ce0),
    .out_data_d0(tdf9_16_U0_out_data_d0),
    .out_data_q0(64'd0),
    .out_data_we0(tdf9_16_U0_out_data_we0),
    .out_data_address1(tdf9_16_U0_out_data_address1),
    .out_data_ce1(tdf9_16_U0_out_data_ce1),
    .out_data_d1(tdf9_16_U0_out_data_d1),
    .out_data_q1(64'd0),
    .out_data_we1(tdf9_16_U0_out_data_we1),
    .filter_data_address0(tdf9_16_U0_filter_data_address0),
    .filter_data_ce0(tdf9_16_U0_filter_data_ce0),
    .filter_data_d0(tdf9_16_U0_filter_data_d0),
    .filter_data_q0(tdf9_filters_q0),
    .filter_data_we0(tdf9_16_U0_filter_data_we0),
    .filter_data_address1(tdf9_16_U0_filter_data_address1),
    .filter_data_ce1(tdf9_16_U0_filter_data_ce1),
    .filter_data_d1(tdf9_16_U0_filter_data_d1),
    .filter_data_q1(16'd0),
    .filter_data_we1(tdf9_16_U0_filter_data_we1),
    .adjustments_address0(tdf9_16_U0_adjustments_address0),
    .adjustments_ce0(tdf9_16_U0_adjustments_ce0),
    .adjustments_d0(tdf9_16_U0_adjustments_d0),
    .adjustments_q0(tdf9_adjustments_q0),
    .adjustments_we0(tdf9_16_U0_adjustments_we0),
    .adjustments_address1(tdf9_16_U0_adjustments_address1),
    .adjustments_ce1(tdf9_16_U0_adjustments_ce1),
    .adjustments_d1(tdf9_16_U0_adjustments_d1),
    .adjustments_q1(48'd0),
    .adjustments_we1(tdf9_16_U0_adjustments_we1),
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .in_data_empty_n(1'b0),
    .in_data_read(tdf9_16_U0_in_data_read),
    .out_data_full_n(tdf10_fmaps_i_full_n),
    .out_data_write(tdf9_16_U0_out_data_write),
    .ap_start(tdf9_16_U0_ap_start),
    .ap_done(tdf9_16_U0_ap_done),
    .ap_ready(tdf9_16_U0_ap_ready),
    .ap_idle(tdf9_16_U0_ap_idle),
    .ap_continue(tdf9_16_U0_ap_continue)
);

td_fused_top_tdf10_15 tdf10_15_U0(
    .in_data_address0(tdf10_15_U0_in_data_address0),
    .in_data_ce0(tdf10_15_U0_in_data_ce0),
    .in_data_d0(tdf10_15_U0_in_data_d0),
    .in_data_q0(tdf10_fmaps_t_q0),
    .in_data_we0(tdf10_15_U0_in_data_we0),
    .in_data_address1(tdf10_15_U0_in_data_address1),
    .in_data_ce1(tdf10_15_U0_in_data_ce1),
    .in_data_d1(tdf10_15_U0_in_data_d1),
    .in_data_q1(64'd0),
    .in_data_we1(tdf10_15_U0_in_data_we1),
    .out_data_address0(tdf10_15_U0_out_data_address0),
    .out_data_ce0(tdf10_15_U0_out_data_ce0),
    .out_data_d0(tdf10_15_U0_out_data_d0),
    .out_data_q0(64'd0),
    .out_data_we0(tdf10_15_U0_out_data_we0),
    .out_data_address1(tdf10_15_U0_out_data_address1),
    .out_data_ce1(tdf10_15_U0_out_data_ce1),
    .out_data_d1(tdf10_15_U0_out_data_d1),
    .out_data_q1(64'd0),
    .out_data_we1(tdf10_15_U0_out_data_we1),
    .l1_filter_data_address0(tdf10_15_U0_l1_filter_data_address0),
    .l1_filter_data_ce0(tdf10_15_U0_l1_filter_data_ce0),
    .l1_filter_data_d0(tdf10_15_U0_l1_filter_data_d0),
    .l1_filter_data_q0(tdf10_filters_q0),
    .l1_filter_data_we0(tdf10_15_U0_l1_filter_data_we0),
    .l1_filter_data_address1(tdf10_15_U0_l1_filter_data_address1),
    .l1_filter_data_ce1(tdf10_15_U0_l1_filter_data_ce1),
    .l1_filter_data_d1(tdf10_15_U0_l1_filter_data_d1),
    .l1_filter_data_q1(64'd0),
    .l1_filter_data_we1(tdf10_15_U0_l1_filter_data_we1),
    .l2_filter_data_address0(tdf10_15_U0_l2_filter_data_address0),
    .l2_filter_data_ce0(tdf10_15_U0_l2_filter_data_ce0),
    .l2_filter_data_d0(tdf10_15_U0_l2_filter_data_d0),
    .l2_filter_data_q0(tdf10_l2_filters_q0),
    .l2_filter_data_we0(tdf10_15_U0_l2_filter_data_we0),
    .l2_filter_data_address1(tdf10_15_U0_l2_filter_data_address1),
    .l2_filter_data_ce1(tdf10_15_U0_l2_filter_data_ce1),
    .l2_filter_data_d1(tdf10_15_U0_l2_filter_data_d1),
    .l2_filter_data_q1(16'd0),
    .l2_filter_data_we1(tdf10_15_U0_l2_filter_data_we1),
    .l1_adjustments_address0(tdf10_15_U0_l1_adjustments_address0),
    .l1_adjustments_ce0(tdf10_15_U0_l1_adjustments_ce0),
    .l1_adjustments_d0(tdf10_15_U0_l1_adjustments_d0),
    .l1_adjustments_q0(tdf10_adjustments_q0),
    .l1_adjustments_we0(tdf10_15_U0_l1_adjustments_we0),
    .l1_adjustments_address1(tdf10_15_U0_l1_adjustments_address1),
    .l1_adjustments_ce1(tdf10_15_U0_l1_adjustments_ce1),
    .l1_adjustments_d1(tdf10_15_U0_l1_adjustments_d1),
    .l1_adjustments_q1(48'd0),
    .l1_adjustments_we1(tdf10_15_U0_l1_adjustments_we1),
    .l2_adjustments_address0(tdf10_15_U0_l2_adjustments_address0),
    .l2_adjustments_ce0(tdf10_15_U0_l2_adjustments_ce0),
    .l2_adjustments_d0(tdf10_15_U0_l2_adjustments_d0),
    .l2_adjustments_q0(tdf10_l2_adjustments_q0),
    .l2_adjustments_we0(tdf10_15_U0_l2_adjustments_we0),
    .l2_adjustments_address1(tdf10_15_U0_l2_adjustments_address1),
    .l2_adjustments_ce1(tdf10_15_U0_l2_adjustments_ce1),
    .l2_adjustments_d1(tdf10_15_U0_l2_adjustments_d1),
    .l2_adjustments_q1(48'd0),
    .l2_adjustments_we1(tdf10_15_U0_l2_adjustments_we1),
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .in_data_empty_n(1'b0),
    .in_data_read(tdf10_15_U0_in_data_read),
    .out_data_full_n(tdf11_fmaps_i_full_n),
    .out_data_write(tdf10_15_U0_out_data_write),
    .ap_start(tdf10_15_U0_ap_start),
    .ap_done(tdf10_15_U0_ap_done),
    .ap_ready(tdf10_15_U0_ap_ready),
    .ap_idle(tdf10_15_U0_ap_idle),
    .ap_continue(tdf10_15_U0_ap_continue)
);

td_fused_top_tdf11_14 tdf11_14_U0(
    .in_data_address0(tdf11_14_U0_in_data_address0),
    .in_data_ce0(tdf11_14_U0_in_data_ce0),
    .in_data_d0(tdf11_14_U0_in_data_d0),
    .in_data_q0(tdf11_fmaps_t_q0),
    .in_data_we0(tdf11_14_U0_in_data_we0),
    .in_data_address1(tdf11_14_U0_in_data_address1),
    .in_data_ce1(tdf11_14_U0_in_data_ce1),
    .in_data_d1(tdf11_14_U0_in_data_d1),
    .in_data_q1(64'd0),
    .in_data_we1(tdf11_14_U0_in_data_we1),
    .out_data_address0(tdf11_14_U0_out_data_address0),
    .out_data_ce0(tdf11_14_U0_out_data_ce0),
    .out_data_d0(tdf11_14_U0_out_data_d0),
    .out_data_q0(64'd0),
    .out_data_we0(tdf11_14_U0_out_data_we0),
    .out_data_address1(tdf11_14_U0_out_data_address1),
    .out_data_ce1(tdf11_14_U0_out_data_ce1),
    .out_data_d1(tdf11_14_U0_out_data_d1),
    .out_data_q1(64'd0),
    .out_data_we1(tdf11_14_U0_out_data_we1),
    .l1_filter_data_address0(tdf11_14_U0_l1_filter_data_address0),
    .l1_filter_data_ce0(tdf11_14_U0_l1_filter_data_ce0),
    .l1_filter_data_d0(tdf11_14_U0_l1_filter_data_d0),
    .l1_filter_data_q0(tdf11_filters_q0),
    .l1_filter_data_we0(tdf11_14_U0_l1_filter_data_we0),
    .l1_filter_data_address1(tdf11_14_U0_l1_filter_data_address1),
    .l1_filter_data_ce1(tdf11_14_U0_l1_filter_data_ce1),
    .l1_filter_data_d1(tdf11_14_U0_l1_filter_data_d1),
    .l1_filter_data_q1(64'd0),
    .l1_filter_data_we1(tdf11_14_U0_l1_filter_data_we1),
    .l2_filter_data_address0(tdf11_14_U0_l2_filter_data_address0),
    .l2_filter_data_ce0(tdf11_14_U0_l2_filter_data_ce0),
    .l2_filter_data_d0(tdf11_14_U0_l2_filter_data_d0),
    .l2_filter_data_q0(tdf11_l2_filters_q0),
    .l2_filter_data_we0(tdf11_14_U0_l2_filter_data_we0),
    .l2_filter_data_address1(tdf11_14_U0_l2_filter_data_address1),
    .l2_filter_data_ce1(tdf11_14_U0_l2_filter_data_ce1),
    .l2_filter_data_d1(tdf11_14_U0_l2_filter_data_d1),
    .l2_filter_data_q1(16'd0),
    .l2_filter_data_we1(tdf11_14_U0_l2_filter_data_we1),
    .l1_adjustments_address0(tdf11_14_U0_l1_adjustments_address0),
    .l1_adjustments_ce0(tdf11_14_U0_l1_adjustments_ce0),
    .l1_adjustments_d0(tdf11_14_U0_l1_adjustments_d0),
    .l1_adjustments_q0(tdf11_adjustments_q0),
    .l1_adjustments_we0(tdf11_14_U0_l1_adjustments_we0),
    .l1_adjustments_address1(tdf11_14_U0_l1_adjustments_address1),
    .l1_adjustments_ce1(tdf11_14_U0_l1_adjustments_ce1),
    .l1_adjustments_d1(tdf11_14_U0_l1_adjustments_d1),
    .l1_adjustments_q1(48'd0),
    .l1_adjustments_we1(tdf11_14_U0_l1_adjustments_we1),
    .l2_adjustments_address0(tdf11_14_U0_l2_adjustments_address0),
    .l2_adjustments_ce0(tdf11_14_U0_l2_adjustments_ce0),
    .l2_adjustments_d0(tdf11_14_U0_l2_adjustments_d0),
    .l2_adjustments_q0(tdf11_l2_adjustments_q0),
    .l2_adjustments_we0(tdf11_14_U0_l2_adjustments_we0),
    .l2_adjustments_address1(tdf11_14_U0_l2_adjustments_address1),
    .l2_adjustments_ce1(tdf11_14_U0_l2_adjustments_ce1),
    .l2_adjustments_d1(tdf11_14_U0_l2_adjustments_d1),
    .l2_adjustments_q1(48'd0),
    .l2_adjustments_we1(tdf11_14_U0_l2_adjustments_we1),
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .in_data_empty_n(1'b0),
    .in_data_read(tdf11_14_U0_in_data_read),
    .out_data_full_n(tdf12_fmaps_i_full_n),
    .out_data_write(tdf11_14_U0_out_data_write),
    .ap_start(tdf11_14_U0_ap_start),
    .ap_done(tdf11_14_U0_ap_done),
    .ap_ready(tdf11_14_U0_ap_ready),
    .ap_idle(tdf11_14_U0_ap_idle),
    .ap_continue(tdf11_14_U0_ap_continue)
);

td_fused_top_tdf12_13 tdf12_13_U0(
    .in_data_address0(tdf12_13_U0_in_data_address0),
    .in_data_ce0(tdf12_13_U0_in_data_ce0),
    .in_data_d0(tdf12_13_U0_in_data_d0),
    .in_data_q0(tdf12_fmaps_t_q0),
    .in_data_we0(tdf12_13_U0_in_data_we0),
    .in_data_address1(tdf12_13_U0_in_data_address1),
    .in_data_ce1(tdf12_13_U0_in_data_ce1),
    .in_data_d1(tdf12_13_U0_in_data_d1),
    .in_data_q1(64'd0),
    .in_data_we1(tdf12_13_U0_in_data_we1),
    .out_data_address0(tdf12_13_U0_out_data_address0),
    .out_data_ce0(tdf12_13_U0_out_data_ce0),
    .out_data_d0(tdf12_13_U0_out_data_d0),
    .out_data_q0(64'd0),
    .out_data_we0(tdf12_13_U0_out_data_we0),
    .out_data_address1(tdf12_13_U0_out_data_address1),
    .out_data_ce1(tdf12_13_U0_out_data_ce1),
    .out_data_d1(tdf12_13_U0_out_data_d1),
    .out_data_q1(64'd0),
    .out_data_we1(tdf12_13_U0_out_data_we1),
    .filter_data_address0(tdf12_13_U0_filter_data_address0),
    .filter_data_ce0(tdf12_13_U0_filter_data_ce0),
    .filter_data_d0(tdf12_13_U0_filter_data_d0),
    .filter_data_q0(tdf12_filters_q0),
    .filter_data_we0(tdf12_13_U0_filter_data_we0),
    .filter_data_address1(tdf12_13_U0_filter_data_address1),
    .filter_data_ce1(tdf12_13_U0_filter_data_ce1),
    .filter_data_d1(tdf12_13_U0_filter_data_d1),
    .filter_data_q1(16'd0),
    .filter_data_we1(tdf12_13_U0_filter_data_we1),
    .adjustments_address0(tdf12_13_U0_adjustments_address0),
    .adjustments_ce0(tdf12_13_U0_adjustments_ce0),
    .adjustments_d0(tdf12_13_U0_adjustments_d0),
    .adjustments_q0(tdf12_adjustments_q0),
    .adjustments_we0(tdf12_13_U0_adjustments_we0),
    .adjustments_address1(tdf12_13_U0_adjustments_address1),
    .adjustments_ce1(tdf12_13_U0_adjustments_ce1),
    .adjustments_d1(tdf12_13_U0_adjustments_d1),
    .adjustments_q1(48'd0),
    .adjustments_we1(tdf12_13_U0_adjustments_we1),
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .in_data_empty_n(1'b0),
    .in_data_read(tdf12_13_U0_in_data_read),
    .out_data_full_n(final_fmaps_i_full_n),
    .out_data_write(tdf12_13_U0_out_data_write),
    .ap_start(tdf12_13_U0_ap_start),
    .ap_done(tdf12_13_U0_ap_done),
    .ap_ready(tdf12_13_U0_ap_ready),
    .ap_idle(tdf12_13_U0_ap_idle),
    .ap_continue(tdf12_13_U0_ap_continue)
);

td_fused_top_td_fused_axi_out td_fused_axi_out_U0(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(td_fused_axi_out_U0_ap_start),
    .ap_done(td_fused_axi_out_U0_ap_done),
    .ap_continue(td_fused_axi_out_U0_ap_continue),
    .ap_idle(td_fused_axi_out_U0_ap_idle),
    .ap_ready(td_fused_axi_out_U0_ap_ready),
    .fmaps_address0(td_fused_axi_out_U0_fmaps_address0),
    .fmaps_ce0(td_fused_axi_out_U0_fmaps_ce0),
    .fmaps_q0(final_fmaps_t_q0),
    .stream_out_TDATA(td_fused_axi_out_U0_stream_out_TDATA),
    .stream_out_TVALID(td_fused_axi_out_U0_stream_out_TVALID),
    .stream_out_TREADY(stream_out_TREADY),
    .stream_out_TKEEP(td_fused_axi_out_U0_stream_out_TKEEP),
    .stream_out_TSTRB(td_fused_axi_out_U0_stream_out_TSTRB),
    .stream_out_TLAST(td_fused_axi_out_U0_stream_out_TLAST)
);

assign ap_channel_done_final_fmaps = tdf12_13_U0_ap_done;

assign ap_channel_done_tdf10_fmaps = tdf9_16_U0_ap_done;

assign ap_channel_done_tdf11_fmaps = tdf10_15_U0_ap_done;

assign ap_channel_done_tdf12_fmaps = tdf11_14_U0_ap_done;

assign ap_channel_done_tdf1_fmaps = td_fused_axi_in_U0_ap_done;

assign ap_channel_done_tdf2_fmaps = tdf1_114_U0_ap_done;

assign ap_channel_done_tdf3_fmaps = tdf2_113_U0_ap_done;

assign ap_channel_done_tdf4_fmaps = tdf3_112_U0_ap_done;

assign ap_channel_done_tdf5_fmaps = tdf4_111_U0_ap_done;

assign ap_channel_done_tdf6_fmaps = tdf5_110_U0_ap_done;

assign ap_channel_done_tdf7_fmaps = tdf6_19_U0_ap_done;

assign ap_channel_done_tdf8_fmaps = tdf7_18_U0_ap_done;

assign ap_channel_done_tdf9_fmaps = tdf8_17_U0_ap_done;

assign ap_done = td_fused_axi_out_U0_ap_done;

assign ap_idle = (tdf9_16_U0_ap_idle & tdf8_17_U0_ap_idle & tdf7_18_U0_ap_idle & tdf6_19_U0_ap_idle & tdf5_110_U0_ap_idle & tdf4_111_U0_ap_idle & tdf3_112_U0_ap_idle & tdf2_113_U0_ap_idle & tdf1_114_U0_ap_idle & tdf12_13_U0_ap_idle & tdf11_14_U0_ap_idle & tdf10_15_U0_ap_idle & td_fused_axi_out_U0_ap_idle & td_fused_axi_in_U0_ap_idle & (final_fmaps_t_empty_n ^ 1'b1) & (tdf12_fmaps_t_empty_n ^ 1'b1) & (tdf11_fmaps_t_empty_n ^ 1'b1) & (tdf10_fmaps_t_empty_n ^ 1'b1) & (tdf9_fmaps_t_empty_n ^ 1'b1) & (tdf8_fmaps_t_empty_n ^ 1'b1) & (tdf7_fmaps_t_empty_n ^ 1'b1) & (tdf6_fmaps_t_empty_n ^ 1'b1) & (tdf5_fmaps_t_empty_n ^ 1'b1) & (tdf4_fmaps_t_empty_n ^ 1'b1) & (tdf3_fmaps_t_empty_n ^ 1'b1) & (tdf2_fmaps_t_empty_n ^ 1'b1) & (tdf1_fmaps_t_empty_n ^ 1'b1));

assign ap_ready = td_fused_axi_in_U0_ap_ready;

assign ap_sync_continue = ap_continue;

assign ap_sync_done = td_fused_axi_out_U0_ap_done;

assign ap_sync_ready = td_fused_axi_in_U0_ap_ready;

assign final_fmaps_t_d0 = 64'd0;

assign final_fmaps_t_we0 = 1'b0;

assign stream_in_TREADY = td_fused_axi_in_U0_stream_in_TREADY;

assign stream_out_TDATA = td_fused_axi_out_U0_stream_out_TDATA;

assign stream_out_TKEEP = td_fused_axi_out_U0_stream_out_TKEEP;

assign stream_out_TLAST = td_fused_axi_out_U0_stream_out_TLAST;

assign stream_out_TSTRB = td_fused_axi_out_U0_stream_out_TSTRB;

assign stream_out_TVALID = td_fused_axi_out_U0_stream_out_TVALID;

assign td_fused_axi_in_U0_ap_continue = tdf1_fmaps_i_full_n;

assign td_fused_axi_in_U0_ap_start = ap_start;

assign td_fused_axi_in_U0_fmaps_full_n = tdf1_fmaps_i_full_n;

assign td_fused_axi_in_U0_start_full_n = 1'b1;

assign td_fused_axi_in_U0_start_write = 1'b0;

assign td_fused_axi_out_U0_ap_continue = ap_continue;

assign td_fused_axi_out_U0_ap_start = final_fmaps_t_empty_n;

assign td_fused_axi_out_U0_start_full_n = 1'b1;

assign td_fused_axi_out_U0_start_write = 1'b0;

assign tdf10_15_U0_ap_continue = tdf10_15_U0_out_data_full_n;

assign tdf10_15_U0_ap_start = tdf10_fmaps_t_empty_n;

assign tdf10_15_U0_out_data_full_n = tdf11_fmaps_i_full_n;

assign tdf10_15_U0_start_full_n = 1'b1;

assign tdf10_15_U0_start_write = 1'b0;

assign tdf10_adjustments_address0 = tdf10_15_U0_l1_adjustments_address0;

assign tdf10_adjustments_address1 = 9'd0;

assign tdf10_adjustments_ce0 = tdf10_15_U0_l1_adjustments_ce0;

assign tdf10_adjustments_ce1 = 1'b0;

assign tdf10_adjustments_d0 = 48'd0;

assign tdf10_adjustments_d1 = 48'd0;

assign tdf10_adjustments_we0 = 1'b0;

assign tdf10_adjustments_we1 = 1'b0;

assign tdf10_filters_address0 = tdf10_15_U0_l1_filter_data_address0;

assign tdf10_filters_address1 = 17'd0;

assign tdf10_filters_ce0 = tdf10_15_U0_l1_filter_data_ce0;

assign tdf10_filters_ce1 = 1'b0;

assign tdf10_filters_d0 = 64'd0;

assign tdf10_filters_d1 = 64'd0;

assign tdf10_filters_we0 = 1'b0;

assign tdf10_filters_we1 = 1'b0;

assign tdf10_fmaps_t_d0 = 64'd0;

assign tdf10_fmaps_t_we0 = 1'b0;

assign tdf10_l2_adjustments_address0 = tdf10_15_U0_l2_adjustments_address0;

assign tdf10_l2_adjustments_address1 = 6'd0;

assign tdf10_l2_adjustments_ce0 = tdf10_15_U0_l2_adjustments_ce0;

assign tdf10_l2_adjustments_ce1 = 1'b0;

assign tdf10_l2_adjustments_d0 = 48'd0;

assign tdf10_l2_adjustments_d1 = 48'd0;

assign tdf10_l2_adjustments_we0 = 1'b0;

assign tdf10_l2_adjustments_we1 = 1'b0;

assign tdf10_l2_filters_address0 = tdf10_15_U0_l2_filter_data_address0;

assign tdf10_l2_filters_address1 = 15'd0;

assign tdf10_l2_filters_ce0 = tdf10_15_U0_l2_filter_data_ce0;

assign tdf10_l2_filters_ce1 = 1'b0;

assign tdf10_l2_filters_d0 = 16'd0;

assign tdf10_l2_filters_d1 = 16'd0;

assign tdf10_l2_filters_we0 = 1'b0;

assign tdf10_l2_filters_we1 = 1'b0;

assign tdf11_14_U0_ap_continue = tdf11_14_U0_out_data_full_n;

assign tdf11_14_U0_ap_start = tdf11_fmaps_t_empty_n;

assign tdf11_14_U0_out_data_full_n = tdf12_fmaps_i_full_n;

assign tdf11_14_U0_start_full_n = 1'b1;

assign tdf11_14_U0_start_write = 1'b0;

assign tdf11_adjustments_address0 = tdf11_14_U0_l1_adjustments_address0;

assign tdf11_adjustments_address1 = 9'd0;

assign tdf11_adjustments_ce0 = tdf11_14_U0_l1_adjustments_ce0;

assign tdf11_adjustments_ce1 = 1'b0;

assign tdf11_adjustments_d0 = 48'd0;

assign tdf11_adjustments_d1 = 48'd0;

assign tdf11_adjustments_we0 = 1'b0;

assign tdf11_adjustments_we1 = 1'b0;

assign tdf11_filters_address0 = tdf11_14_U0_l1_filter_data_address0;

assign tdf11_filters_address1 = 17'd0;

assign tdf11_filters_ce0 = tdf11_14_U0_l1_filter_data_ce0;

assign tdf11_filters_ce1 = 1'b0;

assign tdf11_filters_d0 = 64'd0;

assign tdf11_filters_d1 = 64'd0;

assign tdf11_filters_we0 = 1'b0;

assign tdf11_filters_we1 = 1'b0;

assign tdf11_fmaps_t_d0 = 64'd0;

assign tdf11_fmaps_t_we0 = 1'b0;

assign tdf11_l2_adjustments_address0 = tdf11_14_U0_l2_adjustments_address0;

assign tdf11_l2_adjustments_address1 = 7'd0;

assign tdf11_l2_adjustments_ce0 = tdf11_14_U0_l2_adjustments_ce0;

assign tdf11_l2_adjustments_ce1 = 1'b0;

assign tdf11_l2_adjustments_d0 = 48'd0;

assign tdf11_l2_adjustments_d1 = 48'd0;

assign tdf11_l2_adjustments_we0 = 1'b0;

assign tdf11_l2_adjustments_we1 = 1'b0;

assign tdf11_l2_filters_address0 = tdf11_14_U0_l2_filter_data_address0;

assign tdf11_l2_filters_address1 = 16'd0;

assign tdf11_l2_filters_ce0 = tdf11_14_U0_l2_filter_data_ce0;

assign tdf11_l2_filters_ce1 = 1'b0;

assign tdf11_l2_filters_d0 = 16'd0;

assign tdf11_l2_filters_d1 = 16'd0;

assign tdf11_l2_filters_we0 = 1'b0;

assign tdf11_l2_filters_we1 = 1'b0;

assign tdf12_13_U0_ap_continue = tdf12_13_U0_out_data_full_n;

assign tdf12_13_U0_ap_start = tdf12_fmaps_t_empty_n;

assign tdf12_13_U0_out_data_full_n = final_fmaps_i_full_n;

assign tdf12_13_U0_start_full_n = 1'b1;

assign tdf12_13_U0_start_write = 1'b0;

assign tdf12_adjustments_address0 = tdf12_13_U0_adjustments_address0;

assign tdf12_adjustments_address1 = 10'd0;

assign tdf12_adjustments_ce0 = tdf12_13_U0_adjustments_ce0;

assign tdf12_adjustments_ce1 = 1'b0;

assign tdf12_adjustments_d0 = 48'd0;

assign tdf12_adjustments_d1 = 48'd0;

assign tdf12_adjustments_we0 = 1'b0;

assign tdf12_adjustments_we1 = 1'b0;

assign tdf12_filters_address0 = tdf12_13_U0_filter_data_address0;

assign tdf12_filters_address1 = 17'd0;

assign tdf12_filters_ce0 = tdf12_13_U0_filter_data_ce0;

assign tdf12_filters_ce1 = 1'b0;

assign tdf12_filters_d0 = 16'd0;

assign tdf12_filters_d1 = 16'd0;

assign tdf12_filters_we0 = 1'b0;

assign tdf12_filters_we1 = 1'b0;

assign tdf12_fmaps_t_d0 = 64'd0;

assign tdf12_fmaps_t_we0 = 1'b0;

assign tdf1_114_U0_ap_continue = tdf1_114_U0_out_data_full_n;

assign tdf1_114_U0_ap_start = tdf1_fmaps_t_empty_n;

assign tdf1_114_U0_out_data_full_n = tdf2_fmaps_i_full_n;

assign tdf1_114_U0_start_full_n = 1'b1;

assign tdf1_114_U0_start_write = 1'b0;

assign tdf1_adjustments_address0 = tdf1_114_U0_adjustments_address0;

assign tdf1_adjustments_address1 = 4'd0;

assign tdf1_adjustments_ce0 = tdf1_114_U0_adjustments_ce0;

assign tdf1_adjustments_ce1 = 1'b0;

assign tdf1_adjustments_d0 = 48'd0;

assign tdf1_adjustments_d1 = 48'd0;

assign tdf1_adjustments_we0 = 1'b0;

assign tdf1_adjustments_we1 = 1'b0;

assign tdf1_filters_address0 = tdf1_114_U0_filter_data_address0;

assign tdf1_filters_address1 = 9'd0;

assign tdf1_filters_ce0 = tdf1_114_U0_filter_data_ce0;

assign tdf1_filters_ce1 = 1'b0;

assign tdf1_filters_d0 = 16'd0;

assign tdf1_filters_d1 = 16'd0;

assign tdf1_filters_we0 = 1'b0;

assign tdf1_filters_we1 = 1'b0;

assign tdf1_fmaps_t_d0 = 64'd0;

assign tdf1_fmaps_t_we0 = 1'b0;

assign tdf2_113_U0_ap_continue = tdf2_113_U0_out_data_full_n;

assign tdf2_113_U0_ap_start = tdf2_fmaps_t_empty_n;

assign tdf2_113_U0_out_data_full_n = tdf3_fmaps_i_full_n;

assign tdf2_113_U0_start_full_n = 1'b1;

assign tdf2_113_U0_start_write = 1'b0;

assign tdf2_adjustments_address0 = tdf2_113_U0_adjustments_address0;

assign tdf2_adjustments_address1 = 5'd0;

assign tdf2_adjustments_ce0 = tdf2_113_U0_adjustments_ce0;

assign tdf2_adjustments_ce1 = 1'b0;

assign tdf2_adjustments_d0 = 48'd0;

assign tdf2_adjustments_d1 = 48'd0;

assign tdf2_adjustments_we0 = 1'b0;

assign tdf2_adjustments_we1 = 1'b0;

assign tdf2_filters_address0 = tdf2_113_U0_filter_data_address0;

assign tdf2_filters_address1 = 13'd0;

assign tdf2_filters_ce0 = tdf2_113_U0_filter_data_ce0;

assign tdf2_filters_ce1 = 1'b0;

assign tdf2_filters_d0 = 16'd0;

assign tdf2_filters_d1 = 16'd0;

assign tdf2_filters_we0 = 1'b0;

assign tdf2_filters_we1 = 1'b0;

assign tdf2_fmaps_t_d0 = 64'd0;

assign tdf2_fmaps_t_we0 = 1'b0;

assign tdf3_112_U0_ap_continue = tdf3_112_U0_out_data_full_n;

assign tdf3_112_U0_ap_start = tdf3_fmaps_t_empty_n;

assign tdf3_112_U0_out_data_full_n = tdf4_fmaps_i_full_n;

assign tdf3_112_U0_start_full_n = 1'b1;

assign tdf3_112_U0_start_write = 1'b0;

assign tdf3_adjustments_address0 = tdf3_112_U0_adjustments_address0;

assign tdf3_adjustments_address1 = 4'd0;

assign tdf3_adjustments_ce0 = tdf3_112_U0_adjustments_ce0;

assign tdf3_adjustments_ce1 = 1'b0;

assign tdf3_adjustments_d0 = 48'd0;

assign tdf3_adjustments_d1 = 48'd0;

assign tdf3_adjustments_we0 = 1'b0;

assign tdf3_adjustments_we1 = 1'b0;

assign tdf3_filters_address0 = tdf3_112_U0_filter_data_address0;

assign tdf3_filters_address1 = 9'd0;

assign tdf3_filters_ce0 = tdf3_112_U0_filter_data_ce0;

assign tdf3_filters_ce1 = 1'b0;

assign tdf3_filters_d0 = 16'd0;

assign tdf3_filters_d1 = 16'd0;

assign tdf3_filters_we0 = 1'b0;

assign tdf3_filters_we1 = 1'b0;

assign tdf3_fmaps_t_d0 = 64'd0;

assign tdf3_fmaps_t_we0 = 1'b0;

assign tdf4_111_U0_ap_continue = tdf4_111_U0_out_data_full_n;

assign tdf4_111_U0_ap_start = tdf4_fmaps_t_empty_n;

assign tdf4_111_U0_out_data_full_n = tdf5_fmaps_i_full_n;

assign tdf4_111_U0_start_full_n = 1'b1;

assign tdf4_111_U0_start_write = 1'b0;

assign tdf4_adjustments_address0 = tdf4_111_U0_l1_adjustments_address0;

assign tdf4_adjustments_address1 = 7'd0;

assign tdf4_adjustments_ce0 = tdf4_111_U0_l1_adjustments_ce0;

assign tdf4_adjustments_ce1 = 1'b0;

assign tdf4_adjustments_d0 = 48'd0;

assign tdf4_adjustments_d1 = 48'd0;

assign tdf4_adjustments_we0 = 1'b0;

assign tdf4_adjustments_we1 = 1'b0;

assign tdf4_filters_address0 = tdf4_111_U0_l1_filter_data_address0;

assign tdf4_filters_address1 = 15'd0;

assign tdf4_filters_ce0 = tdf4_111_U0_l1_filter_data_ce0;

assign tdf4_filters_ce1 = 1'b0;

assign tdf4_filters_d0 = 16'd0;

assign tdf4_filters_d1 = 16'd0;

assign tdf4_filters_we0 = 1'b0;

assign tdf4_filters_we1 = 1'b0;

assign tdf4_fmaps_t_d0 = 64'd0;

assign tdf4_fmaps_t_we0 = 1'b0;

assign tdf4_l2_adjustments_address0 = tdf4_111_U0_l2_adjustments_address0;

assign tdf4_l2_adjustments_address1 = 4'd0;

assign tdf4_l2_adjustments_ce0 = tdf4_111_U0_l2_adjustments_ce0;

assign tdf4_l2_adjustments_ce1 = 1'b0;

assign tdf4_l2_adjustments_d0 = 48'd0;

assign tdf4_l2_adjustments_d1 = 48'd0;

assign tdf4_l2_adjustments_we0 = 1'b0;

assign tdf4_l2_adjustments_we1 = 1'b0;

assign tdf4_l2_filters_address0 = tdf4_111_U0_l2_filter_data_address0;

assign tdf4_l2_filters_address1 = 11'd0;

assign tdf4_l2_filters_ce0 = tdf4_111_U0_l2_filter_data_ce0;

assign tdf4_l2_filters_ce1 = 1'b0;

assign tdf4_l2_filters_d0 = 16'd0;

assign tdf4_l2_filters_d1 = 16'd0;

assign tdf4_l2_filters_we0 = 1'b0;

assign tdf4_l2_filters_we1 = 1'b0;

assign tdf5_110_U0_ap_continue = tdf5_110_U0_out_data_full_n;

assign tdf5_110_U0_ap_start = tdf5_fmaps_t_empty_n;

assign tdf5_110_U0_out_data_full_n = tdf6_fmaps_i_full_n;

assign tdf5_110_U0_start_full_n = 1'b1;

assign tdf5_110_U0_start_write = 1'b0;

assign tdf5_adjustments_address0 = tdf5_110_U0_adjustments_address0;

assign tdf5_adjustments_address1 = 7'd0;

assign tdf5_adjustments_ce0 = tdf5_110_U0_adjustments_ce0;

assign tdf5_adjustments_ce1 = 1'b0;

assign tdf5_adjustments_d0 = 48'd0;

assign tdf5_adjustments_d1 = 48'd0;

assign tdf5_adjustments_we0 = 1'b0;

assign tdf5_adjustments_we1 = 1'b0;

assign tdf5_filters_address0 = tdf5_110_U0_filter_data_address0;

assign tdf5_filters_address1 = 15'd0;

assign tdf5_filters_ce0 = tdf5_110_U0_filter_data_ce0;

assign tdf5_filters_ce1 = 1'b0;

assign tdf5_filters_d0 = 16'd0;

assign tdf5_filters_d1 = 16'd0;

assign tdf5_filters_we0 = 1'b0;

assign tdf5_filters_we1 = 1'b0;

assign tdf5_fmaps_t_d0 = 64'd0;

assign tdf5_fmaps_t_we0 = 1'b0;

assign tdf6_19_U0_ap_continue = tdf6_19_U0_out_data_full_n;

assign tdf6_19_U0_ap_start = tdf6_fmaps_t_empty_n;

assign tdf6_19_U0_out_data_full_n = tdf7_fmaps_i_full_n;

assign tdf6_19_U0_start_full_n = 1'b1;

assign tdf6_19_U0_start_write = 1'b0;

assign tdf6_adjustments_address0 = tdf6_19_U0_adjustments_address0;

assign tdf6_adjustments_address1 = 5'd0;

assign tdf6_adjustments_ce0 = tdf6_19_U0_adjustments_ce0;

assign tdf6_adjustments_ce1 = 1'b0;

assign tdf6_adjustments_d0 = 48'd0;

assign tdf6_adjustments_d1 = 48'd0;

assign tdf6_adjustments_we0 = 1'b0;

assign tdf6_adjustments_we1 = 1'b0;

assign tdf6_filters_address0 = tdf6_19_U0_filter_data_address0;

assign tdf6_filters_address1 = 12'd0;

assign tdf6_filters_ce0 = tdf6_19_U0_filter_data_ce0;

assign tdf6_filters_ce1 = 1'b0;

assign tdf6_filters_d0 = 16'd0;

assign tdf6_filters_d1 = 16'd0;

assign tdf6_filters_we0 = 1'b0;

assign tdf6_filters_we1 = 1'b0;

assign tdf6_fmaps_t_d0 = 64'd0;

assign tdf6_fmaps_t_we0 = 1'b0;

assign tdf7_18_U0_ap_continue = tdf7_18_U0_out_data_full_n;

assign tdf7_18_U0_ap_start = tdf7_fmaps_t_empty_n;

assign tdf7_18_U0_out_data_full_n = tdf8_fmaps_i_full_n;

assign tdf7_18_U0_start_full_n = 1'b1;

assign tdf7_18_U0_start_write = 1'b0;

assign tdf7_adjustments_address0 = tdf7_18_U0_l1_adjustments_address0;

assign tdf7_adjustments_address1 = 8'd0;

assign tdf7_adjustments_ce0 = tdf7_18_U0_l1_adjustments_ce0;

assign tdf7_adjustments_ce1 = 1'b0;

assign tdf7_adjustments_d0 = 48'd0;

assign tdf7_adjustments_d1 = 48'd0;

assign tdf7_adjustments_we0 = 1'b0;

assign tdf7_adjustments_we1 = 1'b0;

assign tdf7_filters_address0 = tdf7_18_U0_l1_filter_data_address0;

assign tdf7_filters_address1 = 17'd0;

assign tdf7_filters_ce0 = tdf7_18_U0_l1_filter_data_ce0;

assign tdf7_filters_ce1 = 1'b0;

assign tdf7_filters_d0 = 16'd0;

assign tdf7_filters_d1 = 16'd0;

assign tdf7_filters_we0 = 1'b0;

assign tdf7_filters_we1 = 1'b0;

assign tdf7_fmaps_t_d0 = 64'd0;

assign tdf7_fmaps_t_we0 = 1'b0;

assign tdf7_l2_adjustments_address0 = tdf7_18_U0_l2_adjustments_address0;

assign tdf7_l2_adjustments_address1 = 5'd0;

assign tdf7_l2_adjustments_ce0 = tdf7_18_U0_l2_adjustments_ce0;

assign tdf7_l2_adjustments_ce1 = 1'b0;

assign tdf7_l2_adjustments_d0 = 48'd0;

assign tdf7_l2_adjustments_d1 = 48'd0;

assign tdf7_l2_adjustments_we0 = 1'b0;

assign tdf7_l2_adjustments_we1 = 1'b0;

assign tdf7_l2_filters_address0 = tdf7_18_U0_l2_filter_data_address0;

assign tdf7_l2_filters_address1 = 13'd0;

assign tdf7_l2_filters_ce0 = tdf7_18_U0_l2_filter_data_ce0;

assign tdf7_l2_filters_ce1 = 1'b0;

assign tdf7_l2_filters_d0 = 16'd0;

assign tdf7_l2_filters_d1 = 16'd0;

assign tdf7_l2_filters_we0 = 1'b0;

assign tdf7_l2_filters_we1 = 1'b0;

assign tdf8_17_U0_ap_continue = tdf8_17_U0_out_data_full_n;

assign tdf8_17_U0_ap_start = tdf8_fmaps_t_empty_n;

assign tdf8_17_U0_out_data_full_n = tdf9_fmaps_i_full_n;

assign tdf8_17_U0_start_full_n = 1'b1;

assign tdf8_17_U0_start_write = 1'b0;

assign tdf8_adjustments_address0 = tdf8_17_U0_adjustments_address0;

assign tdf8_adjustments_address1 = 8'd0;

assign tdf8_adjustments_ce0 = tdf8_17_U0_adjustments_ce0;

assign tdf8_adjustments_ce1 = 1'b0;

assign tdf8_adjustments_d0 = 48'd0;

assign tdf8_adjustments_d1 = 48'd0;

assign tdf8_adjustments_we0 = 1'b0;

assign tdf8_adjustments_we1 = 1'b0;

assign tdf8_filters_address0 = tdf8_17_U0_filter_data_address0;

assign tdf8_filters_address1 = 17'd0;

assign tdf8_filters_ce0 = tdf8_17_U0_filter_data_ce0;

assign tdf8_filters_ce1 = 1'b0;

assign tdf8_filters_d0 = 16'd0;

assign tdf8_filters_d1 = 16'd0;

assign tdf8_filters_we0 = 1'b0;

assign tdf8_filters_we1 = 1'b0;

assign tdf8_fmaps_t_d0 = 64'd0;

assign tdf8_fmaps_t_we0 = 1'b0;

assign tdf9_16_U0_ap_continue = tdf9_16_U0_out_data_full_n;

assign tdf9_16_U0_ap_start = tdf9_fmaps_t_empty_n;

assign tdf9_16_U0_out_data_full_n = tdf10_fmaps_i_full_n;

assign tdf9_16_U0_start_full_n = 1'b1;

assign tdf9_16_U0_start_write = 1'b0;

assign tdf9_adjustments_address0 = tdf9_16_U0_adjustments_address0;

assign tdf9_adjustments_address1 = 6'd0;

assign tdf9_adjustments_ce0 = tdf9_16_U0_adjustments_ce0;

assign tdf9_adjustments_ce1 = 1'b0;

assign tdf9_adjustments_d0 = 48'd0;

assign tdf9_adjustments_d1 = 48'd0;

assign tdf9_adjustments_we0 = 1'b0;

assign tdf9_adjustments_we1 = 1'b0;

assign tdf9_filters_address0 = tdf9_16_U0_filter_data_address0;

assign tdf9_filters_address1 = 14'd0;

assign tdf9_filters_ce0 = tdf9_16_U0_filter_data_ce0;

assign tdf9_filters_ce1 = 1'b0;

assign tdf9_filters_d0 = 16'd0;

assign tdf9_filters_d1 = 16'd0;

assign tdf9_filters_we0 = 1'b0;

assign tdf9_filters_we1 = 1'b0;

assign tdf9_fmaps_t_d0 = 64'd0;

assign tdf9_fmaps_t_we0 = 1'b0;

endmodule //td_fused_top_td_fused
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2020.2 (64-bit)
// Version: 2020.2
// Copyright (C) Copyright 1986-2020 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

 

module td_fused_top (
        ap_clk,
        ap_rst_n,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        stream_in_TDATA,
        stream_in_TVALID,
        stream_in_TREADY,
        stream_in_TKEEP,
        stream_in_TSTRB,
        stream_in_TLAST,
        stream_out_TDATA,
        stream_out_TVALID,
        stream_out_TREADY,
        stream_out_TKEEP,
        stream_out_TSTRB,
        stream_out_TLAST
);

parameter    ap_ST_fsm_state1 = 5'd1;
parameter    ap_ST_fsm_state2 = 5'd2;
parameter    ap_ST_fsm_state3 = 5'd4;
parameter    ap_ST_fsm_state4 = 5'd8;
parameter    ap_ST_fsm_state5 = 5'd16;
parameter    ap_const_lv64_0 = 64'd0;

input   ap_clk;
input   ap_rst_n;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
input  [15:0] stream_in_TDATA;
input   stream_in_TVALID;
output   stream_in_TREADY;
input  [1:0] stream_in_TKEEP;
input  [1:0] stream_in_TSTRB;
input  [0:0] stream_in_TLAST;
output  [15:0] stream_out_TDATA;
output   stream_out_TVALID;
input   stream_out_TREADY;
output  [1:0] stream_out_TKEEP;
output  [1:0] stream_out_TSTRB;
output  [0:0] stream_out_TLAST;

reg ap_done;
reg ap_idle;
reg ap_ready;

 reg    ap_rst_n_inv;
  reg   [4:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
wire   [15:0] tmp_data_fu_1262_p1;
wire   [63:0] tmp_fu_1280_p5;
wire   [47:0] trunc_ln151_fu_1294_p1;
reg    tdf1_filters_ce0;
wire   [15:0] tdf1_filters_q0;
wire   [8:0] tdf1_filters_address1;
reg    tdf1_filters_ce1;
reg    tdf1_filters_we1;
reg    tdf2_filters_ce0;
wire   [15:0] tdf2_filters_q0;
wire   [12:0] tdf2_filters_address1;
reg    tdf2_filters_ce1;
reg    tdf2_filters_we1;
reg    tdf3_filters_ce0;
wire   [15:0] tdf3_filters_q0;
wire   [8:0] tdf3_filters_address1;
reg    tdf3_filters_ce1;
reg    tdf3_filters_we1;
reg    tdf4_filters_ce0;
wire   [15:0] tdf4_filters_q0;
wire   [14:0] tdf4_filters_address1;
reg    tdf4_filters_ce1;
reg    tdf4_filters_we1;
reg    tdf4_l2_filters_ce0;
wire   [15:0] tdf4_l2_filters_q0;
wire   [10:0] tdf4_l2_filters_address1;
reg    tdf4_l2_filters_ce1;
reg    tdf4_l2_filters_we1;
reg    tdf5_filters_ce0;
wire   [15:0] tdf5_filters_q0;
wire   [14:0] tdf5_filters_address1;
reg    tdf5_filters_ce1;
reg    tdf5_filters_we1;
reg    tdf6_filters_ce0;
wire   [15:0] tdf6_filters_q0;
wire   [11:0] tdf6_filters_address1;
reg    tdf6_filters_ce1;
reg    tdf6_filters_we1;
reg    tdf7_filters_ce0;
wire   [15:0] tdf7_filters_q0;
wire   [16:0] tdf7_filters_address1;
reg    tdf7_filters_ce1;
reg    tdf7_filters_we1;
reg    tdf7_l2_filters_ce0;
wire   [15:0] tdf7_l2_filters_q0;
wire   [12:0] tdf7_l2_filters_address1;
reg    tdf7_l2_filters_ce1;
reg    tdf7_l2_filters_we1;
reg    tdf8_filters_ce0;
wire   [15:0] tdf8_filters_q0;
wire   [16:0] tdf8_filters_address1;
reg    tdf8_filters_ce1;
reg    tdf8_filters_we1;
reg    tdf9_filters_ce0;
wire   [15:0] tdf9_filters_q0;
wire   [13:0] tdf9_filters_address1;
reg    tdf9_filters_ce1;
reg    tdf9_filters_we1;
reg    tdf10_filters_ce0;
wire   [63:0] tdf10_filters_q0;
wire   [16:0] tdf10_filters_address1;
reg    tdf10_filters_ce1;
reg    tdf10_filters_we1;
reg    tdf10_l2_filters_ce0;
wire   [15:0] tdf10_l2_filters_q0;
wire   [14:0] tdf10_l2_filters_address1;
reg    tdf10_l2_filters_ce1;
reg    tdf10_l2_filters_we1;
reg    tdf11_filters_ce0;
wire   [63:0] tdf11_filters_q0;
wire   [16:0] tdf11_filters_address1;
reg    tdf11_filters_ce1;
reg    tdf11_filters_we1;
reg    tdf11_l2_filters_ce0;
wire   [15:0] tdf11_l2_filters_q0;
wire   [15:0] tdf11_l2_filters_address1;
reg    tdf11_l2_filters_ce1;
reg    tdf11_l2_filters_we1;
reg    tdf12_filters_ce0;
wire   [15:0] tdf12_filters_q0;
wire   [16:0] tdf12_filters_address1;
reg    tdf12_filters_ce1;
reg    tdf12_filters_we1;
reg    tdf1_adjustments_ce0;
wire   [47:0] tdf1_adjustments_q0;
wire   [3:0] tdf1_adjustments_address1;
reg    tdf1_adjustments_ce1;
reg    tdf1_adjustments_we1;
reg    tdf2_adjustments_ce0;
wire   [47:0] tdf2_adjustments_q0;
wire   [4:0] tdf2_adjustments_address1;
reg    tdf2_adjustments_ce1;
reg    tdf2_adjustments_we1;
reg    tdf3_adjustments_ce0;
wire   [47:0] tdf3_adjustments_q0;
wire   [3:0] tdf3_adjustments_address1;
reg    tdf3_adjustments_ce1;
reg    tdf3_adjustments_we1;
reg    tdf4_adjustments_ce0;
wire   [47:0] tdf4_adjustments_q0;
wire   [6:0] tdf4_adjustments_address1;
reg    tdf4_adjustments_ce1;
reg    tdf4_adjustments_we1;
reg    tdf4_l2_adjustments_ce0;
wire   [47:0] tdf4_l2_adjustments_q0;
wire   [3:0] tdf4_l2_adjustments_address1;
reg    tdf4_l2_adjustments_ce1;
reg    tdf4_l2_adjustments_we1;
reg    tdf5_adjustments_ce0;
wire   [47:0] tdf5_adjustments_q0;
wire   [6:0] tdf5_adjustments_address1;
reg    tdf5_adjustments_ce1;
reg    tdf5_adjustments_we1;
reg    tdf6_adjustments_ce0;
wire   [47:0] tdf6_adjustments_q0;
wire   [4:0] tdf6_adjustments_address1;
reg    tdf6_adjustments_ce1;
reg    tdf6_adjustments_we1;
reg    tdf7_adjustments_ce0;
wire   [47:0] tdf7_adjustments_q0;
wire   [7:0] tdf7_adjustments_address1;
reg    tdf7_adjustments_ce1;
reg    tdf7_adjustments_we1;
reg    tdf7_l2_adjustments_ce0;
wire   [47:0] tdf7_l2_adjustments_q0;
wire   [4:0] tdf7_l2_adjustments_address1;
reg    tdf7_l2_adjustments_ce1;
reg    tdf7_l2_adjustments_we1;
reg    tdf8_adjustments_ce0;
wire   [47:0] tdf8_adjustments_q0;
wire   [7:0] tdf8_adjustments_address1;
reg    tdf8_adjustments_ce1;
reg    tdf8_adjustments_we1;
reg    tdf9_adjustments_ce0;
wire   [47:0] tdf9_adjustments_q0;
wire   [5:0] tdf9_adjustments_address1;
reg    tdf9_adjustments_ce1;
reg    tdf9_adjustments_we1;
reg    tdf10_adjustments_ce0;
wire   [47:0] tdf10_adjustments_q0;
wire   [8:0] tdf10_adjustments_address1;
reg    tdf10_adjustments_ce1;
reg    tdf10_adjustments_we1;
reg    tdf10_l2_adjustments_ce0;
wire   [47:0] tdf10_l2_adjustments_q0;
wire   [5:0] tdf10_l2_adjustments_address1;
reg    tdf10_l2_adjustments_ce1;
reg    tdf10_l2_adjustments_we1;
reg    tdf11_adjustments_ce0;
wire   [47:0] tdf11_adjustments_q0;
wire   [8:0] tdf11_adjustments_address1;
reg    tdf11_adjustments_ce1;
reg    tdf11_adjustments_we1;
reg    tdf11_l2_adjustments_ce0;
wire   [47:0] tdf11_l2_adjustments_q0;
wire   [6:0] tdf11_l2_adjustments_address1;
reg    tdf11_l2_adjustments_ce1;
reg    tdf11_l2_adjustments_we1;
reg    tdf12_adjustments_ce0;
wire   [47:0] tdf12_adjustments_q0;
wire   [9:0] tdf12_adjustments_address1;
reg    tdf12_adjustments_ce1;
reg    tdf12_adjustments_we1;
wire   [8:0] grp_td_fused_fu_990_tdf1_filters_address0;
wire    grp_td_fused_fu_990_tdf1_filters_ce0;
wire   [15:0] grp_td_fused_fu_990_tdf1_filters_d0;
wire    grp_td_fused_fu_990_tdf1_filters_we0;
wire   [8:0] grp_td_fused_fu_990_tdf1_filters_address1;
wire    grp_td_fused_fu_990_tdf1_filters_ce1;
wire   [15:0] grp_td_fused_fu_990_tdf1_filters_d1;
wire    grp_td_fused_fu_990_tdf1_filters_we1;
wire   [12:0] grp_td_fused_fu_990_tdf2_filters_address0;
wire    grp_td_fused_fu_990_tdf2_filters_ce0;
wire   [15:0] grp_td_fused_fu_990_tdf2_filters_d0;
wire    grp_td_fused_fu_990_tdf2_filters_we0;
wire   [12:0] grp_td_fused_fu_990_tdf2_filters_address1;
wire    grp_td_fused_fu_990_tdf2_filters_ce1;
wire   [15:0] grp_td_fused_fu_990_tdf2_filters_d1;
wire    grp_td_fused_fu_990_tdf2_filters_we1;
wire   [8:0] grp_td_fused_fu_990_tdf3_filters_address0;
wire    grp_td_fused_fu_990_tdf3_filters_ce0;
wire   [15:0] grp_td_fused_fu_990_tdf3_filters_d0;
wire    grp_td_fused_fu_990_tdf3_filters_we0;
wire   [8:0] grp_td_fused_fu_990_tdf3_filters_address1;
wire    grp_td_fused_fu_990_tdf3_filters_ce1;
wire   [15:0] grp_td_fused_fu_990_tdf3_filters_d1;
wire    grp_td_fused_fu_990_tdf3_filters_we1;
wire   [14:0] grp_td_fused_fu_990_tdf4_filters_address0;
wire    grp_td_fused_fu_990_tdf4_filters_ce0;
wire   [15:0] grp_td_fused_fu_990_tdf4_filters_d0;
wire    grp_td_fused_fu_990_tdf4_filters_we0;
wire   [14:0] grp_td_fused_fu_990_tdf4_filters_address1;
wire    grp_td_fused_fu_990_tdf4_filters_ce1;
wire   [15:0] grp_td_fused_fu_990_tdf4_filters_d1;
wire    grp_td_fused_fu_990_tdf4_filters_we1;
wire   [10:0] grp_td_fused_fu_990_tdf4_l2_filters_address0;
wire    grp_td_fused_fu_990_tdf4_l2_filters_ce0;
wire   [15:0] grp_td_fused_fu_990_tdf4_l2_filters_d0;
wire    grp_td_fused_fu_990_tdf4_l2_filters_we0;
wire   [10:0] grp_td_fused_fu_990_tdf4_l2_filters_address1;
wire    grp_td_fused_fu_990_tdf4_l2_filters_ce1;
wire   [15:0] grp_td_fused_fu_990_tdf4_l2_filters_d1;
wire    grp_td_fused_fu_990_tdf4_l2_filters_we1;
wire   [14:0] grp_td_fused_fu_990_tdf5_filters_address0;
wire    grp_td_fused_fu_990_tdf5_filters_ce0;
wire   [15:0] grp_td_fused_fu_990_tdf5_filters_d0;
wire    grp_td_fused_fu_990_tdf5_filters_we0;
wire   [14:0] grp_td_fused_fu_990_tdf5_filters_address1;
wire    grp_td_fused_fu_990_tdf5_filters_ce1;
wire   [15:0] grp_td_fused_fu_990_tdf5_filters_d1;
wire    grp_td_fused_fu_990_tdf5_filters_we1;
wire   [11:0] grp_td_fused_fu_990_tdf6_filters_address0;
wire    grp_td_fused_fu_990_tdf6_filters_ce0;
wire   [15:0] grp_td_fused_fu_990_tdf6_filters_d0;
wire    grp_td_fused_fu_990_tdf6_filters_we0;
wire   [11:0] grp_td_fused_fu_990_tdf6_filters_address1;
wire    grp_td_fused_fu_990_tdf6_filters_ce1;
wire   [15:0] grp_td_fused_fu_990_tdf6_filters_d1;
wire    grp_td_fused_fu_990_tdf6_filters_we1;
wire   [16:0] grp_td_fused_fu_990_tdf7_filters_address0;
wire    grp_td_fused_fu_990_tdf7_filters_ce0;
wire   [15:0] grp_td_fused_fu_990_tdf7_filters_d0;
wire    grp_td_fused_fu_990_tdf7_filters_we0;
wire   [16:0] grp_td_fused_fu_990_tdf7_filters_address1;
wire    grp_td_fused_fu_990_tdf7_filters_ce1;
wire   [15:0] grp_td_fused_fu_990_tdf7_filters_d1;
wire    grp_td_fused_fu_990_tdf7_filters_we1;
wire   [12:0] grp_td_fused_fu_990_tdf7_l2_filters_address0;
wire    grp_td_fused_fu_990_tdf7_l2_filters_ce0;
wire   [15:0] grp_td_fused_fu_990_tdf7_l2_filters_d0;
wire    grp_td_fused_fu_990_tdf7_l2_filters_we0;
wire   [12:0] grp_td_fused_fu_990_tdf7_l2_filters_address1;
wire    grp_td_fused_fu_990_tdf7_l2_filters_ce1;
wire   [15:0] grp_td_fused_fu_990_tdf7_l2_filters_d1;
wire    grp_td_fused_fu_990_tdf7_l2_filters_we1;
wire   [16:0] grp_td_fused_fu_990_tdf8_filters_address0;
wire    grp_td_fused_fu_990_tdf8_filters_ce0;
wire   [15:0] grp_td_fused_fu_990_tdf8_filters_d0;
wire    grp_td_fused_fu_990_tdf8_filters_we0;
wire   [16:0] grp_td_fused_fu_990_tdf8_filters_address1;
wire    grp_td_fused_fu_990_tdf8_filters_ce1;
wire   [15:0] grp_td_fused_fu_990_tdf8_filters_d1;
wire    grp_td_fused_fu_990_tdf8_filters_we1;
wire   [13:0] grp_td_fused_fu_990_tdf9_filters_address0;
wire    grp_td_fused_fu_990_tdf9_filters_ce0;
wire   [15:0] grp_td_fused_fu_990_tdf9_filters_d0;
wire    grp_td_fused_fu_990_tdf9_filters_we0;
wire   [13:0] grp_td_fused_fu_990_tdf9_filters_address1;
wire    grp_td_fused_fu_990_tdf9_filters_ce1;
wire   [15:0] grp_td_fused_fu_990_tdf9_filters_d1;
wire    grp_td_fused_fu_990_tdf9_filters_we1;
wire   [16:0] grp_td_fused_fu_990_tdf10_filters_address0;
wire    grp_td_fused_fu_990_tdf10_filters_ce0;
wire   [63:0] grp_td_fused_fu_990_tdf10_filters_d0;
wire    grp_td_fused_fu_990_tdf10_filters_we0;
wire   [16:0] grp_td_fused_fu_990_tdf10_filters_address1;
wire    grp_td_fused_fu_990_tdf10_filters_ce1;
wire   [63:0] grp_td_fused_fu_990_tdf10_filters_d1;
wire    grp_td_fused_fu_990_tdf10_filters_we1;
wire   [14:0] grp_td_fused_fu_990_tdf10_l2_filters_address0;
wire    grp_td_fused_fu_990_tdf10_l2_filters_ce0;
wire   [15:0] grp_td_fused_fu_990_tdf10_l2_filters_d0;
wire    grp_td_fused_fu_990_tdf10_l2_filters_we0;
wire   [14:0] grp_td_fused_fu_990_tdf10_l2_filters_address1;
wire    grp_td_fused_fu_990_tdf10_l2_filters_ce1;
wire   [15:0] grp_td_fused_fu_990_tdf10_l2_filters_d1;
wire    grp_td_fused_fu_990_tdf10_l2_filters_we1;
wire   [16:0] grp_td_fused_fu_990_tdf11_filters_address0;
wire    grp_td_fused_fu_990_tdf11_filters_ce0;
wire   [63:0] grp_td_fused_fu_990_tdf11_filters_d0;
wire    grp_td_fused_fu_990_tdf11_filters_we0;
wire   [16:0] grp_td_fused_fu_990_tdf11_filters_address1;
wire    grp_td_fused_fu_990_tdf11_filters_ce1;
wire   [63:0] grp_td_fused_fu_990_tdf11_filters_d1;
wire    grp_td_fused_fu_990_tdf11_filters_we1;
wire   [15:0] grp_td_fused_fu_990_tdf11_l2_filters_address0;
wire    grp_td_fused_fu_990_tdf11_l2_filters_ce0;
wire   [15:0] grp_td_fused_fu_990_tdf11_l2_filters_d0;
wire    grp_td_fused_fu_990_tdf11_l2_filters_we0;
wire   [15:0] grp_td_fused_fu_990_tdf11_l2_filters_address1;
wire    grp_td_fused_fu_990_tdf11_l2_filters_ce1;
wire   [15:0] grp_td_fused_fu_990_tdf11_l2_filters_d1;
wire    grp_td_fused_fu_990_tdf11_l2_filters_we1;
wire   [16:0] grp_td_fused_fu_990_tdf12_filters_address0;
wire    grp_td_fused_fu_990_tdf12_filters_ce0;
wire   [15:0] grp_td_fused_fu_990_tdf12_filters_d0;
wire    grp_td_fused_fu_990_tdf12_filters_we0;
wire   [16:0] grp_td_fused_fu_990_tdf12_filters_address1;
wire    grp_td_fused_fu_990_tdf12_filters_ce1;
wire   [15:0] grp_td_fused_fu_990_tdf12_filters_d1;
wire    grp_td_fused_fu_990_tdf12_filters_we1;
wire   [3:0] grp_td_fused_fu_990_tdf1_adjustments_address0;
wire    grp_td_fused_fu_990_tdf1_adjustments_ce0;
wire   [47:0] grp_td_fused_fu_990_tdf1_adjustments_d0;
wire    grp_td_fused_fu_990_tdf1_adjustments_we0;
wire   [3:0] grp_td_fused_fu_990_tdf1_adjustments_address1;
wire    grp_td_fused_fu_990_tdf1_adjustments_ce1;
wire   [47:0] grp_td_fused_fu_990_tdf1_adjustments_d1;
wire    grp_td_fused_fu_990_tdf1_adjustments_we1;
wire   [4:0] grp_td_fused_fu_990_tdf2_adjustments_address0;
wire    grp_td_fused_fu_990_tdf2_adjustments_ce0;
wire   [47:0] grp_td_fused_fu_990_tdf2_adjustments_d0;
wire    grp_td_fused_fu_990_tdf2_adjustments_we0;
wire   [4:0] grp_td_fused_fu_990_tdf2_adjustments_address1;
wire    grp_td_fused_fu_990_tdf2_adjustments_ce1;
wire   [47:0] grp_td_fused_fu_990_tdf2_adjustments_d1;
wire    grp_td_fused_fu_990_tdf2_adjustments_we1;
wire   [3:0] grp_td_fused_fu_990_tdf3_adjustments_address0;
wire    grp_td_fused_fu_990_tdf3_adjustments_ce0;
wire   [47:0] grp_td_fused_fu_990_tdf3_adjustments_d0;
wire    grp_td_fused_fu_990_tdf3_adjustments_we0;
wire   [3:0] grp_td_fused_fu_990_tdf3_adjustments_address1;
wire    grp_td_fused_fu_990_tdf3_adjustments_ce1;
wire   [47:0] grp_td_fused_fu_990_tdf3_adjustments_d1;
wire    grp_td_fused_fu_990_tdf3_adjustments_we1;
wire   [6:0] grp_td_fused_fu_990_tdf4_adjustments_address0;
wire    grp_td_fused_fu_990_tdf4_adjustments_ce0;
wire   [47:0] grp_td_fused_fu_990_tdf4_adjustments_d0;
wire    grp_td_fused_fu_990_tdf4_adjustments_we0;
wire   [6:0] grp_td_fused_fu_990_tdf4_adjustments_address1;
wire    grp_td_fused_fu_990_tdf4_adjustments_ce1;
wire   [47:0] grp_td_fused_fu_990_tdf4_adjustments_d1;
wire    grp_td_fused_fu_990_tdf4_adjustments_we1;
wire   [3:0] grp_td_fused_fu_990_tdf4_l2_adjustments_address0;
wire    grp_td_fused_fu_990_tdf4_l2_adjustments_ce0;
wire   [47:0] grp_td_fused_fu_990_tdf4_l2_adjustments_d0;
wire    grp_td_fused_fu_990_tdf4_l2_adjustments_we0;
wire   [3:0] grp_td_fused_fu_990_tdf4_l2_adjustments_address1;
wire    grp_td_fused_fu_990_tdf4_l2_adjustments_ce1;
wire   [47:0] grp_td_fused_fu_990_tdf4_l2_adjustments_d1;
wire    grp_td_fused_fu_990_tdf4_l2_adjustments_we1;
wire   [6:0] grp_td_fused_fu_990_tdf5_adjustments_address0;
wire    grp_td_fused_fu_990_tdf5_adjustments_ce0;
wire   [47:0] grp_td_fused_fu_990_tdf5_adjustments_d0;
wire    grp_td_fused_fu_990_tdf5_adjustments_we0;
wire   [6:0] grp_td_fused_fu_990_tdf5_adjustments_address1;
wire    grp_td_fused_fu_990_tdf5_adjustments_ce1;
wire   [47:0] grp_td_fused_fu_990_tdf5_adjustments_d1;
wire    grp_td_fused_fu_990_tdf5_adjustments_we1;
wire   [4:0] grp_td_fused_fu_990_tdf6_adjustments_address0;
wire    grp_td_fused_fu_990_tdf6_adjustments_ce0;
wire   [47:0] grp_td_fused_fu_990_tdf6_adjustments_d0;
wire    grp_td_fused_fu_990_tdf6_adjustments_we0;
wire   [4:0] grp_td_fused_fu_990_tdf6_adjustments_address1;
wire    grp_td_fused_fu_990_tdf6_adjustments_ce1;
wire   [47:0] grp_td_fused_fu_990_tdf6_adjustments_d1;
wire    grp_td_fused_fu_990_tdf6_adjustments_we1;
wire   [7:0] grp_td_fused_fu_990_tdf7_adjustments_address0;
wire    grp_td_fused_fu_990_tdf7_adjustments_ce0;
wire   [47:0] grp_td_fused_fu_990_tdf7_adjustments_d0;
wire    grp_td_fused_fu_990_tdf7_adjustments_we0;
wire   [7:0] grp_td_fused_fu_990_tdf7_adjustments_address1;
wire    grp_td_fused_fu_990_tdf7_adjustments_ce1;
wire   [47:0] grp_td_fused_fu_990_tdf7_adjustments_d1;
wire    grp_td_fused_fu_990_tdf7_adjustments_we1;
wire   [4:0] grp_td_fused_fu_990_tdf7_l2_adjustments_address0;
wire    grp_td_fused_fu_990_tdf7_l2_adjustments_ce0;
wire   [47:0] grp_td_fused_fu_990_tdf7_l2_adjustments_d0;
wire    grp_td_fused_fu_990_tdf7_l2_adjustments_we0;
wire   [4:0] grp_td_fused_fu_990_tdf7_l2_adjustments_address1;
wire    grp_td_fused_fu_990_tdf7_l2_adjustments_ce1;
wire   [47:0] grp_td_fused_fu_990_tdf7_l2_adjustments_d1;
wire    grp_td_fused_fu_990_tdf7_l2_adjustments_we1;
wire   [7:0] grp_td_fused_fu_990_tdf8_adjustments_address0;
wire    grp_td_fused_fu_990_tdf8_adjustments_ce0;
wire   [47:0] grp_td_fused_fu_990_tdf8_adjustments_d0;
wire    grp_td_fused_fu_990_tdf8_adjustments_we0;
wire   [7:0] grp_td_fused_fu_990_tdf8_adjustments_address1;
wire    grp_td_fused_fu_990_tdf8_adjustments_ce1;
wire   [47:0] grp_td_fused_fu_990_tdf8_adjustments_d1;
wire    grp_td_fused_fu_990_tdf8_adjustments_we1;
wire   [5:0] grp_td_fused_fu_990_tdf9_adjustments_address0;
wire    grp_td_fused_fu_990_tdf9_adjustments_ce0;
wire   [47:0] grp_td_fused_fu_990_tdf9_adjustments_d0;
wire    grp_td_fused_fu_990_tdf9_adjustments_we0;
wire   [5:0] grp_td_fused_fu_990_tdf9_adjustments_address1;
wire    grp_td_fused_fu_990_tdf9_adjustments_ce1;
wire   [47:0] grp_td_fused_fu_990_tdf9_adjustments_d1;
wire    grp_td_fused_fu_990_tdf9_adjustments_we1;
wire   [8:0] grp_td_fused_fu_990_tdf10_adjustments_address0;
wire    grp_td_fused_fu_990_tdf10_adjustments_ce0;
wire   [47:0] grp_td_fused_fu_990_tdf10_adjustments_d0;
wire    grp_td_fused_fu_990_tdf10_adjustments_we0;
wire   [8:0] grp_td_fused_fu_990_tdf10_adjustments_address1;
wire    grp_td_fused_fu_990_tdf10_adjustments_ce1;
wire   [47:0] grp_td_fused_fu_990_tdf10_adjustments_d1;
wire    grp_td_fused_fu_990_tdf10_adjustments_we1;
wire   [5:0] grp_td_fused_fu_990_tdf10_l2_adjustments_address0;
wire    grp_td_fused_fu_990_tdf10_l2_adjustments_ce0;
wire   [47:0] grp_td_fused_fu_990_tdf10_l2_adjustments_d0;
wire    grp_td_fused_fu_990_tdf10_l2_adjustments_we0;
wire   [5:0] grp_td_fused_fu_990_tdf10_l2_adjustments_address1;
wire    grp_td_fused_fu_990_tdf10_l2_adjustments_ce1;
wire   [47:0] grp_td_fused_fu_990_tdf10_l2_adjustments_d1;
wire    grp_td_fused_fu_990_tdf10_l2_adjustments_we1;
wire   [8:0] grp_td_fused_fu_990_tdf11_adjustments_address0;
wire    grp_td_fused_fu_990_tdf11_adjustments_ce0;
wire   [47:0] grp_td_fused_fu_990_tdf11_adjustments_d0;
wire    grp_td_fused_fu_990_tdf11_adjustments_we0;
wire   [8:0] grp_td_fused_fu_990_tdf11_adjustments_address1;
wire    grp_td_fused_fu_990_tdf11_adjustments_ce1;
wire   [47:0] grp_td_fused_fu_990_tdf11_adjustments_d1;
wire    grp_td_fused_fu_990_tdf11_adjustments_we1;
wire   [6:0] grp_td_fused_fu_990_tdf11_l2_adjustments_address0;
wire    grp_td_fused_fu_990_tdf11_l2_adjustments_ce0;
wire   [47:0] grp_td_fused_fu_990_tdf11_l2_adjustments_d0;
wire    grp_td_fused_fu_990_tdf11_l2_adjustments_we0;
wire   [6:0] grp_td_fused_fu_990_tdf11_l2_adjustments_address1;
wire    grp_td_fused_fu_990_tdf11_l2_adjustments_ce1;
wire   [47:0] grp_td_fused_fu_990_tdf11_l2_adjustments_d1;
wire    grp_td_fused_fu_990_tdf11_l2_adjustments_we1;
wire   [9:0] grp_td_fused_fu_990_tdf12_adjustments_address0;
wire    grp_td_fused_fu_990_tdf12_adjustments_ce0;
wire   [47:0] grp_td_fused_fu_990_tdf12_adjustments_d0;
wire    grp_td_fused_fu_990_tdf12_adjustments_we0;
wire   [9:0] grp_td_fused_fu_990_tdf12_adjustments_address1;
wire    grp_td_fused_fu_990_tdf12_adjustments_ce1;
wire   [47:0] grp_td_fused_fu_990_tdf12_adjustments_d1;
wire    grp_td_fused_fu_990_tdf12_adjustments_we1;
wire   [15:0] grp_td_fused_fu_990_stream_out_TDATA;
wire   [1:0] grp_td_fused_fu_990_stream_out_TKEEP;
wire   [1:0] grp_td_fused_fu_990_stream_out_TSTRB;
wire   [0:0] grp_td_fused_fu_990_stream_out_TLAST;
wire    grp_td_fused_fu_990_stream_in_TREADY;
wire    grp_td_fused_fu_990_ap_start;
wire    grp_td_fused_fu_990_stream_out_TVALID;
wire    grp_td_fused_fu_990_stream_out_TREADY;
wire    grp_td_fused_fu_990_ap_done;
wire    grp_td_fused_fu_990_ap_ready;
wire    grp_td_fused_fu_990_ap_idle;
reg    grp_td_fused_fu_990_ap_continue;
reg    grp_td_fused_fu_990_ap_start_reg;
wire    ap_CS_fsm_state3;
wire    ap_CS_fsm_state4;
wire    ap_sync_grp_td_fused_fu_990_ap_ready;
wire    ap_sync_grp_td_fused_fu_990_ap_done;
reg    ap_block_state4_on_subcall_done;
reg    ap_sync_reg_grp_td_fused_fu_990_ap_ready;
reg    ap_sync_reg_grp_td_fused_fu_990_ap_done;
wire    ap_CS_fsm_state2;
wire    ap_CS_fsm_state5;
wire    regslice_both_stream_out_V_data_V_U_apdone_blk;
reg   [4:0] ap_NS_fsm;
wire    regslice_both_stream_in_V_data_V_U_apdone_blk;
wire   [15:0] stream_in_TDATA_int_regslice;
wire    stream_in_TVALID_int_regslice;
reg    stream_in_TREADY_int_regslice;
wire    regslice_both_stream_in_V_data_V_U_ack_in;
wire    regslice_both_stream_in_V_keep_V_U_apdone_blk;
wire   [1:0] stream_in_TKEEP_int_regslice;
wire    regslice_both_stream_in_V_keep_V_U_vld_out;
wire    regslice_both_stream_in_V_keep_V_U_ack_in;
wire    regslice_both_stream_in_V_strb_V_U_apdone_blk;
wire   [1:0] stream_in_TSTRB_int_regslice;
wire    regslice_both_stream_in_V_strb_V_U_vld_out;
wire    regslice_both_stream_in_V_strb_V_U_ack_in;
wire    regslice_both_stream_in_V_last_V_U_apdone_blk;
wire   [0:0] stream_in_TLAST_int_regslice;
wire    regslice_both_stream_in_V_last_V_U_vld_out;
wire    regslice_both_stream_in_V_last_V_U_ack_in;
wire    stream_out_TREADY_int_regslice;
wire    regslice_both_stream_out_V_data_V_U_vld_out;
wire    regslice_both_stream_out_V_keep_V_U_apdone_blk;
wire    regslice_both_stream_out_V_keep_V_U_ack_in_dummy;
wire    regslice_both_stream_out_V_keep_V_U_vld_out;
wire    regslice_both_stream_out_V_strb_V_U_apdone_blk;
wire    regslice_both_stream_out_V_strb_V_U_ack_in_dummy;
wire    regslice_both_stream_out_V_strb_V_U_vld_out;
wire    regslice_both_stream_out_V_last_V_U_apdone_blk;
wire    regslice_both_stream_out_V_last_V_U_ack_in_dummy;
wire    regslice_both_stream_out_V_last_V_U_vld_out;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_CS_fsm = 5'd1;
#0 grp_td_fused_fu_990_ap_start_reg = 1'b0;
#0 ap_sync_reg_grp_td_fused_fu_990_ap_ready = 1'b0;
#0 ap_sync_reg_grp_td_fused_fu_990_ap_done = 1'b0;
end

td_fused_top_tdf1_filters #(
    .DataWidth( 16 ),
    .AddressRange( 432 ),
    .AddressWidth( 9 ))
tdf1_filters_U(
    .reset(ap_rst_n_inv),
    .clk(ap_clk),
    .address0(grp_td_fused_fu_990_tdf1_filters_address0),
    .ce0(tdf1_filters_ce0),
    .q0(tdf1_filters_q0),
    .address1(tdf1_filters_address1),
    .ce1(tdf1_filters_ce1),
    .we1(tdf1_filters_we1),
    .d1(tmp_data_fu_1262_p1)
);

td_fused_top_tdf2_filters #(
    .DataWidth( 16 ),
    .AddressRange( 4608 ),
    .AddressWidth( 13 ))
tdf2_filters_U(
    .reset(ap_rst_n_inv),
    .clk(ap_clk),
    .address0(grp_td_fused_fu_990_tdf2_filters_address0),
    .ce0(tdf2_filters_ce0),
    .q0(tdf2_filters_q0),
    .address1(tdf2_filters_address1),
    .ce1(tdf2_filters_ce1),
    .we1(tdf2_filters_we1),
    .d1(tmp_data_fu_1262_p1)
);

td_fused_top_tdf3_filters #(
    .DataWidth( 16 ),
    .AddressRange( 512 ),
    .AddressWidth( 9 ))
tdf3_filters_U(
    .reset(ap_rst_n_inv),
    .clk(ap_clk),
    .address0(grp_td_fused_fu_990_tdf3_filters_address0),
    .ce0(tdf3_filters_ce0),
    .q0(tdf3_filters_q0),
    .address1(tdf3_filters_address1),
    .ce1(tdf3_filters_ce1),
    .we1(tdf3_filters_we1),
    .d1(tmp_data_fu_1262_p1)
);

td_fused_top_tdf4_filters #(
    .DataWidth( 16 ),
    .AddressRange( 18432 ),
    .AddressWidth( 15 ))
tdf4_filters_U(
    .reset(ap_rst_n_inv),
    .clk(ap_clk),
    .address0(grp_td_fused_fu_990_tdf4_filters_address0),
    .ce0(tdf4_filters_ce0),
    .q0(tdf4_filters_q0),
    .address1(tdf4_filters_address1),
    .ce1(tdf4_filters_ce1),
    .we1(tdf4_filters_we1),
    .d1(tmp_data_fu_1262_p1)
);

td_fused_top_tdf4_l2_filters #(
    .DataWidth( 16 ),
    .AddressRange( 2048 ),
    .AddressWidth( 11 ))
tdf4_l2_filters_U(
    .reset(ap_rst_n_inv),
    .clk(ap_clk),
    .address0(grp_td_fused_fu_990_tdf4_l2_filters_address0),
    .ce0(tdf4_l2_filters_ce0),
    .q0(tdf4_l2_filters_q0),
    .address1(tdf4_l2_filters_address1),
    .ce1(tdf4_l2_filters_ce1),
    .we1(tdf4_l2_filters_we1),
    .d1(tmp_data_fu_1262_p1)
);

td_fused_top_tdf4_filters #(
    .DataWidth( 16 ),
    .AddressRange( 18432 ),
    .AddressWidth( 15 ))
tdf5_filters_U(
    .reset(ap_rst_n_inv),
    .clk(ap_clk),
    .address0(grp_td_fused_fu_990_tdf5_filters_address0),
    .ce0(tdf5_filters_ce0),
    .q0(tdf5_filters_q0),
    .address1(tdf5_filters_address1),
    .ce1(tdf5_filters_ce1),
    .we1(tdf5_filters_we1),
    .d1(tmp_data_fu_1262_p1)
);

td_fused_top_tdf6_filters #(
    .DataWidth( 16 ),
    .AddressRange( 4096 ),
    .AddressWidth( 12 ))
tdf6_filters_U(
    .reset(ap_rst_n_inv),
    .clk(ap_clk),
    .address0(grp_td_fused_fu_990_tdf6_filters_address0),
    .ce0(tdf6_filters_ce0),
    .q0(tdf6_filters_q0),
    .address1(tdf6_filters_address1),
    .ce1(tdf6_filters_ce1),
    .we1(tdf6_filters_we1),
    .d1(tmp_data_fu_1262_p1)
);

td_fused_top_tdf7_filters #(
    .DataWidth( 16 ),
    .AddressRange( 73728 ),
    .AddressWidth( 17 ))
tdf7_filters_U(
    .reset(ap_rst_n_inv),
    .clk(ap_clk),
    .address0(grp_td_fused_fu_990_tdf7_filters_address0),
    .ce0(tdf7_filters_ce0),
    .q0(tdf7_filters_q0),
    .address1(tdf7_filters_address1),
    .ce1(tdf7_filters_ce1),
    .we1(tdf7_filters_we1),
    .d1(tmp_data_fu_1262_p1)
);

td_fused_top_tdf7_l2_filters #(
    .DataWidth( 16 ),
    .AddressRange( 8192 ),
    .AddressWidth( 13 ))
tdf7_l2_filters_U(
    .reset(ap_rst_n_inv),
    .clk(ap_clk),
    .address0(grp_td_fused_fu_990_tdf7_l2_filters_address0),
    .ce0(tdf7_l2_filters_ce0),
    .q0(tdf7_l2_filters_q0),
    .address1(tdf7_l2_filters_address1),
    .ce1(tdf7_l2_filters_ce1),
    .we1(tdf7_l2_filters_we1),
    .d1(tmp_data_fu_1262_p1)
);

td_fused_top_tdf7_filters #(
    .DataWidth( 16 ),
    .AddressRange( 73728 ),
    .AddressWidth( 17 ))
tdf8_filters_U(
    .reset(ap_rst_n_inv),
    .clk(ap_clk),
    .address0(grp_td_fused_fu_990_tdf8_filters_address0),
    .ce0(tdf8_filters_ce0),
    .q0(tdf8_filters_q0),
    .address1(tdf8_filters_address1),
    .ce1(tdf8_filters_ce1),
    .we1(tdf8_filters_we1),
    .d1(tmp_data_fu_1262_p1)
);

td_fused_top_tdf9_filters #(
    .DataWidth( 16 ),
    .AddressRange( 16384 ),
    .AddressWidth( 14 ))
tdf9_filters_U(
    .reset(ap_rst_n_inv),
    .clk(ap_clk),
    .address0(grp_td_fused_fu_990_tdf9_filters_address0),
    .ce0(tdf9_filters_ce0),
    .q0(tdf9_filters_q0),
    .address1(tdf9_filters_address1),
    .ce1(tdf9_filters_ce1),
    .we1(tdf9_filters_we1),
    .d1(tmp_data_fu_1262_p1)
);

td_fused_top_tdf10_filters #(
    .DataWidth( 64 ),
    .AddressRange( 73728 ),
    .AddressWidth( 17 ))
tdf10_filters_U(
    .reset(ap_rst_n_inv),
    .clk(ap_clk),
    .address0(grp_td_fused_fu_990_tdf10_filters_address0),
    .ce0(tdf10_filters_ce0),
    .q0(tdf10_filters_q0),
    .address1(tdf10_filters_address1),
    .ce1(tdf10_filters_ce1),
    .we1(tdf10_filters_we1),
    .d1(tmp_fu_1280_p5)
);

td_fused_top_tdf10_l2_filters #(
    .DataWidth( 16 ),
    .AddressRange( 32768 ),
    .AddressWidth( 15 ))
tdf10_l2_filters_U(
    .reset(ap_rst_n_inv),
    .clk(ap_clk),
    .address0(grp_td_fused_fu_990_tdf10_l2_filters_address0),
    .ce0(tdf10_l2_filters_ce0),
    .q0(tdf10_l2_filters_q0),
    .address1(tdf10_l2_filters_address1),
    .ce1(tdf10_l2_filters_ce1),
    .we1(tdf10_l2_filters_we1),
    .d1(tmp_data_fu_1262_p1)
);

td_fused_top_tdf10_filters #(
    .DataWidth( 64 ),
    .AddressRange( 73728 ),
    .AddressWidth( 17 ))
tdf11_filters_U(
    .reset(ap_rst_n_inv),
    .clk(ap_clk),
    .address0(grp_td_fused_fu_990_tdf11_filters_address0),
    .ce0(tdf11_filters_ce0),
    .q0(tdf11_filters_q0),
    .address1(tdf11_filters_address1),
    .ce1(tdf11_filters_ce1),
    .we1(tdf11_filters_we1),
    .d1(tmp_fu_1280_p5)
);

td_fused_top_tdf11_l2_filters #(
    .DataWidth( 16 ),
    .AddressRange( 65536 ),
    .AddressWidth( 16 ))
tdf11_l2_filters_U(
    .reset(ap_rst_n_inv),
    .clk(ap_clk),
    .address0(grp_td_fused_fu_990_tdf11_l2_filters_address0),
    .ce0(tdf11_l2_filters_ce0),
    .q0(tdf11_l2_filters_q0),
    .address1(tdf11_l2_filters_address1),
    .ce1(tdf11_l2_filters_ce1),
    .we1(tdf11_l2_filters_we1),
    .d1(tmp_data_fu_1262_p1)
);

td_fused_top_tdf12_filters #(
    .DataWidth( 16 ),
    .AddressRange( 128000 ),
    .AddressWidth( 17 ))
tdf12_filters_U(
    .reset(ap_rst_n_inv),
    .clk(ap_clk),
    .address0(grp_td_fused_fu_990_tdf12_filters_address0),
    .ce0(tdf12_filters_ce0),
    .q0(tdf12_filters_q0),
    .address1(tdf12_filters_address1),
    .ce1(tdf12_filters_ce1),
    .we1(tdf12_filters_we1),
    .d1(tmp_data_fu_1262_p1)
);

td_fused_top_tdf1_adjustments #(
    .DataWidth( 48 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
tdf1_adjustments_U(
    .reset(ap_rst_n_inv),
    .clk(ap_clk),
    .address0(grp_td_fused_fu_990_tdf1_adjustments_address0),
    .ce0(tdf1_adjustments_ce0),
    .q0(tdf1_adjustments_q0),
    .address1(tdf1_adjustments_address1),
    .ce1(tdf1_adjustments_ce1),
    .we1(tdf1_adjustments_we1),
    .d1(trunc_ln151_fu_1294_p1)
);

td_fused_top_tdf2_adjustments #(
    .DataWidth( 48 ),
    .AddressRange( 32 ),
    .AddressWidth( 5 ))
tdf2_adjustments_U(
    .reset(ap_rst_n_inv),
    .clk(ap_clk),
    .address0(grp_td_fused_fu_990_tdf2_adjustments_address0),
    .ce0(tdf2_adjustments_ce0),
    .q0(tdf2_adjustments_q0),
    .address1(tdf2_adjustments_address1),
    .ce1(tdf2_adjustments_ce1),
    .we1(tdf2_adjustments_we1),
    .d1(trunc_ln151_fu_1294_p1)
);

td_fused_top_tdf1_adjustments #(
    .DataWidth( 48 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
tdf3_adjustments_U(
    .reset(ap_rst_n_inv),
    .clk(ap_clk),
    .address0(grp_td_fused_fu_990_tdf3_adjustments_address0),
    .ce0(tdf3_adjustments_ce0),
    .q0(tdf3_adjustments_q0),
    .address1(tdf3_adjustments_address1),
    .ce1(tdf3_adjustments_ce1),
    .we1(tdf3_adjustments_we1),
    .d1(trunc_ln151_fu_1294_p1)
);

td_fused_top_tdf4_adjustments #(
    .DataWidth( 48 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
tdf4_adjustments_U(
    .reset(ap_rst_n_inv),
    .clk(ap_clk),
    .address0(grp_td_fused_fu_990_tdf4_adjustments_address0),
    .ce0(tdf4_adjustments_ce0),
    .q0(tdf4_adjustments_q0),
    .address1(tdf4_adjustments_address1),
    .ce1(tdf4_adjustments_ce1),
    .we1(tdf4_adjustments_we1),
    .d1(trunc_ln151_fu_1294_p1)
);

td_fused_top_tdf1_adjustments #(
    .DataWidth( 48 ),
    .AddressRange( 16 ),
    .AddressWidth( 4 ))
tdf4_l2_adjustments_U(
    .reset(ap_rst_n_inv),
    .clk(ap_clk),
    .address0(grp_td_fused_fu_990_tdf4_l2_adjustments_address0),
    .ce0(tdf4_l2_adjustments_ce0),
    .q0(tdf4_l2_adjustments_q0),
    .address1(tdf4_l2_adjustments_address1),
    .ce1(tdf4_l2_adjustments_ce1),
    .we1(tdf4_l2_adjustments_we1),
    .d1(trunc_ln151_fu_1294_p1)
);

td_fused_top_tdf4_adjustments #(
    .DataWidth( 48 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
tdf5_adjustments_U(
    .reset(ap_rst_n_inv),
    .clk(ap_clk),
    .address0(grp_td_fused_fu_990_tdf5_adjustments_address0),
    .ce0(tdf5_adjustments_ce0),
    .q0(tdf5_adjustments_q0),
    .address1(tdf5_adjustments_address1),
    .ce1(tdf5_adjustments_ce1),
    .we1(tdf5_adjustments_we1),
    .d1(trunc_ln151_fu_1294_p1)
);

td_fused_top_tdf2_adjustments #(
    .DataWidth( 48 ),
    .AddressRange( 32 ),
    .AddressWidth( 5 ))
tdf6_adjustments_U(
    .reset(ap_rst_n_inv),
    .clk(ap_clk),
    .address0(grp_td_fused_fu_990_tdf6_adjustments_address0),
    .ce0(tdf6_adjustments_ce0),
    .q0(tdf6_adjustments_q0),
    .address1(tdf6_adjustments_address1),
    .ce1(tdf6_adjustments_ce1),
    .we1(tdf6_adjustments_we1),
    .d1(trunc_ln151_fu_1294_p1)
);

td_fused_top_tdf7_adjustments #(
    .DataWidth( 48 ),
    .AddressRange( 256 ),
    .AddressWidth( 8 ))
tdf7_adjustments_U(
    .reset(ap_rst_n_inv),
    .clk(ap_clk),
    .address0(grp_td_fused_fu_990_tdf7_adjustments_address0),
    .ce0(tdf7_adjustments_ce0),
    .q0(tdf7_adjustments_q0),
    .address1(tdf7_adjustments_address1),
    .ce1(tdf7_adjustments_ce1),
    .we1(tdf7_adjustments_we1),
    .d1(trunc_ln151_fu_1294_p1)
);

td_fused_top_tdf2_adjustments #(
    .DataWidth( 48 ),
    .AddressRange( 32 ),
    .AddressWidth( 5 ))
tdf7_l2_adjustments_U(
    .reset(ap_rst_n_inv),
    .clk(ap_clk),
    .address0(grp_td_fused_fu_990_tdf7_l2_adjustments_address0),
    .ce0(tdf7_l2_adjustments_ce0),
    .q0(tdf7_l2_adjustments_q0),
    .address1(tdf7_l2_adjustments_address1),
    .ce1(tdf7_l2_adjustments_ce1),
    .we1(tdf7_l2_adjustments_we1),
    .d1(trunc_ln151_fu_1294_p1)
);

td_fused_top_tdf7_adjustments #(
    .DataWidth( 48 ),
    .AddressRange( 256 ),
    .AddressWidth( 8 ))
tdf8_adjustments_U(
    .reset(ap_rst_n_inv),
    .clk(ap_clk),
    .address0(grp_td_fused_fu_990_tdf8_adjustments_address0),
    .ce0(tdf8_adjustments_ce0),
    .q0(tdf8_adjustments_q0),
    .address1(tdf8_adjustments_address1),
    .ce1(tdf8_adjustments_ce1),
    .we1(tdf8_adjustments_we1),
    .d1(trunc_ln151_fu_1294_p1)
);

td_fused_top_tdf9_adjustments #(
    .DataWidth( 48 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
tdf9_adjustments_U(
    .reset(ap_rst_n_inv),
    .clk(ap_clk),
    .address0(grp_td_fused_fu_990_tdf9_adjustments_address0),
    .ce0(tdf9_adjustments_ce0),
    .q0(tdf9_adjustments_q0),
    .address1(tdf9_adjustments_address1),
    .ce1(tdf9_adjustments_ce1),
    .we1(tdf9_adjustments_we1),
    .d1(trunc_ln151_fu_1294_p1)
);

td_fused_top_tdf10_adjustments #(
    .DataWidth( 48 ),
    .AddressRange( 512 ),
    .AddressWidth( 9 ))
tdf10_adjustments_U(
    .reset(ap_rst_n_inv),
    .clk(ap_clk),
    .address0(grp_td_fused_fu_990_tdf10_adjustments_address0),
    .ce0(tdf10_adjustments_ce0),
    .q0(tdf10_adjustments_q0),
    .address1(tdf10_adjustments_address1),
    .ce1(tdf10_adjustments_ce1),
    .we1(tdf10_adjustments_we1),
    .d1(trunc_ln151_fu_1294_p1)
);

td_fused_top_tdf9_adjustments #(
    .DataWidth( 48 ),
    .AddressRange( 64 ),
    .AddressWidth( 6 ))
tdf10_l2_adjustments_U(
    .reset(ap_rst_n_inv),
    .clk(ap_clk),
    .address0(grp_td_fused_fu_990_tdf10_l2_adjustments_address0),
    .ce0(tdf10_l2_adjustments_ce0),
    .q0(tdf10_l2_adjustments_q0),
    .address1(tdf10_l2_adjustments_address1),
    .ce1(tdf10_l2_adjustments_ce1),
    .we1(tdf10_l2_adjustments_we1),
    .d1(trunc_ln151_fu_1294_p1)
);

td_fused_top_tdf10_adjustments #(
    .DataWidth( 48 ),
    .AddressRange( 512 ),
    .AddressWidth( 9 ))
tdf11_adjustments_U(
    .reset(ap_rst_n_inv),
    .clk(ap_clk),
    .address0(grp_td_fused_fu_990_tdf11_adjustments_address0),
    .ce0(tdf11_adjustments_ce0),
    .q0(tdf11_adjustments_q0),
    .address1(tdf11_adjustments_address1),
    .ce1(tdf11_adjustments_ce1),
    .we1(tdf11_adjustments_we1),
    .d1(trunc_ln151_fu_1294_p1)
);

td_fused_top_tdf4_adjustments #(
    .DataWidth( 48 ),
    .AddressRange( 128 ),
    .AddressWidth( 7 ))
tdf11_l2_adjustments_U(
    .reset(ap_rst_n_inv),
    .clk(ap_clk),
    .address0(grp_td_fused_fu_990_tdf11_l2_adjustments_address0),
    .ce0(tdf11_l2_adjustments_ce0),
    .q0(tdf11_l2_adjustments_q0),
    .address1(tdf11_l2_adjustments_address1),
    .ce1(tdf11_l2_adjustments_ce1),
    .we1(tdf11_l2_adjustments_we1),
    .d1(trunc_ln151_fu_1294_p1)
);

td_fused_top_tdf12_adjustments #(
    .DataWidth( 48 ),
    .AddressRange( 1000 ),
    .AddressWidth( 10 ))
tdf12_adjustments_U(
    .reset(ap_rst_n_inv),
    .clk(ap_clk),
    .address0(grp_td_fused_fu_990_tdf12_adjustments_address0),
    .ce0(tdf12_adjustments_ce0),
    .q0(tdf12_adjustments_q0),
    .address1(tdf12_adjustments_address1),
    .ce1(tdf12_adjustments_ce1),
    .we1(tdf12_adjustments_we1),
    .d1(trunc_ln151_fu_1294_p1)
);

td_fused_top_td_fused grp_td_fused_fu_990(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .tdf1_filters_address0(grp_td_fused_fu_990_tdf1_filters_address0),
    .tdf1_filters_ce0(grp_td_fused_fu_990_tdf1_filters_ce0),
    .tdf1_filters_d0(grp_td_fused_fu_990_tdf1_filters_d0),
    .tdf1_filters_q0(tdf1_filters_q0),
    .tdf1_filters_we0(grp_td_fused_fu_990_tdf1_filters_we0),
    .tdf1_filters_address1(grp_td_fused_fu_990_tdf1_filters_address1),
    .tdf1_filters_ce1(grp_td_fused_fu_990_tdf1_filters_ce1),
    .tdf1_filters_d1(grp_td_fused_fu_990_tdf1_filters_d1),
    .tdf1_filters_q1(16'd0),
    .tdf1_filters_we1(grp_td_fused_fu_990_tdf1_filters_we1),
    .tdf2_filters_address0(grp_td_fused_fu_990_tdf2_filters_address0),
    .tdf2_filters_ce0(grp_td_fused_fu_990_tdf2_filters_ce0),
    .tdf2_filters_d0(grp_td_fused_fu_990_tdf2_filters_d0),
    .tdf2_filters_q0(tdf2_filters_q0),
    .tdf2_filters_we0(grp_td_fused_fu_990_tdf2_filters_we0),
    .tdf2_filters_address1(grp_td_fused_fu_990_tdf2_filters_address1),
    .tdf2_filters_ce1(grp_td_fused_fu_990_tdf2_filters_ce1),
    .tdf2_filters_d1(grp_td_fused_fu_990_tdf2_filters_d1),
    .tdf2_filters_q1(16'd0),
    .tdf2_filters_we1(grp_td_fused_fu_990_tdf2_filters_we1),
    .tdf3_filters_address0(grp_td_fused_fu_990_tdf3_filters_address0),
    .tdf3_filters_ce0(grp_td_fused_fu_990_tdf3_filters_ce0),
    .tdf3_filters_d0(grp_td_fused_fu_990_tdf3_filters_d0),
    .tdf3_filters_q0(tdf3_filters_q0),
    .tdf3_filters_we0(grp_td_fused_fu_990_tdf3_filters_we0),
    .tdf3_filters_address1(grp_td_fused_fu_990_tdf3_filters_address1),
    .tdf3_filters_ce1(grp_td_fused_fu_990_tdf3_filters_ce1),
    .tdf3_filters_d1(grp_td_fused_fu_990_tdf3_filters_d1),
    .tdf3_filters_q1(16'd0),
    .tdf3_filters_we1(grp_td_fused_fu_990_tdf3_filters_we1),
    .tdf4_filters_address0(grp_td_fused_fu_990_tdf4_filters_address0),
    .tdf4_filters_ce0(grp_td_fused_fu_990_tdf4_filters_ce0),
    .tdf4_filters_d0(grp_td_fused_fu_990_tdf4_filters_d0),
    .tdf4_filters_q0(tdf4_filters_q0),
    .tdf4_filters_we0(grp_td_fused_fu_990_tdf4_filters_we0),
    .tdf4_filters_address1(grp_td_fused_fu_990_tdf4_filters_address1),
    .tdf4_filters_ce1(grp_td_fused_fu_990_tdf4_filters_ce1),
    .tdf4_filters_d1(grp_td_fused_fu_990_tdf4_filters_d1),
    .tdf4_filters_q1(16'd0),
    .tdf4_filters_we1(grp_td_fused_fu_990_tdf4_filters_we1),
    .tdf4_l2_filters_address0(grp_td_fused_fu_990_tdf4_l2_filters_address0),
    .tdf4_l2_filters_ce0(grp_td_fused_fu_990_tdf4_l2_filters_ce0),
    .tdf4_l2_filters_d0(grp_td_fused_fu_990_tdf4_l2_filters_d0),
    .tdf4_l2_filters_q0(tdf4_l2_filters_q0),
    .tdf4_l2_filters_we0(grp_td_fused_fu_990_tdf4_l2_filters_we0),
    .tdf4_l2_filters_address1(grp_td_fused_fu_990_tdf4_l2_filters_address1),
    .tdf4_l2_filters_ce1(grp_td_fused_fu_990_tdf4_l2_filters_ce1),
    .tdf4_l2_filters_d1(grp_td_fused_fu_990_tdf4_l2_filters_d1),
    .tdf4_l2_filters_q1(16'd0),
    .tdf4_l2_filters_we1(grp_td_fused_fu_990_tdf4_l2_filters_we1),
    .tdf5_filters_address0(grp_td_fused_fu_990_tdf5_filters_address0),
    .tdf5_filters_ce0(grp_td_fused_fu_990_tdf5_filters_ce0),
    .tdf5_filters_d0(grp_td_fused_fu_990_tdf5_filters_d0),
    .tdf5_filters_q0(tdf5_filters_q0),
    .tdf5_filters_we0(grp_td_fused_fu_990_tdf5_filters_we0),
    .tdf5_filters_address1(grp_td_fused_fu_990_tdf5_filters_address1),
    .tdf5_filters_ce1(grp_td_fused_fu_990_tdf5_filters_ce1),
    .tdf5_filters_d1(grp_td_fused_fu_990_tdf5_filters_d1),
    .tdf5_filters_q1(16'd0),
    .tdf5_filters_we1(grp_td_fused_fu_990_tdf5_filters_we1),
    .tdf6_filters_address0(grp_td_fused_fu_990_tdf6_filters_address0),
    .tdf6_filters_ce0(grp_td_fused_fu_990_tdf6_filters_ce0),
    .tdf6_filters_d0(grp_td_fused_fu_990_tdf6_filters_d0),
    .tdf6_filters_q0(tdf6_filters_q0),
    .tdf6_filters_we0(grp_td_fused_fu_990_tdf6_filters_we0),
    .tdf6_filters_address1(grp_td_fused_fu_990_tdf6_filters_address1),
    .tdf6_filters_ce1(grp_td_fused_fu_990_tdf6_filters_ce1),
    .tdf6_filters_d1(grp_td_fused_fu_990_tdf6_filters_d1),
    .tdf6_filters_q1(16'd0),
    .tdf6_filters_we1(grp_td_fused_fu_990_tdf6_filters_we1),
    .tdf7_filters_address0(grp_td_fused_fu_990_tdf7_filters_address0),
    .tdf7_filters_ce0(grp_td_fused_fu_990_tdf7_filters_ce0),
    .tdf7_filters_d0(grp_td_fused_fu_990_tdf7_filters_d0),
    .tdf7_filters_q0(tdf7_filters_q0),
    .tdf7_filters_we0(grp_td_fused_fu_990_tdf7_filters_we0),
    .tdf7_filters_address1(grp_td_fused_fu_990_tdf7_filters_address1),
    .tdf7_filters_ce1(grp_td_fused_fu_990_tdf7_filters_ce1),
    .tdf7_filters_d1(grp_td_fused_fu_990_tdf7_filters_d1),
    .tdf7_filters_q1(16'd0),
    .tdf7_filters_we1(grp_td_fused_fu_990_tdf7_filters_we1),
    .tdf7_l2_filters_address0(grp_td_fused_fu_990_tdf7_l2_filters_address0),
    .tdf7_l2_filters_ce0(grp_td_fused_fu_990_tdf7_l2_filters_ce0),
    .tdf7_l2_filters_d0(grp_td_fused_fu_990_tdf7_l2_filters_d0),
    .tdf7_l2_filters_q0(tdf7_l2_filters_q0),
    .tdf7_l2_filters_we0(grp_td_fused_fu_990_tdf7_l2_filters_we0),
    .tdf7_l2_filters_address1(grp_td_fused_fu_990_tdf7_l2_filters_address1),
    .tdf7_l2_filters_ce1(grp_td_fused_fu_990_tdf7_l2_filters_ce1),
    .tdf7_l2_filters_d1(grp_td_fused_fu_990_tdf7_l2_filters_d1),
    .tdf7_l2_filters_q1(16'd0),
    .tdf7_l2_filters_we1(grp_td_fused_fu_990_tdf7_l2_filters_we1),
    .tdf8_filters_address0(grp_td_fused_fu_990_tdf8_filters_address0),
    .tdf8_filters_ce0(grp_td_fused_fu_990_tdf8_filters_ce0),
    .tdf8_filters_d0(grp_td_fused_fu_990_tdf8_filters_d0),
    .tdf8_filters_q0(tdf8_filters_q0),
    .tdf8_filters_we0(grp_td_fused_fu_990_tdf8_filters_we0),
    .tdf8_filters_address1(grp_td_fused_fu_990_tdf8_filters_address1),
    .tdf8_filters_ce1(grp_td_fused_fu_990_tdf8_filters_ce1),
    .tdf8_filters_d1(grp_td_fused_fu_990_tdf8_filters_d1),
    .tdf8_filters_q1(16'd0),
    .tdf8_filters_we1(grp_td_fused_fu_990_tdf8_filters_we1),
    .tdf9_filters_address0(grp_td_fused_fu_990_tdf9_filters_address0),
    .tdf9_filters_ce0(grp_td_fused_fu_990_tdf9_filters_ce0),
    .tdf9_filters_d0(grp_td_fused_fu_990_tdf9_filters_d0),
    .tdf9_filters_q0(tdf9_filters_q0),
    .tdf9_filters_we0(grp_td_fused_fu_990_tdf9_filters_we0),
    .tdf9_filters_address1(grp_td_fused_fu_990_tdf9_filters_address1),
    .tdf9_filters_ce1(grp_td_fused_fu_990_tdf9_filters_ce1),
    .tdf9_filters_d1(grp_td_fused_fu_990_tdf9_filters_d1),
    .tdf9_filters_q1(16'd0),
    .tdf9_filters_we1(grp_td_fused_fu_990_tdf9_filters_we1),
    .tdf10_filters_address0(grp_td_fused_fu_990_tdf10_filters_address0),
    .tdf10_filters_ce0(grp_td_fused_fu_990_tdf10_filters_ce0),
    .tdf10_filters_d0(grp_td_fused_fu_990_tdf10_filters_d0),
    .tdf10_filters_q0(tdf10_filters_q0),
    .tdf10_filters_we0(grp_td_fused_fu_990_tdf10_filters_we0),
    .tdf10_filters_address1(grp_td_fused_fu_990_tdf10_filters_address1),
    .tdf10_filters_ce1(grp_td_fused_fu_990_tdf10_filters_ce1),
    .tdf10_filters_d1(grp_td_fused_fu_990_tdf10_filters_d1),
    .tdf10_filters_q1(64'd0),
    .tdf10_filters_we1(grp_td_fused_fu_990_tdf10_filters_we1),
    .tdf10_l2_filters_address0(grp_td_fused_fu_990_tdf10_l2_filters_address0),
    .tdf10_l2_filters_ce0(grp_td_fused_fu_990_tdf10_l2_filters_ce0),
    .tdf10_l2_filters_d0(grp_td_fused_fu_990_tdf10_l2_filters_d0),
    .tdf10_l2_filters_q0(tdf10_l2_filters_q0),
    .tdf10_l2_filters_we0(grp_td_fused_fu_990_tdf10_l2_filters_we0),
    .tdf10_l2_filters_address1(grp_td_fused_fu_990_tdf10_l2_filters_address1),
    .tdf10_l2_filters_ce1(grp_td_fused_fu_990_tdf10_l2_filters_ce1),
    .tdf10_l2_filters_d1(grp_td_fused_fu_990_tdf10_l2_filters_d1),
    .tdf10_l2_filters_q1(16'd0),
    .tdf10_l2_filters_we1(grp_td_fused_fu_990_tdf10_l2_filters_we1),
    .tdf11_filters_address0(grp_td_fused_fu_990_tdf11_filters_address0),
    .tdf11_filters_ce0(grp_td_fused_fu_990_tdf11_filters_ce0),
    .tdf11_filters_d0(grp_td_fused_fu_990_tdf11_filters_d0),
    .tdf11_filters_q0(tdf11_filters_q0),
    .tdf11_filters_we0(grp_td_fused_fu_990_tdf11_filters_we0),
    .tdf11_filters_address1(grp_td_fused_fu_990_tdf11_filters_address1),
    .tdf11_filters_ce1(grp_td_fused_fu_990_tdf11_filters_ce1),
    .tdf11_filters_d1(grp_td_fused_fu_990_tdf11_filters_d1),
    .tdf11_filters_q1(64'd0),
    .tdf11_filters_we1(grp_td_fused_fu_990_tdf11_filters_we1),
    .tdf11_l2_filters_address0(grp_td_fused_fu_990_tdf11_l2_filters_address0),
    .tdf11_l2_filters_ce0(grp_td_fused_fu_990_tdf11_l2_filters_ce0),
    .tdf11_l2_filters_d0(grp_td_fused_fu_990_tdf11_l2_filters_d0),
    .tdf11_l2_filters_q0(tdf11_l2_filters_q0),
    .tdf11_l2_filters_we0(grp_td_fused_fu_990_tdf11_l2_filters_we0),
    .tdf11_l2_filters_address1(grp_td_fused_fu_990_tdf11_l2_filters_address1),
    .tdf11_l2_filters_ce1(grp_td_fused_fu_990_tdf11_l2_filters_ce1),
    .tdf11_l2_filters_d1(grp_td_fused_fu_990_tdf11_l2_filters_d1),
    .tdf11_l2_filters_q1(16'd0),
    .tdf11_l2_filters_we1(grp_td_fused_fu_990_tdf11_l2_filters_we1),
    .tdf12_filters_address0(grp_td_fused_fu_990_tdf12_filters_address0),
    .tdf12_filters_ce0(grp_td_fused_fu_990_tdf12_filters_ce0),
    .tdf12_filters_d0(grp_td_fused_fu_990_tdf12_filters_d0),
    .tdf12_filters_q0(tdf12_filters_q0),
    .tdf12_filters_we0(grp_td_fused_fu_990_tdf12_filters_we0),
    .tdf12_filters_address1(grp_td_fused_fu_990_tdf12_filters_address1),
    .tdf12_filters_ce1(grp_td_fused_fu_990_tdf12_filters_ce1),
    .tdf12_filters_d1(grp_td_fused_fu_990_tdf12_filters_d1),
    .tdf12_filters_q1(16'd0),
    .tdf12_filters_we1(grp_td_fused_fu_990_tdf12_filters_we1),
    .tdf1_adjustments_address0(grp_td_fused_fu_990_tdf1_adjustments_address0),
    .tdf1_adjustments_ce0(grp_td_fused_fu_990_tdf1_adjustments_ce0),
    .tdf1_adjustments_d0(grp_td_fused_fu_990_tdf1_adjustments_d0),
    .tdf1_adjustments_q0(tdf1_adjustments_q0),
    .tdf1_adjustments_we0(grp_td_fused_fu_990_tdf1_adjustments_we0),
    .tdf1_adjustments_address1(grp_td_fused_fu_990_tdf1_adjustments_address1),
    .tdf1_adjustments_ce1(grp_td_fused_fu_990_tdf1_adjustments_ce1),
    .tdf1_adjustments_d1(grp_td_fused_fu_990_tdf1_adjustments_d1),
    .tdf1_adjustments_q1(48'd0),
    .tdf1_adjustments_we1(grp_td_fused_fu_990_tdf1_adjustments_we1),
    .tdf2_adjustments_address0(grp_td_fused_fu_990_tdf2_adjustments_address0),
    .tdf2_adjustments_ce0(grp_td_fused_fu_990_tdf2_adjustments_ce0),
    .tdf2_adjustments_d0(grp_td_fused_fu_990_tdf2_adjustments_d0),
    .tdf2_adjustments_q0(tdf2_adjustments_q0),
    .tdf2_adjustments_we0(grp_td_fused_fu_990_tdf2_adjustments_we0),
    .tdf2_adjustments_address1(grp_td_fused_fu_990_tdf2_adjustments_address1),
    .tdf2_adjustments_ce1(grp_td_fused_fu_990_tdf2_adjustments_ce1),
    .tdf2_adjustments_d1(grp_td_fused_fu_990_tdf2_adjustments_d1),
    .tdf2_adjustments_q1(48'd0),
    .tdf2_adjustments_we1(grp_td_fused_fu_990_tdf2_adjustments_we1),
    .tdf3_adjustments_address0(grp_td_fused_fu_990_tdf3_adjustments_address0),
    .tdf3_adjustments_ce0(grp_td_fused_fu_990_tdf3_adjustments_ce0),
    .tdf3_adjustments_d0(grp_td_fused_fu_990_tdf3_adjustments_d0),
    .tdf3_adjustments_q0(tdf3_adjustments_q0),
    .tdf3_adjustments_we0(grp_td_fused_fu_990_tdf3_adjustments_we0),
    .tdf3_adjustments_address1(grp_td_fused_fu_990_tdf3_adjustments_address1),
    .tdf3_adjustments_ce1(grp_td_fused_fu_990_tdf3_adjustments_ce1),
    .tdf3_adjustments_d1(grp_td_fused_fu_990_tdf3_adjustments_d1),
    .tdf3_adjustments_q1(48'd0),
    .tdf3_adjustments_we1(grp_td_fused_fu_990_tdf3_adjustments_we1),
    .tdf4_adjustments_address0(grp_td_fused_fu_990_tdf4_adjustments_address0),
    .tdf4_adjustments_ce0(grp_td_fused_fu_990_tdf4_adjustments_ce0),
    .tdf4_adjustments_d0(grp_td_fused_fu_990_tdf4_adjustments_d0),
    .tdf4_adjustments_q0(tdf4_adjustments_q0),
    .tdf4_adjustments_we0(grp_td_fused_fu_990_tdf4_adjustments_we0),
    .tdf4_adjustments_address1(grp_td_fused_fu_990_tdf4_adjustments_address1),
    .tdf4_adjustments_ce1(grp_td_fused_fu_990_tdf4_adjustments_ce1),
    .tdf4_adjustments_d1(grp_td_fused_fu_990_tdf4_adjustments_d1),
    .tdf4_adjustments_q1(48'd0),
    .tdf4_adjustments_we1(grp_td_fused_fu_990_tdf4_adjustments_we1),
    .tdf4_l2_adjustments_address0(grp_td_fused_fu_990_tdf4_l2_adjustments_address0),
    .tdf4_l2_adjustments_ce0(grp_td_fused_fu_990_tdf4_l2_adjustments_ce0),
    .tdf4_l2_adjustments_d0(grp_td_fused_fu_990_tdf4_l2_adjustments_d0),
    .tdf4_l2_adjustments_q0(tdf4_l2_adjustments_q0),
    .tdf4_l2_adjustments_we0(grp_td_fused_fu_990_tdf4_l2_adjustments_we0),
    .tdf4_l2_adjustments_address1(grp_td_fused_fu_990_tdf4_l2_adjustments_address1),
    .tdf4_l2_adjustments_ce1(grp_td_fused_fu_990_tdf4_l2_adjustments_ce1),
    .tdf4_l2_adjustments_d1(grp_td_fused_fu_990_tdf4_l2_adjustments_d1),
    .tdf4_l2_adjustments_q1(48'd0),
    .tdf4_l2_adjustments_we1(grp_td_fused_fu_990_tdf4_l2_adjustments_we1),
    .tdf5_adjustments_address0(grp_td_fused_fu_990_tdf5_adjustments_address0),
    .tdf5_adjustments_ce0(grp_td_fused_fu_990_tdf5_adjustments_ce0),
    .tdf5_adjustments_d0(grp_td_fused_fu_990_tdf5_adjustments_d0),
    .tdf5_adjustments_q0(tdf5_adjustments_q0),
    .tdf5_adjustments_we0(grp_td_fused_fu_990_tdf5_adjustments_we0),
    .tdf5_adjustments_address1(grp_td_fused_fu_990_tdf5_adjustments_address1),
    .tdf5_adjustments_ce1(grp_td_fused_fu_990_tdf5_adjustments_ce1),
    .tdf5_adjustments_d1(grp_td_fused_fu_990_tdf5_adjustments_d1),
    .tdf5_adjustments_q1(48'd0),
    .tdf5_adjustments_we1(grp_td_fused_fu_990_tdf5_adjustments_we1),
    .tdf6_adjustments_address0(grp_td_fused_fu_990_tdf6_adjustments_address0),
    .tdf6_adjustments_ce0(grp_td_fused_fu_990_tdf6_adjustments_ce0),
    .tdf6_adjustments_d0(grp_td_fused_fu_990_tdf6_adjustments_d0),
    .tdf6_adjustments_q0(tdf6_adjustments_q0),
    .tdf6_adjustments_we0(grp_td_fused_fu_990_tdf6_adjustments_we0),
    .tdf6_adjustments_address1(grp_td_fused_fu_990_tdf6_adjustments_address1),
    .tdf6_adjustments_ce1(grp_td_fused_fu_990_tdf6_adjustments_ce1),
    .tdf6_adjustments_d1(grp_td_fused_fu_990_tdf6_adjustments_d1),
    .tdf6_adjustments_q1(48'd0),
    .tdf6_adjustments_we1(grp_td_fused_fu_990_tdf6_adjustments_we1),
    .tdf7_adjustments_address0(grp_td_fused_fu_990_tdf7_adjustments_address0),
    .tdf7_adjustments_ce0(grp_td_fused_fu_990_tdf7_adjustments_ce0),
    .tdf7_adjustments_d0(grp_td_fused_fu_990_tdf7_adjustments_d0),
    .tdf7_adjustments_q0(tdf7_adjustments_q0),
    .tdf7_adjustments_we0(grp_td_fused_fu_990_tdf7_adjustments_we0),
    .tdf7_adjustments_address1(grp_td_fused_fu_990_tdf7_adjustments_address1),
    .tdf7_adjustments_ce1(grp_td_fused_fu_990_tdf7_adjustments_ce1),
    .tdf7_adjustments_d1(grp_td_fused_fu_990_tdf7_adjustments_d1),
    .tdf7_adjustments_q1(48'd0),
    .tdf7_adjustments_we1(grp_td_fused_fu_990_tdf7_adjustments_we1),
    .tdf7_l2_adjustments_address0(grp_td_fused_fu_990_tdf7_l2_adjustments_address0),
    .tdf7_l2_adjustments_ce0(grp_td_fused_fu_990_tdf7_l2_adjustments_ce0),
    .tdf7_l2_adjustments_d0(grp_td_fused_fu_990_tdf7_l2_adjustments_d0),
    .tdf7_l2_adjustments_q0(tdf7_l2_adjustments_q0),
    .tdf7_l2_adjustments_we0(grp_td_fused_fu_990_tdf7_l2_adjustments_we0),
    .tdf7_l2_adjustments_address1(grp_td_fused_fu_990_tdf7_l2_adjustments_address1),
    .tdf7_l2_adjustments_ce1(grp_td_fused_fu_990_tdf7_l2_adjustments_ce1),
    .tdf7_l2_adjustments_d1(grp_td_fused_fu_990_tdf7_l2_adjustments_d1),
    .tdf7_l2_adjustments_q1(48'd0),
    .tdf7_l2_adjustments_we1(grp_td_fused_fu_990_tdf7_l2_adjustments_we1),
    .tdf8_adjustments_address0(grp_td_fused_fu_990_tdf8_adjustments_address0),
    .tdf8_adjustments_ce0(grp_td_fused_fu_990_tdf8_adjustments_ce0),
    .tdf8_adjustments_d0(grp_td_fused_fu_990_tdf8_adjustments_d0),
    .tdf8_adjustments_q0(tdf8_adjustments_q0),
    .tdf8_adjustments_we0(grp_td_fused_fu_990_tdf8_adjustments_we0),
    .tdf8_adjustments_address1(grp_td_fused_fu_990_tdf8_adjustments_address1),
    .tdf8_adjustments_ce1(grp_td_fused_fu_990_tdf8_adjustments_ce1),
    .tdf8_adjustments_d1(grp_td_fused_fu_990_tdf8_adjustments_d1),
    .tdf8_adjustments_q1(48'd0),
    .tdf8_adjustments_we1(grp_td_fused_fu_990_tdf8_adjustments_we1),
    .tdf9_adjustments_address0(grp_td_fused_fu_990_tdf9_adjustments_address0),
    .tdf9_adjustments_ce0(grp_td_fused_fu_990_tdf9_adjustments_ce0),
    .tdf9_adjustments_d0(grp_td_fused_fu_990_tdf9_adjustments_d0),
    .tdf9_adjustments_q0(tdf9_adjustments_q0),
    .tdf9_adjustments_we0(grp_td_fused_fu_990_tdf9_adjustments_we0),
    .tdf9_adjustments_address1(grp_td_fused_fu_990_tdf9_adjustments_address1),
    .tdf9_adjustments_ce1(grp_td_fused_fu_990_tdf9_adjustments_ce1),
    .tdf9_adjustments_d1(grp_td_fused_fu_990_tdf9_adjustments_d1),
    .tdf9_adjustments_q1(48'd0),
    .tdf9_adjustments_we1(grp_td_fused_fu_990_tdf9_adjustments_we1),
    .tdf10_adjustments_address0(grp_td_fused_fu_990_tdf10_adjustments_address0),
    .tdf10_adjustments_ce0(grp_td_fused_fu_990_tdf10_adjustments_ce0),
    .tdf10_adjustments_d0(grp_td_fused_fu_990_tdf10_adjustments_d0),
    .tdf10_adjustments_q0(tdf10_adjustments_q0),
    .tdf10_adjustments_we0(grp_td_fused_fu_990_tdf10_adjustments_we0),
    .tdf10_adjustments_address1(grp_td_fused_fu_990_tdf10_adjustments_address1),
    .tdf10_adjustments_ce1(grp_td_fused_fu_990_tdf10_adjustments_ce1),
    .tdf10_adjustments_d1(grp_td_fused_fu_990_tdf10_adjustments_d1),
    .tdf10_adjustments_q1(48'd0),
    .tdf10_adjustments_we1(grp_td_fused_fu_990_tdf10_adjustments_we1),
    .tdf10_l2_adjustments_address0(grp_td_fused_fu_990_tdf10_l2_adjustments_address0),
    .tdf10_l2_adjustments_ce0(grp_td_fused_fu_990_tdf10_l2_adjustments_ce0),
    .tdf10_l2_adjustments_d0(grp_td_fused_fu_990_tdf10_l2_adjustments_d0),
    .tdf10_l2_adjustments_q0(tdf10_l2_adjustments_q0),
    .tdf10_l2_adjustments_we0(grp_td_fused_fu_990_tdf10_l2_adjustments_we0),
    .tdf10_l2_adjustments_address1(grp_td_fused_fu_990_tdf10_l2_adjustments_address1),
    .tdf10_l2_adjustments_ce1(grp_td_fused_fu_990_tdf10_l2_adjustments_ce1),
    .tdf10_l2_adjustments_d1(grp_td_fused_fu_990_tdf10_l2_adjustments_d1),
    .tdf10_l2_adjustments_q1(48'd0),
    .tdf10_l2_adjustments_we1(grp_td_fused_fu_990_tdf10_l2_adjustments_we1),
    .tdf11_adjustments_address0(grp_td_fused_fu_990_tdf11_adjustments_address0),
    .tdf11_adjustments_ce0(grp_td_fused_fu_990_tdf11_adjustments_ce0),
    .tdf11_adjustments_d0(grp_td_fused_fu_990_tdf11_adjustments_d0),
    .tdf11_adjustments_q0(tdf11_adjustments_q0),
    .tdf11_adjustments_we0(grp_td_fused_fu_990_tdf11_adjustments_we0),
    .tdf11_adjustments_address1(grp_td_fused_fu_990_tdf11_adjustments_address1),
    .tdf11_adjustments_ce1(grp_td_fused_fu_990_tdf11_adjustments_ce1),
    .tdf11_adjustments_d1(grp_td_fused_fu_990_tdf11_adjustments_d1),
    .tdf11_adjustments_q1(48'd0),
    .tdf11_adjustments_we1(grp_td_fused_fu_990_tdf11_adjustments_we1),
    .tdf11_l2_adjustments_address0(grp_td_fused_fu_990_tdf11_l2_adjustments_address0),
    .tdf11_l2_adjustments_ce0(grp_td_fused_fu_990_tdf11_l2_adjustments_ce0),
    .tdf11_l2_adjustments_d0(grp_td_fused_fu_990_tdf11_l2_adjustments_d0),
    .tdf11_l2_adjustments_q0(tdf11_l2_adjustments_q0),
    .tdf11_l2_adjustments_we0(grp_td_fused_fu_990_tdf11_l2_adjustments_we0),
    .tdf11_l2_adjustments_address1(grp_td_fused_fu_990_tdf11_l2_adjustments_address1),
    .tdf11_l2_adjustments_ce1(grp_td_fused_fu_990_tdf11_l2_adjustments_ce1),
    .tdf11_l2_adjustments_d1(grp_td_fused_fu_990_tdf11_l2_adjustments_d1),
    .tdf11_l2_adjustments_q1(48'd0),
    .tdf11_l2_adjustments_we1(grp_td_fused_fu_990_tdf11_l2_adjustments_we1),
    .tdf12_adjustments_address0(grp_td_fused_fu_990_tdf12_adjustments_address0),
    .tdf12_adjustments_ce0(grp_td_fused_fu_990_tdf12_adjustments_ce0),
    .tdf12_adjustments_d0(grp_td_fused_fu_990_tdf12_adjustments_d0),
    .tdf12_adjustments_q0(tdf12_adjustments_q0),
    .tdf12_adjustments_we0(grp_td_fused_fu_990_tdf12_adjustments_we0),
    .tdf12_adjustments_address1(grp_td_fused_fu_990_tdf12_adjustments_address1),
    .tdf12_adjustments_ce1(grp_td_fused_fu_990_tdf12_adjustments_ce1),
    .tdf12_adjustments_d1(grp_td_fused_fu_990_tdf12_adjustments_d1),
    .tdf12_adjustments_q1(48'd0),
    .tdf12_adjustments_we1(grp_td_fused_fu_990_tdf12_adjustments_we1),
    .stream_in_TDATA(stream_in_TDATA_int_regslice),
    .stream_in_TKEEP(stream_in_TKEEP_int_regslice),
    .stream_in_TSTRB(stream_in_TSTRB_int_regslice),
    .stream_in_TLAST(stream_in_TLAST_int_regslice),
    .stream_out_TDATA(grp_td_fused_fu_990_stream_out_TDATA),
    .stream_out_TKEEP(grp_td_fused_fu_990_stream_out_TKEEP),
    .stream_out_TSTRB(grp_td_fused_fu_990_stream_out_TSTRB),
    .stream_out_TLAST(grp_td_fused_fu_990_stream_out_TLAST),
    .stream_in_TVALID(stream_in_TVALID_int_regslice),
    .stream_in_TREADY(grp_td_fused_fu_990_stream_in_TREADY),
    .ap_start(grp_td_fused_fu_990_ap_start),
    .stream_out_TVALID(grp_td_fused_fu_990_stream_out_TVALID),
    .stream_out_TREADY(grp_td_fused_fu_990_stream_out_TREADY),
    .ap_done(grp_td_fused_fu_990_ap_done),
    .ap_ready(grp_td_fused_fu_990_ap_ready),
    .ap_idle(grp_td_fused_fu_990_ap_idle),
    .ap_continue(grp_td_fused_fu_990_ap_continue)
);

td_fused_top_regslice_both #(
    .DataWidth( 16 ))
regslice_both_stream_in_V_data_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(stream_in_TDATA),
    .vld_in(stream_in_TVALID),
    .ack_in(regslice_both_stream_in_V_data_V_U_ack_in),
    .data_out(stream_in_TDATA_int_regslice),
    .vld_out(stream_in_TVALID_int_regslice),
    .ack_out(stream_in_TREADY_int_regslice),
    .apdone_blk(regslice_both_stream_in_V_data_V_U_apdone_blk)
);

td_fused_top_regslice_both #(
    .DataWidth( 2 ))
regslice_both_stream_in_V_keep_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(stream_in_TKEEP),
    .vld_in(stream_in_TVALID),
    .ack_in(regslice_both_stream_in_V_keep_V_U_ack_in),
    .data_out(stream_in_TKEEP_int_regslice),
    .vld_out(regslice_both_stream_in_V_keep_V_U_vld_out),
    .ack_out(stream_in_TREADY_int_regslice),
    .apdone_blk(regslice_both_stream_in_V_keep_V_U_apdone_blk)
);

td_fused_top_regslice_both #(
    .DataWidth( 2 ))
regslice_both_stream_in_V_strb_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(stream_in_TSTRB),
    .vld_in(stream_in_TVALID),
    .ack_in(regslice_both_stream_in_V_strb_V_U_ack_in),
    .data_out(stream_in_TSTRB_int_regslice),
    .vld_out(regslice_both_stream_in_V_strb_V_U_vld_out),
    .ack_out(stream_in_TREADY_int_regslice),
    .apdone_blk(regslice_both_stream_in_V_strb_V_U_apdone_blk)
);

td_fused_top_regslice_both #(
    .DataWidth( 1 ))
regslice_both_stream_in_V_last_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(stream_in_TLAST),
    .vld_in(stream_in_TVALID),
    .ack_in(regslice_both_stream_in_V_last_V_U_ack_in),
    .data_out(stream_in_TLAST_int_regslice),
    .vld_out(regslice_both_stream_in_V_last_V_U_vld_out),
    .ack_out(stream_in_TREADY_int_regslice),
    .apdone_blk(regslice_both_stream_in_V_last_V_U_apdone_blk)
);

td_fused_top_regslice_both #(
    .DataWidth( 16 ))
regslice_both_stream_out_V_data_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(grp_td_fused_fu_990_stream_out_TDATA),
    .vld_in(grp_td_fused_fu_990_stream_out_TVALID),
    .ack_in(stream_out_TREADY_int_regslice),
    .data_out(stream_out_TDATA),
    .vld_out(regslice_both_stream_out_V_data_V_U_vld_out),
    .ack_out(stream_out_TREADY),
    .apdone_blk(regslice_both_stream_out_V_data_V_U_apdone_blk)
);

td_fused_top_regslice_both #(
    .DataWidth( 2 ))
regslice_both_stream_out_V_keep_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(grp_td_fused_fu_990_stream_out_TKEEP),
    .vld_in(grp_td_fused_fu_990_stream_out_TVALID),
    .ack_in(regslice_both_stream_out_V_keep_V_U_ack_in_dummy),
    .data_out(stream_out_TKEEP),
    .vld_out(regslice_both_stream_out_V_keep_V_U_vld_out),
    .ack_out(stream_out_TREADY),
    .apdone_blk(regslice_both_stream_out_V_keep_V_U_apdone_blk)
);

td_fused_top_regslice_both #(
    .DataWidth( 2 ))
regslice_both_stream_out_V_strb_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(grp_td_fused_fu_990_stream_out_TSTRB),
    .vld_in(grp_td_fused_fu_990_stream_out_TVALID),
    .ack_in(regslice_both_stream_out_V_strb_V_U_ack_in_dummy),
    .data_out(stream_out_TSTRB),
    .vld_out(regslice_both_stream_out_V_strb_V_U_vld_out),
    .ack_out(stream_out_TREADY),
    .apdone_blk(regslice_both_stream_out_V_strb_V_U_apdone_blk)
);

td_fused_top_regslice_both #(
    .DataWidth( 1 ))
regslice_both_stream_out_V_last_V_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .data_in(grp_td_fused_fu_990_stream_out_TLAST),
    .vld_in(grp_td_fused_fu_990_stream_out_TVALID),
    .ack_in(regslice_both_stream_out_V_last_V_U_ack_in_dummy),
    .data_out(stream_out_TLAST),
    .vld_out(regslice_both_stream_out_V_last_V_U_vld_out),
    .ack_out(stream_out_TREADY),
    .apdone_blk(regslice_both_stream_out_V_last_V_U_apdone_blk)
);

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        ap_sync_reg_grp_td_fused_fu_990_ap_done <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_state4_on_subcall_done) & (1'b1 == ap_CS_fsm_state4))) begin
            ap_sync_reg_grp_td_fused_fu_990_ap_done <= 1'b0;
        end else if ((grp_td_fused_fu_990_ap_done == 1'b1)) begin
            ap_sync_reg_grp_td_fused_fu_990_ap_done <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        ap_sync_reg_grp_td_fused_fu_990_ap_ready <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_state4_on_subcall_done) & (1'b1 == ap_CS_fsm_state4))) begin
            ap_sync_reg_grp_td_fused_fu_990_ap_ready <= 1'b0;
        end else if ((grp_td_fused_fu_990_ap_ready == 1'b1)) begin
            ap_sync_reg_grp_td_fused_fu_990_ap_ready <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        grp_td_fused_fu_990_ap_start_reg <= 1'b0;
    end else begin
        if (((1'b1 == ap_CS_fsm_state3) | ((ap_sync_grp_td_fused_fu_990_ap_ready == 1'b0) & (1'b1 == ap_CS_fsm_state4)))) begin
            grp_td_fused_fu_990_ap_start_reg <= 1'b1;
        end else if ((grp_td_fused_fu_990_ap_ready == 1'b1)) begin
            grp_td_fused_fu_990_ap_start_reg <= 1'b0;
        end
    end
end

always @ (*) begin
    if (((regslice_both_stream_out_V_data_V_U_apdone_blk == 1'b0) & (1'b1 == ap_CS_fsm_state5))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((regslice_both_stream_out_V_data_V_U_apdone_blk == 1'b0) & (1'b1 == ap_CS_fsm_state5))) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_state4_on_subcall_done) & (1'b1 == ap_CS_fsm_state4))) begin
        grp_td_fused_fu_990_ap_continue = 1'b1;
    end else begin
        grp_td_fused_fu_990_ap_continue = 1'b0;
    end
end

always @ (*) begin
    if (((stream_in_TVALID_int_regslice == 1'b1) & (1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1))) begin
        stream_in_TREADY_int_regslice = 1'b1;
    end else if ((1'b1 == ap_CS_fsm_state4)) begin
        stream_in_TREADY_int_regslice = grp_td_fused_fu_990_stream_in_TREADY;
    end else begin
        stream_in_TREADY_int_regslice = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        tdf10_adjustments_ce0 = grp_td_fused_fu_990_tdf10_adjustments_ce0;
    end else begin
        tdf10_adjustments_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state2) | ((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)))) begin
        tdf10_adjustments_ce1 = 1'b1;
    end else begin
        tdf10_adjustments_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1))) begin
        tdf10_adjustments_we1 = 1'b1;
    end else begin
        tdf10_adjustments_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        tdf10_filters_ce0 = grp_td_fused_fu_990_tdf10_filters_ce0;
    end else begin
        tdf10_filters_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state2) | ((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)))) begin
        tdf10_filters_ce1 = 1'b1;
    end else begin
        tdf10_filters_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1))) begin
        tdf10_filters_we1 = 1'b1;
    end else begin
        tdf10_filters_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        tdf10_l2_adjustments_ce0 = grp_td_fused_fu_990_tdf10_l2_adjustments_ce0;
    end else begin
        tdf10_l2_adjustments_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state2) | ((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)))) begin
        tdf10_l2_adjustments_ce1 = 1'b1;
    end else begin
        tdf10_l2_adjustments_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1))) begin
        tdf10_l2_adjustments_we1 = 1'b1;
    end else begin
        tdf10_l2_adjustments_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        tdf10_l2_filters_ce0 = grp_td_fused_fu_990_tdf10_l2_filters_ce0;
    end else begin
        tdf10_l2_filters_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state2) | ((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)))) begin
        tdf10_l2_filters_ce1 = 1'b1;
    end else begin
        tdf10_l2_filters_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1))) begin
        tdf10_l2_filters_we1 = 1'b1;
    end else begin
        tdf10_l2_filters_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        tdf11_adjustments_ce0 = grp_td_fused_fu_990_tdf11_adjustments_ce0;
    end else begin
        tdf11_adjustments_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state2) | ((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)))) begin
        tdf11_adjustments_ce1 = 1'b1;
    end else begin
        tdf11_adjustments_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1))) begin
        tdf11_adjustments_we1 = 1'b1;
    end else begin
        tdf11_adjustments_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        tdf11_filters_ce0 = grp_td_fused_fu_990_tdf11_filters_ce0;
    end else begin
        tdf11_filters_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state2) | ((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)))) begin
        tdf11_filters_ce1 = 1'b1;
    end else begin
        tdf11_filters_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1))) begin
        tdf11_filters_we1 = 1'b1;
    end else begin
        tdf11_filters_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        tdf11_l2_adjustments_ce0 = grp_td_fused_fu_990_tdf11_l2_adjustments_ce0;
    end else begin
        tdf11_l2_adjustments_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state2) | ((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)))) begin
        tdf11_l2_adjustments_ce1 = 1'b1;
    end else begin
        tdf11_l2_adjustments_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1))) begin
        tdf11_l2_adjustments_we1 = 1'b1;
    end else begin
        tdf11_l2_adjustments_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        tdf11_l2_filters_ce0 = grp_td_fused_fu_990_tdf11_l2_filters_ce0;
    end else begin
        tdf11_l2_filters_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state2) | ((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)))) begin
        tdf11_l2_filters_ce1 = 1'b1;
    end else begin
        tdf11_l2_filters_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1))) begin
        tdf11_l2_filters_we1 = 1'b1;
    end else begin
        tdf11_l2_filters_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        tdf12_adjustments_ce0 = grp_td_fused_fu_990_tdf12_adjustments_ce0;
    end else begin
        tdf12_adjustments_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state2) | ((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)))) begin
        tdf12_adjustments_ce1 = 1'b1;
    end else begin
        tdf12_adjustments_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1))) begin
        tdf12_adjustments_we1 = 1'b1;
    end else begin
        tdf12_adjustments_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        tdf12_filters_ce0 = grp_td_fused_fu_990_tdf12_filters_ce0;
    end else begin
        tdf12_filters_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state2) | ((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)))) begin
        tdf12_filters_ce1 = 1'b1;
    end else begin
        tdf12_filters_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1))) begin
        tdf12_filters_we1 = 1'b1;
    end else begin
        tdf12_filters_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        tdf1_adjustments_ce0 = grp_td_fused_fu_990_tdf1_adjustments_ce0;
    end else begin
        tdf1_adjustments_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state2) | ((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)))) begin
        tdf1_adjustments_ce1 = 1'b1;
    end else begin
        tdf1_adjustments_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1))) begin
        tdf1_adjustments_we1 = 1'b1;
    end else begin
        tdf1_adjustments_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        tdf1_filters_ce0 = grp_td_fused_fu_990_tdf1_filters_ce0;
    end else begin
        tdf1_filters_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state2) | ((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)))) begin
        tdf1_filters_ce1 = 1'b1;
    end else begin
        tdf1_filters_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1))) begin
        tdf1_filters_we1 = 1'b1;
    end else begin
        tdf1_filters_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        tdf2_adjustments_ce0 = grp_td_fused_fu_990_tdf2_adjustments_ce0;
    end else begin
        tdf2_adjustments_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state2) | ((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)))) begin
        tdf2_adjustments_ce1 = 1'b1;
    end else begin
        tdf2_adjustments_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1))) begin
        tdf2_adjustments_we1 = 1'b1;
    end else begin
        tdf2_adjustments_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        tdf2_filters_ce0 = grp_td_fused_fu_990_tdf2_filters_ce0;
    end else begin
        tdf2_filters_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state2) | ((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)))) begin
        tdf2_filters_ce1 = 1'b1;
    end else begin
        tdf2_filters_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1))) begin
        tdf2_filters_we1 = 1'b1;
    end else begin
        tdf2_filters_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        tdf3_adjustments_ce0 = grp_td_fused_fu_990_tdf3_adjustments_ce0;
    end else begin
        tdf3_adjustments_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state2) | ((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)))) begin
        tdf3_adjustments_ce1 = 1'b1;
    end else begin
        tdf3_adjustments_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1))) begin
        tdf3_adjustments_we1 = 1'b1;
    end else begin
        tdf3_adjustments_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        tdf3_filters_ce0 = grp_td_fused_fu_990_tdf3_filters_ce0;
    end else begin
        tdf3_filters_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state2) | ((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)))) begin
        tdf3_filters_ce1 = 1'b1;
    end else begin
        tdf3_filters_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1))) begin
        tdf3_filters_we1 = 1'b1;
    end else begin
        tdf3_filters_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        tdf4_adjustments_ce0 = grp_td_fused_fu_990_tdf4_adjustments_ce0;
    end else begin
        tdf4_adjustments_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state2) | ((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)))) begin
        tdf4_adjustments_ce1 = 1'b1;
    end else begin
        tdf4_adjustments_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1))) begin
        tdf4_adjustments_we1 = 1'b1;
    end else begin
        tdf4_adjustments_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        tdf4_filters_ce0 = grp_td_fused_fu_990_tdf4_filters_ce0;
    end else begin
        tdf4_filters_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state2) | ((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)))) begin
        tdf4_filters_ce1 = 1'b1;
    end else begin
        tdf4_filters_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1))) begin
        tdf4_filters_we1 = 1'b1;
    end else begin
        tdf4_filters_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        tdf4_l2_adjustments_ce0 = grp_td_fused_fu_990_tdf4_l2_adjustments_ce0;
    end else begin
        tdf4_l2_adjustments_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state2) | ((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)))) begin
        tdf4_l2_adjustments_ce1 = 1'b1;
    end else begin
        tdf4_l2_adjustments_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1))) begin
        tdf4_l2_adjustments_we1 = 1'b1;
    end else begin
        tdf4_l2_adjustments_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        tdf4_l2_filters_ce0 = grp_td_fused_fu_990_tdf4_l2_filters_ce0;
    end else begin
        tdf4_l2_filters_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state2) | ((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)))) begin
        tdf4_l2_filters_ce1 = 1'b1;
    end else begin
        tdf4_l2_filters_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1))) begin
        tdf4_l2_filters_we1 = 1'b1;
    end else begin
        tdf4_l2_filters_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        tdf5_adjustments_ce0 = grp_td_fused_fu_990_tdf5_adjustments_ce0;
    end else begin
        tdf5_adjustments_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state2) | ((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)))) begin
        tdf5_adjustments_ce1 = 1'b1;
    end else begin
        tdf5_adjustments_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1))) begin
        tdf5_adjustments_we1 = 1'b1;
    end else begin
        tdf5_adjustments_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        tdf5_filters_ce0 = grp_td_fused_fu_990_tdf5_filters_ce0;
    end else begin
        tdf5_filters_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state2) | ((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)))) begin
        tdf5_filters_ce1 = 1'b1;
    end else begin
        tdf5_filters_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1))) begin
        tdf5_filters_we1 = 1'b1;
    end else begin
        tdf5_filters_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        tdf6_adjustments_ce0 = grp_td_fused_fu_990_tdf6_adjustments_ce0;
    end else begin
        tdf6_adjustments_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state2) | ((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)))) begin
        tdf6_adjustments_ce1 = 1'b1;
    end else begin
        tdf6_adjustments_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1))) begin
        tdf6_adjustments_we1 = 1'b1;
    end else begin
        tdf6_adjustments_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        tdf6_filters_ce0 = grp_td_fused_fu_990_tdf6_filters_ce0;
    end else begin
        tdf6_filters_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state2) | ((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)))) begin
        tdf6_filters_ce1 = 1'b1;
    end else begin
        tdf6_filters_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1))) begin
        tdf6_filters_we1 = 1'b1;
    end else begin
        tdf6_filters_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        tdf7_adjustments_ce0 = grp_td_fused_fu_990_tdf7_adjustments_ce0;
    end else begin
        tdf7_adjustments_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state2) | ((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)))) begin
        tdf7_adjustments_ce1 = 1'b1;
    end else begin
        tdf7_adjustments_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1))) begin
        tdf7_adjustments_we1 = 1'b1;
    end else begin
        tdf7_adjustments_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        tdf7_filters_ce0 = grp_td_fused_fu_990_tdf7_filters_ce0;
    end else begin
        tdf7_filters_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state2) | ((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)))) begin
        tdf7_filters_ce1 = 1'b1;
    end else begin
        tdf7_filters_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1))) begin
        tdf7_filters_we1 = 1'b1;
    end else begin
        tdf7_filters_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        tdf7_l2_adjustments_ce0 = grp_td_fused_fu_990_tdf7_l2_adjustments_ce0;
    end else begin
        tdf7_l2_adjustments_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state2) | ((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)))) begin
        tdf7_l2_adjustments_ce1 = 1'b1;
    end else begin
        tdf7_l2_adjustments_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1))) begin
        tdf7_l2_adjustments_we1 = 1'b1;
    end else begin
        tdf7_l2_adjustments_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        tdf7_l2_filters_ce0 = grp_td_fused_fu_990_tdf7_l2_filters_ce0;
    end else begin
        tdf7_l2_filters_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state2) | ((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)))) begin
        tdf7_l2_filters_ce1 = 1'b1;
    end else begin
        tdf7_l2_filters_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1))) begin
        tdf7_l2_filters_we1 = 1'b1;
    end else begin
        tdf7_l2_filters_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        tdf8_adjustments_ce0 = grp_td_fused_fu_990_tdf8_adjustments_ce0;
    end else begin
        tdf8_adjustments_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state2) | ((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)))) begin
        tdf8_adjustments_ce1 = 1'b1;
    end else begin
        tdf8_adjustments_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1))) begin
        tdf8_adjustments_we1 = 1'b1;
    end else begin
        tdf8_adjustments_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        tdf8_filters_ce0 = grp_td_fused_fu_990_tdf8_filters_ce0;
    end else begin
        tdf8_filters_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state2) | ((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)))) begin
        tdf8_filters_ce1 = 1'b1;
    end else begin
        tdf8_filters_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1))) begin
        tdf8_filters_we1 = 1'b1;
    end else begin
        tdf8_filters_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        tdf9_adjustments_ce0 = grp_td_fused_fu_990_tdf9_adjustments_ce0;
    end else begin
        tdf9_adjustments_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state2) | ((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)))) begin
        tdf9_adjustments_ce1 = 1'b1;
    end else begin
        tdf9_adjustments_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1))) begin
        tdf9_adjustments_we1 = 1'b1;
    end else begin
        tdf9_adjustments_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        tdf9_filters_ce0 = grp_td_fused_fu_990_tdf9_filters_ce0;
    end else begin
        tdf9_filters_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state2) | ((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)))) begin
        tdf9_filters_ce1 = 1'b1;
    end else begin
        tdf9_filters_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1))) begin
        tdf9_filters_we1 = 1'b1;
    end else begin
        tdf9_filters_we1 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_state2 : begin
            ap_NS_fsm = ap_ST_fsm_state3;
        end
        ap_ST_fsm_state3 : begin
            ap_NS_fsm = ap_ST_fsm_state4;
        end
        ap_ST_fsm_state4 : begin
            if (((1'b0 == ap_block_state4_on_subcall_done) & (1'b1 == ap_CS_fsm_state4))) begin
                ap_NS_fsm = ap_ST_fsm_state5;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end
        end
        ap_ST_fsm_state5 : begin
            if (((regslice_both_stream_out_V_data_V_U_apdone_blk == 1'b0) & (1'b1 == ap_CS_fsm_state5))) begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state5;
            end
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

assign ap_CS_fsm_state5 = ap_CS_fsm[32'd4];

always @ (*) begin
    ap_block_state4_on_subcall_done = ((ap_sync_grp_td_fused_fu_990_ap_ready & ap_sync_grp_td_fused_fu_990_ap_done) == 1'b0);
end

always @ (*) begin
    ap_rst_n_inv = ~ap_rst_n;
end

assign ap_sync_grp_td_fused_fu_990_ap_done = (grp_td_fused_fu_990_ap_done | ap_sync_reg_grp_td_fused_fu_990_ap_done);

assign ap_sync_grp_td_fused_fu_990_ap_ready = (grp_td_fused_fu_990_ap_ready | ap_sync_reg_grp_td_fused_fu_990_ap_ready);

assign grp_td_fused_fu_990_ap_start = grp_td_fused_fu_990_ap_start_reg;

assign grp_td_fused_fu_990_stream_out_TREADY = (stream_out_TREADY_int_regslice & ap_CS_fsm_state4);

assign stream_in_TREADY = regslice_both_stream_in_V_data_V_U_ack_in;

assign stream_out_TVALID = regslice_both_stream_out_V_data_V_U_vld_out;

assign tdf10_adjustments_address1 = 64'd0;

assign tdf10_filters_address1 = 64'd0;

assign tdf10_l2_adjustments_address1 = 64'd0;

assign tdf10_l2_filters_address1 = 64'd0;

assign tdf11_adjustments_address1 = 64'd0;

assign tdf11_filters_address1 = 64'd0;

assign tdf11_l2_adjustments_address1 = 64'd0;

assign tdf11_l2_filters_address1 = 64'd0;

assign tdf12_adjustments_address1 = 64'd0;

assign tdf12_filters_address1 = 64'd0;

assign tdf1_adjustments_address1 = 64'd0;

assign tdf1_filters_address1 = 64'd0;

assign tdf2_adjustments_address1 = 64'd0;

assign tdf2_filters_address1 = 64'd0;

assign tdf3_adjustments_address1 = 64'd0;

assign tdf3_filters_address1 = 64'd0;

assign tdf4_adjustments_address1 = 64'd0;

assign tdf4_filters_address1 = 64'd0;

assign tdf4_l2_adjustments_address1 = 64'd0;

assign tdf4_l2_filters_address1 = 64'd0;

assign tdf5_adjustments_address1 = 64'd0;

assign tdf5_filters_address1 = 64'd0;

assign tdf6_adjustments_address1 = 64'd0;

assign tdf6_filters_address1 = 64'd0;

assign tdf7_adjustments_address1 = 64'd0;

assign tdf7_filters_address1 = 64'd0;

assign tdf7_l2_adjustments_address1 = 64'd0;

assign tdf7_l2_filters_address1 = 64'd0;

assign tdf8_adjustments_address1 = 64'd0;

assign tdf8_filters_address1 = 64'd0;

assign tdf9_adjustments_address1 = 64'd0;

assign tdf9_filters_address1 = 64'd0;

assign tmp_data_fu_1262_p1 = stream_in_TDATA_int_regslice;

assign tmp_fu_1280_p5 = {{ap_const_lv64_0[63:16]}, {stream_in_TDATA_int_regslice}};

assign trunc_ln151_fu_1294_p1 = tmp_fu_1280_p5[47:0];

endmodule //td_fused_top


//////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////
// Floating point 16-bit multiplier
// This is a heavily modified version of:
// https://github.com/fbrosser/DSP48E1-FP/tree/master/src/FPMult
// Original author: Fredrik Brosser
// Abridged by: Samidh Mehta
//////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////

`ifndef complex_dsp

`define EXPONENT 5
`define MANTISSA 10
`define ACTUAL_MANTISSA 11
`define EXPONENT_LSB 10
`define EXPONENT_MSB 14
`define MANTISSA_LSB 0
`define MANTISSA_MSB 9
`define MANTISSA_MUL_SPLIT_LSB 3
`define MANTISSA_MUL_SPLIT_MSB 9
`define SIGN 1
`define SIGN_LOC 15
`define DWIDTH (`SIGN+`EXPONENT+`MANTISSA)
`define IEEE_COMPLIANCE 1

module FPMult_16(
		clk,
		rst,
		a,
		b,
		result,
		flags
    );
	
	// Input Ports
	input clk ;							// Clock
	input rst ;							// Reset signal
	input [`DWIDTH-1:0] a;					// Input A, a 32-bit floating point number
	input [`DWIDTH-1:0] b;					// Input B, a 32-bit floating point number
	
	// Output ports
	output [`DWIDTH-1:0] result ;					// Product, result of the operation, 32-bit FP number
	output [4:0] flags ;				// Flags indicating exceptions according to IEEE754
	
	// Internal signals
	wire [31:0] Z_int ;				// Product, result of the operation, 32-bit FP number
	wire [4:0] Flags_int ;			// Flags indicating exceptions according to IEEE754
	
	wire Sa ;							// A's sign
	wire Sb ;							// B's sign
	wire Sp ;							// Product sign
	wire [`EXPONENT-1:0] Ea ;					// A's exponent
	wire [`EXPONENT-1:0] Eb ;					// B's exponent
	wire [2*`MANTISSA+1:0] Mp ;					// Product mantissa
	wire [4:0] InputExc ;			// Exceptions in inputs
	wire [`MANTISSA-1:0] NormM ;				// Normalized mantissa
	wire [`EXPONENT:0] NormE ;				// Normalized exponent
	wire [`MANTISSA:0] RoundM ;				// Normalized mantissa
	wire [`EXPONENT:0] RoundE ;				// Normalized exponent
	wire [`MANTISSA:0] RoundMP ;				// Normalized mantissa
	wire [`EXPONENT:0] RoundEP ;				// Normalized exponent
	wire GRS ;

	//reg [63:0] pipe_0;			// Pipeline register Input->Prep
	reg [2*`DWIDTH-1:0] pipe_0;			// Pipeline register Input->Prep

	//reg [92:0] pipe_1;			// Pipeline register Prep->Execute
	reg [3*`MANTISSA+2*`EXPONENT+7:0] pipe_1;			// Pipeline register Prep->Execute

	//reg [38:0] pipe_2;			// Pipeline register Execute->Normalize
	reg [`MANTISSA+`EXPONENT+7:0] pipe_2;			// Pipeline register Execute->Normalize
	
	//reg [72:0] pipe_3;			// Pipeline register Normalize->Round
	reg [2*`MANTISSA+2*`EXPONENT+10:0] pipe_3;			// Pipeline register Normalize->Round

	//reg [36:0] pipe_4;			// Pipeline register Round->Output
	reg [`DWIDTH+4:0] pipe_4;			// Pipeline register Round->Output
	
	assign result = pipe_4[`DWIDTH+4:5] ;
	assign flags = pipe_4[4:0] ;
	
	// Prepare the operands for alignment and check for exceptions
	FPMult_PrepModule PrepModule(clk, rst, pipe_0[2*`DWIDTH-1:`DWIDTH], pipe_0[`DWIDTH-1:0], Sa, Sb, Ea[`EXPONENT-1:0], Eb[`EXPONENT-1:0], Mp[2*`MANTISSA+1:0], InputExc[4:0]) ;

	// Perform (unsigned) mantissa multiplication
	FPMult_ExecuteModule ExecuteModule(pipe_1[3*`MANTISSA+`EXPONENT*2+7:2*`MANTISSA+2*`EXPONENT+8], pipe_1[2*`MANTISSA+2*`EXPONENT+7:2*`MANTISSA+7], pipe_1[2*`MANTISSA+6:5], pipe_1[2*`MANTISSA+2*`EXPONENT+6:2*`MANTISSA+`EXPONENT+7], pipe_1[2*`MANTISSA+`EXPONENT+6:2*`MANTISSA+7], pipe_1[2*`MANTISSA+2*`EXPONENT+8], pipe_1[2*`MANTISSA+2*`EXPONENT+7], Sp, NormE[`EXPONENT:0], NormM[`MANTISSA-1:0], GRS) ;

	// Round result and if necessary, perform a second (post-rounding) normalization step
	FPMult_NormalizeModule NormalizeModule(pipe_2[`MANTISSA-1:0], pipe_2[`MANTISSA+`EXPONENT:`MANTISSA], RoundE[`EXPONENT:0], RoundEP[`EXPONENT:0], RoundM[`MANTISSA:0], RoundMP[`MANTISSA:0]) ;		

	// Round result and if necessary, perform a second (post-rounding) normalization step
	//FPMult_RoundModule RoundModule(pipe_3[47:24], pipe_3[23:0], pipe_3[65:57], pipe_3[56:48], pipe_3[66], pipe_3[67], pipe_3[72:68], Z_int[31:0], Flags_int[4:0]) ;		
	FPMult_RoundModule RoundModule(pipe_3[2*`MANTISSA+1:`MANTISSA+1], pipe_3[`MANTISSA:0], pipe_3[2*`MANTISSA+2*`EXPONENT+3:2*`MANTISSA+`EXPONENT+3], pipe_3[2*`MANTISSA+`EXPONENT+2:2*`MANTISSA+2], pipe_3[2*`MANTISSA+2*`EXPONENT+4], pipe_3[2*`MANTISSA+2*`EXPONENT+5], pipe_3[2*`MANTISSA+2*`EXPONENT+10:2*`MANTISSA+2*`EXPONENT+6], Z_int[`DWIDTH-1:0], Flags_int[4:0]) ;		

	always @ (*) begin	
		if(rst) begin
			pipe_0 = 0;
			pipe_1 = 0;
			pipe_2 = 0; 
			pipe_3 = 0;
			pipe_4 = 0;
		end 
		else begin		
			/* PIPE 0
				[63:32] A
				[31:0] B
			*/
      pipe_0 = {a, b} ;

			/* PIPE 1
				[70] Sa
				[69] Sb
				[68:61] Ea
				[60:53] Eb
				[52:5] Mp
				[4:0] InputExc
			*/
			//pipe_1 <= {pipe_0[`DWIDTH+`MANTISSA-1:`DWIDTH], pipe_0[`MANTISSA_MUL_SPLIT_LSB-1:0], Sa, Sb, Ea[`EXPONENT-1:0], Eb[`EXPONENT-1:0], Mp[2*`MANTISSA-1:0], InputExc[4:0]} ;
			pipe_1 = {pipe_0[`DWIDTH+`MANTISSA-1:`DWIDTH], pipe_0[8:0], Sa, Sb, Ea[`EXPONENT-1:0], Eb[`EXPONENT-1:0], Mp[2*`MANTISSA+1:0], InputExc[4:0]} ;
			/* PIPE 2
				[38:34] InputExc
				[33] GRS
				[32] Sp
				[31:23] NormE
				[22:0] NormM
			*/
			pipe_2 = {pipe_1[4:0], GRS, Sp, NormE[`EXPONENT:0], NormM[`MANTISSA-1:0]} ;
			/* PIPE 3
				[72:68] InputExc
				[67] GRS
				[66] Sp	
				[65:57] RoundE
				[56:48] RoundEP
				[47:24] RoundM
				[23:0] RoundMP
			*/
			pipe_3 = {pipe_2[`EXPONENT+`MANTISSA+7:`EXPONENT+`MANTISSA+1], RoundE[`EXPONENT:0], RoundEP[`EXPONENT:0], RoundM[`MANTISSA:0], RoundMP[`MANTISSA:0]} ;
			/* PIPE 4
				[36:5] Z
				[4:0] Flags
			*/				
			pipe_4 = {Z_int[`DWIDTH-1:0], Flags_int[4:0]} ;
		end
	end
		
endmodule


module FPMult_PrepModule (
		clk,
		rst,
		a,
		b,
		Sa,
		Sb,
		Ea,
		Eb,
		Mp,
		InputExc
	);
	
	// Input ports
	input clk ;
	input rst ;
	input [`DWIDTH-1:0] a ;								// Input A, a 32-bit floating point number
	input [`DWIDTH-1:0] b ;								// Input B, a 32-bit floating point number
	
	// Output ports
	output Sa ;										// A's sign
	output Sb ;										// B's sign
	output [`EXPONENT-1:0] Ea ;								// A's exponent
	output [`EXPONENT-1:0] Eb ;								// B's exponent
	output [2*`MANTISSA+1:0] Mp ;							// Mantissa product
	output [4:0] InputExc ;						// Input numbers are exceptions
	
	// Internal signals							// If signal is high...
	wire ANaN ;										// A is a signalling NaN
	wire BNaN ;										// B is a signalling NaN
	wire AInf ;										// A is infinity
	wire BInf ;										// B is infinity
    wire [`MANTISSA-1:0] Ma;
    wire [`MANTISSA-1:0] Mb;
	
	assign ANaN = &(a[`DWIDTH-2:`MANTISSA]) &  |(a[`DWIDTH-2:`MANTISSA]) ;			// All one exponent and not all zero mantissa - NaN
	assign BNaN = &(b[`DWIDTH-2:`MANTISSA]) &  |(b[`MANTISSA-1:0]);			// All one exponent and not all zero mantissa - NaN
	assign AInf = &(a[`DWIDTH-2:`MANTISSA]) & ~|(a[`DWIDTH-2:`MANTISSA]) ;		// All one exponent and all zero mantissa - Infinity
	assign BInf = &(b[`DWIDTH-2:`MANTISSA]) & ~|(b[`DWIDTH-2:`MANTISSA]) ;		// All one exponent and all zero mantissa - Infinity
	
	// Check for any exceptions and put all flags into exception vector
	assign InputExc = {(ANaN | BNaN | AInf | BInf), ANaN, BNaN, AInf, BInf} ;
	//assign InputExc = {(ANaN | ANaN | BNaN |BNaN), ANaN, ANaN, BNaN,BNaN} ;
	
	// Take input numbers apart
	assign Sa = a[`DWIDTH-1] ;							// A's sign
	assign Sb = b[`DWIDTH-1] ;							// B's sign
	assign Ea = a[`DWIDTH-2:`MANTISSA];						// Store A's exponent in Ea, unless A is an exception
	assign Eb = b[`DWIDTH-2:`MANTISSA];						// Store B's exponent in Eb, unless B is an exception	
//    assign Ma = a[`MANTISSA_MSB:`MANTISSA_LSB];
  //  assign Mb = b[`MANTISSA_MSB:`MANTISSA_LSB];
	


	//assign Mp = ({4'b0001, a[`MANTISSA-1:0]}*{4'b0001, b[`MANTISSA-1:9]}) ;
	assign Mp = ({1'b1,a[`MANTISSA-1:0]}*{1'b1, b[`MANTISSA-1:0]}) ;

	
    //We multiply part of the mantissa here
    //Full mantissa of A
    //Bits MANTISSA_MUL_SPLIT_MSB:MANTISSA_MUL_SPLIT_LSB of B
   // wire [`ACTUAL_MANTISSA-1:0] inp_A;
   // wire [`ACTUAL_MANTISSA-1:0] inp_B;
   // assign inp_A = {1'b1, Ma};
   // assign inp_B = {{(`MANTISSA-(`MANTISSA_MUL_SPLIT_MSB-`MANTISSA_MUL_SPLIT_LSB+1)){1'b0}}, 1'b1, Mb[`MANTISSA_MUL_SPLIT_MSB:`MANTISSA_MUL_SPLIT_LSB]};
   // DW02_mult #(`ACTUAL_MANTISSA,`ACTUAL_MANTISSA) u_mult(.A(inp_A), .B(inp_B), .TC(1'b0), .PRODUCT(Mp));
endmodule


module FPMult_ExecuteModule(
		a,
		b,
		MpC,
		Ea,
		Eb,
		Sa,
		Sb,
		Sp,
		NormE,
		NormM,
		GRS
    );

	// Input ports
	input [`MANTISSA-1:0] a ;
	input [2*`EXPONENT:0] b ;
	input [2*`MANTISSA+1:0] MpC ;
	input [`EXPONENT-1:0] Ea ;						// A's exponent
	input [`EXPONENT-1:0] Eb ;						// B's exponent
	input Sa ;								// A's sign
	input Sb ;								// B's sign
	
	// Output ports
	output Sp ;								// Product sign
	output [`EXPONENT:0] NormE ;													// Normalized exponent
	output [`MANTISSA-1:0] NormM ;												// Normalized mantissa
	output GRS ;
	
	wire [2*`MANTISSA+1:0] Mp ;
	
	assign Sp = (Sa ^ Sb) ;												// Equal signs give a positive product
	
   // wire [`ACTUAL_MANTISSA-1:0] inp_a;
   // wire [`ACTUAL_MANTISSA-1:0] inp_b;
   // assign inp_a = {1'b1, a};
   // assign inp_b = {{(`MANTISSA-`MANTISSA_MUL_SPLIT_LSB){1'b0}}, 1'b0, b};
   // DW02_mult #(`ACTUAL_MANTISSA,`ACTUAL_MANTISSA) u_mult(.A(inp_a), .B(inp_b), .TC(1'b0), .PRODUCT(Mp_temp));
   // DW01_add #(2*`ACTUAL_MANTISSA) u_add(.A(Mp_temp), .B(MpC<<`MANTISSA_MUL_SPLIT_LSB), .CI(1'b0), .SUM(Mp), .CO());

	//assign Mp = (MpC<<(2*`EXPONENT+1)) + ({4'b0001, a[`MANTISSA-1:0]}*{1'b0, b[2*`EXPONENT:0]}) ;
	assign Mp = MpC;


	assign NormM = (Mp[2*`MANTISSA+1] ? Mp[2*`MANTISSA:`MANTISSA+1] : Mp[2*`MANTISSA-1:`MANTISSA]); 	// Check for overflow
	assign NormE = (Ea + Eb + Mp[2*`MANTISSA+1]);								// If so, increment exponent
	
	assign GRS = ((Mp[`MANTISSA]&(Mp[`MANTISSA+1]))|(|Mp[`MANTISSA-1:0])) ;
	
endmodule

module FPMult_NormalizeModule(
		NormM,
		NormE,
		RoundE,
		RoundEP,
		RoundM,
		RoundMP
    );

	// Input Ports
	input [`MANTISSA-1:0] NormM ;									// Normalized mantissa
	input [`EXPONENT:0] NormE ;									// Normalized exponent

	// Output Ports
	output [`EXPONENT:0] RoundE ;
	output [`EXPONENT:0] RoundEP ;
	output [`MANTISSA:0] RoundM ;
	output [`MANTISSA:0] RoundMP ; 
	
	assign RoundE = NormE - 15 ;
	assign RoundEP = NormE - 14 ;
	assign RoundM = NormM ;
	assign RoundMP = NormM ;

endmodule

module FPMult_RoundModule(
		RoundM,
		RoundMP,
		RoundE,
		RoundEP,
		Sp,
		GRS,
		InputExc,
		Z,
		Flags
    );

	// Input Ports
	input [`MANTISSA:0] RoundM ;									// Normalized mantissa
	input [`MANTISSA:0] RoundMP ;									// Normalized exponent
	input [`EXPONENT:0] RoundE ;									// Normalized mantissa + 1
	input [`EXPONENT:0] RoundEP ;									// Normalized exponent + 1
	input Sp ;												// Product sign
	input GRS ;
	input [4:0] InputExc ;
	
	// Output Ports
	output [`DWIDTH-1:0] Z ;										// Final product
	output [4:0] Flags ;
	
	// Internal Signals
	wire [`EXPONENT:0] FinalE ;									// Rounded exponent
	wire [`MANTISSA:0] FinalM;
	wire [`MANTISSA:0] PreShiftM;
	
	assign PreShiftM = GRS ? RoundMP : RoundM ;	// Round up if R and (G or S)
	
	// Post rounding normalization (potential one bit shift> use shifted mantissa if there is overflow)
	assign FinalM = (PreShiftM[`MANTISSA] ? {1'b0, PreShiftM[`MANTISSA:1]} : PreShiftM[`MANTISSA:0]) ;
	
	assign FinalE = (PreShiftM[`MANTISSA] ? RoundEP : RoundE) ; // Increment exponent if a shift was done
	
	assign Z = {Sp, FinalE[`EXPONENT-1:0], FinalM[`MANTISSA-1:0]} ;   // Putting the pieces together
	assign Flags = InputExc[4:0];

endmodule

//////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////
// Definition of a 16-bit floating point adder/subtractor
// This is a heavily modified version of:
// https://github.com/fbrosser/DSP48E1-FP/tree/master/src/FP_AddSub
// Original author: Fredrik Brosser
// Abridged by: Samidh Mehta
//////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////

module FPAddSub(
		clk,
		rst,
		a,
		b,
		operation,			// 0 add, 1 sub
		result,
		flags
	);
	
	// Clock and reset
	input clk ;										// Clock signal
	input rst ;										// Reset (active high, resets pipeline registers)
	
	// Input ports
	input [`DWIDTH-1:0] a ;								// Input A, a 32-bit floating point number
	input [`DWIDTH-1:0] b ;								// Input B, a 32-bit floating point number
	input operation ;								// Operation select signal
	
	// Output ports
	output [`DWIDTH-1:0] result ;						// Result of the operation
	output [4:0] flags ;							// Flags indicating exceptions according to IEEE754
	
	// Pipeline Registers
	//reg [79:0] pipe_1;							// Pipeline register PreAlign->Align1
	reg [`DWIDTH*2+15:0] pipe_1;							// Pipeline register PreAlign->Align1

	//reg [67:0] pipe_2;							// Pipeline register Align1->Align3
	reg [`MANTISSA*2+`EXPONENT+13:0] pipe_2;							// Pipeline register Align1->Align3

	//reg [76:0] pipe_3;	68						// Pipeline register Align1->Align3
	reg [`MANTISSA*2+`EXPONENT+14:0] pipe_3;							// Pipeline register Align1->Align3

	//reg [69:0] pipe_4;							// Pipeline register Align3->Execute
	reg [`MANTISSA*2+`EXPONENT+15:0] pipe_4;							// Pipeline register Align3->Execute

	//reg [51:0] pipe_5;							// Pipeline register Execute->Normalize
	reg [`DWIDTH+`EXPONENT+11:0] pipe_5;							// Pipeline register Execute->Normalize

	//reg [56:0] pipe_6;							// Pipeline register Nomalize->NormalizeShift1
	reg [`DWIDTH+`EXPONENT+16:0] pipe_6;							// Pipeline register Nomalize->NormalizeShift1

	//reg [56:0] pipe_7;							// Pipeline register NormalizeShift2->NormalizeShift3
	reg [`DWIDTH+`EXPONENT+16:0] pipe_7;							// Pipeline register NormalizeShift2->NormalizeShift3

	//reg [54:0] pipe_8;							// Pipeline register NormalizeShift3->Round
	reg [`EXPONENT*2+`MANTISSA+15:0] pipe_8;							// Pipeline register NormalizeShift3->Round

	//reg [40:0] pipe_9;							// Pipeline register NormalizeShift3->Round
	reg [`DWIDTH+8:0] pipe_9;							// Pipeline register NormalizeShift3->Round
	
	// Internal wires between modules
	wire [`DWIDTH-2:0] Aout_0 ;							// A - sign
	wire [`DWIDTH-2:0] Bout_0 ;							// B - sign
	wire Opout_0 ;									// A's sign
	wire Sa_0 ;										// A's sign
	wire Sb_0 ;										// B's sign
	wire MaxAB_1 ;									// Indicates the larger of A and B(0/A, 1/B)
	wire [`EXPONENT-1:0] CExp_1 ;							// Common Exponent
	wire [4:0] Shift_1 ;							// Number of steps to smaller mantissa shift right (align)
	wire [`MANTISSA-1:0] Mmax_1 ;							// Larger mantissa
	wire [4:0] InputExc_0 ;						// Input numbers are exceptions
	wire [9:0] ShiftDet_0 ;
	wire [`MANTISSA-1:0] MminS_1 ;						// Smaller mantissa after 0/16 shift
	wire [`MANTISSA:0] MminS_2 ;						// Smaller mantissa after 0/4/8/12 shift
	wire [`MANTISSA:0] Mmin_3 ;							// Smaller mantissa after 0/1/2/3 shift
	wire [`DWIDTH:0] Sum_4 ;
	wire PSgn_4 ;
	wire Opr_4 ;
	wire [4:0] Shift_5 ;							// Number of steps to shift sum left (normalize)
	wire [`DWIDTH:0] SumS_5 ;							// Sum after 0/16 shift
	wire [`DWIDTH:0] SumS_6 ;							// Sum after 0/16 shift
	wire [`DWIDTH:0] SumS_7 ;							// Sum after 0/16 shift
	wire [`MANTISSA-1:0] NormM_8 ;						// Normalized mantissa
	wire [`EXPONENT:0] NormE_8;							// Adjusted exponent
	wire ZeroSum_8 ;								// Zero flag
	wire NegE_8 ;									// Flag indicating negative exponent
	wire R_8 ;										// Round bit
	wire S_8 ;										// Final sticky bit
	wire FG_8 ;										// Final sticky bit
	wire [`DWIDTH-1:0] P_int ;
	wire EOF ;
	
	// Prepare the operands for alignment and check for exceptions
	FPAddSub_PrealignModule PrealignModule
	(	// Inputs
		a, b, operation,
		// Outputs
		Sa_0, Sb_0, ShiftDet_0[9:0], InputExc_0[4:0], Aout_0[`DWIDTH-2:0], Bout_0[`DWIDTH-2:0], Opout_0) ;
		
	// Prepare the operands for alignment and check for exceptions
	FPAddSub_AlignModule AlignModule
	(	// Inputs
		pipe_1[14+2*`DWIDTH:16+`DWIDTH], pipe_1[15+`DWIDTH:17], pipe_1[14:5],
		// Outputs
		CExp_1[`EXPONENT-1:0], MaxAB_1, Shift_1[4:0], MminS_1[`MANTISSA-1:0], Mmax_1[`MANTISSA-1:0]) ;	

	// Alignment Shift Stage 1
	FPAddSub_AlignShift1 AlignShift1
	(  // Inputs
		pipe_2[`MANTISSA-1:0], pipe_2[2*`MANTISSA+9:2*`MANTISSA+7],
		// Outputs
		MminS_2[`MANTISSA:0]) ;

	// Alignment Shift Stage 3 and compution of guard and sticky bits
	FPAddSub_AlignShift2 AlignShift2  
	(  // Inputs
		pipe_3[`MANTISSA:0], pipe_3[2*`MANTISSA+7:2*`MANTISSA+6],
		// Outputs
		Mmin_3[`MANTISSA:0]) ;
						
	// Perform mantissa addition
	FPAddSub_ExecutionModule ExecutionModule
	(  // Inputs
		pipe_4[`MANTISSA*2+5:`MANTISSA+6], pipe_4[`MANTISSA:0], pipe_4[`MANTISSA*2+`EXPONENT+13], pipe_4[`MANTISSA*2+`EXPONENT+12], pipe_4[`MANTISSA*2+`EXPONENT+11], pipe_4[`MANTISSA*2+`EXPONENT+14],
		// Outputs
		Sum_4[`DWIDTH:0], PSgn_4, Opr_4) ;
	
	// Prepare normalization of result
	FPAddSub_NormalizeModule NormalizeModule
	(  // Inputs
		pipe_5[`DWIDTH:0], 
		// Outputs
		SumS_5[`DWIDTH:0], Shift_5[4:0]) ;
					
	// Normalization Shift Stage 1
	FPAddSub_NormalizeShift1 NormalizeShift1
	(  // Inputs
		pipe_6[`DWIDTH:0], pipe_6[`DWIDTH+`EXPONENT+14:`DWIDTH+`EXPONENT+11],
		// Outputs
		SumS_7[`DWIDTH:0]) ;
		
	// Normalization Shift Stage 3 and final guard, sticky and round bits
	FPAddSub_NormalizeShift2 NormalizeShift2
	(  // Inputs
		pipe_7[`DWIDTH:0], pipe_7[`DWIDTH+`EXPONENT+5:`DWIDTH+6], pipe_7[`DWIDTH+`EXPONENT+15:`DWIDTH+`EXPONENT+11],
		// Outputs
		NormM_8[`MANTISSA-1:0], NormE_8[`EXPONENT:0], ZeroSum_8, NegE_8, R_8, S_8, FG_8) ;

	// Round and put result together
	FPAddSub_RoundModule RoundModule
	(  // Inputs
		 pipe_8[3], pipe_8[4+`EXPONENT:4], pipe_8[`EXPONENT+`MANTISSA+4:5+`EXPONENT], pipe_8[1], pipe_8[0], pipe_8[`EXPONENT*2+`MANTISSA+15], pipe_8[`EXPONENT*2+`MANTISSA+12], pipe_8[`EXPONENT*2+`MANTISSA+11], pipe_8[`EXPONENT*2+`MANTISSA+14], pipe_8[`EXPONENT*2+`MANTISSA+10], 
		// Outputs
		P_int[`DWIDTH-1:0], EOF) ;
	
	// Check for exceptions
	FPAddSub_ExceptionModule Exceptionmodule
	(  // Inputs
		pipe_9[8+`DWIDTH:9], pipe_9[8], pipe_9[7], pipe_9[6], pipe_9[5:1], pipe_9[0], 
		// Outputs
		result[`DWIDTH-1:0], flags[4:0]) ;			
	
	always @ (*) begin	
		if(rst) begin
			pipe_1 = 0;
			pipe_2 = 0;
			pipe_3 = 0;
			pipe_4 = 0;
			pipe_5 = 0;
			pipe_6 = 0;
			pipe_7 = 0;
			pipe_8 = 0;
			pipe_9 = 0;
		end 
		else begin
		
			pipe_1 = {Opout_0, Aout_0[`DWIDTH-2:0], Bout_0[`DWIDTH-2:0], Sa_0, Sb_0, ShiftDet_0[9:0], InputExc_0[4:0]} ;	
			// PIPE_2 :
			//[67] operation
			//[66] Sa_0
			//[65] Sb_0
			//[64] MaxAB_0
			//[63:56] CExp_0
			//[55:51] Shift_0
			//[50:28] Mmax_0
			//[27:23] InputExc_0
			//[22:0] MminS_1
			//
			pipe_2 = {pipe_1[`DWIDTH*2+15], pipe_1[16:15], MaxAB_1, CExp_1[`EXPONENT-1:0], Shift_1[4:0], Mmax_1[`MANTISSA-1:0], pipe_1[4:0], MminS_1[`MANTISSA-1:0]} ;	
			// PIPE_3 :
			//[68] operation
			//[67] Sa_0
			//[66] Sb_0
			//[65] MaxAB_0
			//[64:57] CExp_0
			//[56:52] Shift_0
			//[51:29] Mmax_0
			//[28:24] InputExc_0
			//[23:0] MminS_1
			//
			pipe_3 = {pipe_2[`MANTISSA*2+`EXPONENT+13:`MANTISSA], MminS_2[`MANTISSA:0]} ;	
			// PIPE_4 :
			//[68] operation
			//[67] Sa_0
			//[66] Sb_0
			//[65] MaxAB_0
			//[64:57] CExp_0
			//[56:52] Shift_0
			//[51:29] Mmax_0
			//[28:24] InputExc_0
			//[23:0] Mmin_3
			//					
			pipe_4 = {pipe_3[`MANTISSA*2+`EXPONENT+14:`MANTISSA+1], Mmin_3[`MANTISSA:0]} ;	
			// PIPE_5 :
			//[51] operation
			//[50] PSgn_4
			//[49] Opr_4
			//[48] Sa_0
			//[47] Sb_0
			//[46] MaxAB_0
			//[45:38] CExp_0
			//[37:33] InputExc_0
			//[32:0] Sum_4
			//					
			pipe_5 = {pipe_4[2*`MANTISSA+`EXPONENT+14], PSgn_4, Opr_4, pipe_4[2*`MANTISSA+`EXPONENT+13:2*`MANTISSA+11], pipe_4[`MANTISSA+5:`MANTISSA+1], Sum_4[`DWIDTH:0]} ;
			// PIPE_6 :
			//[56] operation
			//[55:51] Shift_5
			//[50] PSgn_4
			//[49] Opr_4
			//[48] Sa_0
			//[47] Sb_0
			//[46] MaxAB_0
			//[45:38] CExp_0
			//[37:33] InputExc_0
			//[32:0] Sum_4
			//					
			pipe_6 = {pipe_5[`EXPONENT+`EXPONENT+11], Shift_5[4:0], pipe_5[`DWIDTH+`EXPONENT+10:`DWIDTH+1], SumS_5[`DWIDTH:0]} ;	
			// pipe_7 :
			//[56] operation
			//[55:51] Shift_5
			//[50] PSgn_4
			//[49] Opr_4
			//[48] Sa_0
			//[47] Sb_0
			//[46] MaxAB_0
			//[45:38] CExp_0
			//[37:33] InputExc_0
			//[32:0] Sum_4
			//						
			pipe_7 = {pipe_6[`DWIDTH+`EXPONENT+16:`DWIDTH+1], SumS_7[`DWIDTH:0]} ;	
			// pipe_8:
			//[54] FG_8 
			//[53] operation
			//[52] PSgn_4
			//[51] Sa_0
			//[50] Sb_0
			//[49] MaxAB_0
			//[48:41] CExp_0
			//[40:36] InputExc_8
			//[35:13] NormM_8 
			//[12:4] NormE_8
			//[3] ZeroSum_8
			//[2] NegE_8
			//[1] R_8
			//[0] S_8
			//				
			pipe_8 = {FG_8, pipe_7[`DWIDTH+`EXPONENT+16], pipe_7[`DWIDTH+`EXPONENT+10], pipe_7[`DWIDTH+`EXPONENT+8:`DWIDTH+1], NormM_8[`MANTISSA-1:0], NormE_8[`EXPONENT:0], ZeroSum_8, NegE_8, R_8, S_8} ;	
			// pipe_9:
			//[40:9] P_int
			//[8] NegE_8
			//[7] R_8
			//[6] S_8
			//[5:1] InputExc_8
			//[0] EOF
			//				
			pipe_9 = {P_int[`DWIDTH-1:0], pipe_8[2], pipe_8[1], pipe_8[0], pipe_8[`EXPONENT+`MANTISSA+9:`EXPONENT+`MANTISSA+5], EOF} ;	
		end
	end		
	
endmodule

// Description:	 	The pre-alignment module is responsible for taking the inputs
//							apart and checking the parts for exceptions.
//							The exponent difference is also calculated in this module.

module FPAddSub_PrealignModule(
		A,
		B,
		operation,
		Sa,
		Sb,
		ShiftDet,
		InputExc,
		Aout,
		Bout,
		Opout
	);
	
	// Input ports
	input [`DWIDTH-1:0] A ;										// Input A, a 32-bit floating point number
	input [`DWIDTH-1:0] B ;										// Input B, a 32-bit floating point number
	input operation ;
	
	// Output ports
	output Sa ;												// A's sign
	output Sb ;												// B's sign
	output [9:0] ShiftDet ;
	output [4:0] InputExc ;								// Input numbers are exceptions
	output [`DWIDTH-2:0] Aout ;
	output [`DWIDTH-2:0] Bout ;
	output Opout ;
	
	// Internal signals									// If signal is high...
	wire ANaN ;												// A is a NaN (Not-a-Number)
	wire BNaN ;												// B is a NaN
	wire AInf ;												// A is infinity
	wire BInf ;												// B is infinity
	wire [`EXPONENT-1:0] DAB ;										// ExpA - ExpB					
	wire [`EXPONENT-1:0] DBA ;										// ExpB - ExpA	
	
	assign ANaN = &(A[`DWIDTH-2:`DWIDTH-1-`EXPONENT]) & |(A[`MANTISSA-1:0]) ;		// All one exponent and not all zero mantissa - NaN
	assign BNaN = &(B[`DWIDTH-2:`DWIDTH-1-`EXPONENT]) & |(B[`MANTISSA-1:0]);		// All one exponent and not all zero mantissa - NaN
	assign AInf = &(A[`DWIDTH-2:`DWIDTH-1-`EXPONENT]) & ~|(A[`MANTISSA-1:0]) ;	// All one exponent and all zero mantissa - Infinity
	assign BInf = &(B[`DWIDTH-2:`DWIDTH-1-`EXPONENT]) & ~|(B[`MANTISSA-1:0]) ;	// All one exponent and all zero mantissa - Infinity
	
	// Put all flags into exception vector
	assign InputExc = {(ANaN | BNaN | AInf | BInf), ANaN, BNaN, AInf, BInf} ;
	
	//assign DAB = (A[30:23] - B[30:23]) ;
	//assign DBA = (B[30:23] - A[30:23]) ;
	assign DAB = (A[`DWIDTH-2:`MANTISSA] + ~(B[`DWIDTH-2:`MANTISSA]) + 1) ;
	assign DBA = (B[`DWIDTH-2:`MANTISSA] + ~(A[`DWIDTH-2:`MANTISSA]) + 1) ;
	
	assign Sa = A[`DWIDTH-1] ;									// A's sign bit
	assign Sb = B[`DWIDTH-1] ;									// B's sign	bit
	assign ShiftDet = {DBA[4:0], DAB[4:0]} ;		// Shift data
	assign Opout = operation ;
	assign Aout = A[`DWIDTH-2:0] ;
	assign Bout = B[`DWIDTH-2:0] ;
	
endmodule

// Description:	 	The alignment module determines the larger input operand and
//							sets the mantissas, shift and common exponent accordingly.

module FPAddSub_AlignModule (
		A,
		B,
		ShiftDet,
		CExp,
		MaxAB,
		Shift,
		Mmin,
		Mmax
	);
	
	// Input ports
	input [`DWIDTH-2:0] A ;								// Input A, a 32-bit floating point number
	input [`DWIDTH-2:0] B ;								// Input B, a 32-bit floating point number
	input [9:0] ShiftDet ;
	
	// Output ports
	output [`EXPONENT-1:0] CExp ;							// Common Exponent
	output MaxAB ;									// Incidates larger of A and B (0/A, 1/B)
	output [4:0] Shift ;							// Number of steps to smaller mantissa shift right
	output [`MANTISSA-1:0] Mmin ;							// Smaller mantissa 
	output [`MANTISSA-1:0] Mmax ;							// Larger mantissa
	
	// Internal signals
	//wire BOF ;										// Check for shifting overflow if B is larger
	//wire AOF ;										// Check for shifting overflow if A is larger
	
	assign MaxAB = (A[`DWIDTH-2:0] < B[`DWIDTH-2:0]) ;	
	//assign BOF = ShiftDet[9:5] < 25 ;		// Cannot shift more than 25 bits
	//assign AOF = ShiftDet[4:0] < 25 ;		// Cannot shift more than 25 bits
	
	// Determine final shift value
	//assign Shift = MaxAB ? (BOF ? ShiftDet[9:5] : 5'b11001) : (AOF ? ShiftDet[4:0] : 5'b11001) ;
	
	assign Shift = MaxAB ? ShiftDet[9:5] : ShiftDet[4:0] ;
	
	// Take out smaller mantissa and append shift space
	assign Mmin = MaxAB ? A[`MANTISSA-1:0] : B[`MANTISSA-1:0] ; 
	
	// Take out larger mantissa	
	assign Mmax = MaxAB ? B[`MANTISSA-1:0]: A[`MANTISSA-1:0] ;	
	
	// Common exponent
	assign CExp = (MaxAB ? B[`MANTISSA+`EXPONENT-1:`MANTISSA] : A[`MANTISSA+`EXPONENT-1:`MANTISSA]) ;		
	
endmodule

// Description:	 Alignment shift stage 1, performs 16|12|8|4 shift

module FPAddSub_AlignShift1(
		MminP,
		Shift,
		Mmin
	);
	
	// Input ports
	input [`MANTISSA-1:0] MminP ;						// Smaller mantissa after 16|12|8|4 shift
	input [2:0] Shift ;						// Shift amount
	
	// Output ports
	output [`MANTISSA:0] Mmin ;						// The smaller mantissa
	
	// Internal signals
	reg	  [`MANTISSA:0]		Lvl1;
	reg	  [`MANTISSA:0]		Lvl2;
	wire    [2*`MANTISSA+1:0]    Stage1;	
	integer           i;                // Loop variable
	
	always @(*) begin						
		// Rotate by 16?
		//Lvl1 <= Shift[2] ? {17'b00000000000000001, MminP[22:16]} : {1'b1, MminP}; 
		Lvl1 <= Shift[2] ? {11'b0000000000} : {1'b1, MminP}; 
		
	end
	
	assign Stage1 = { 11'b0, Lvl1};
	
	always @(*) begin    					// Rotate {0 | 4 | 8 | 12} bits
	  case (Shift[1:0])
			// Rotate by 0	
			2'b00:  Lvl2 <= Stage1[`MANTISSA:0];       			
			// Rotate by 4	
			2'b01:  begin for (i=0; i<=`MANTISSA; i=i+1) begin Lvl2[i] <= Stage1[i+4]; end /*Lvl2[`MANTISSA:`MANTISSA-3] <= 0;*/ end
			// Rotate by 8
			2'b10:  begin for (i=0; i<=`MANTISSA; i=i+1) begin Lvl2[i] <= Stage1[i+8]; end /*Lvl2[`MANTISSA:`MANTISSA-7] <= 0;*/ end
			// Rotate by 12	
			2'b11: Lvl2[`MANTISSA: 0] <= 0; 
			//2'b11:  begin for (i=0; i<=`MANTISSA; i=i+1) begin Lvl2[i] <= Stage1[i+12]; end Lvl2[`MANTISSA:`MANTISSA-12] <= 0; end
	  endcase
	end
	
	// Assign output to next shift stage
	assign Mmin = Lvl2;
	
endmodule

// Description:	 Alignment shift stage 2, performs 3|2|1 shift

module FPAddSub_AlignShift2(
		MminP,
		Shift,
		Mmin
	);
	
	// Input ports
	input [`MANTISSA:0] MminP ;						// Smaller mantissa after 16|12|8|4 shift
	input [1:0] Shift ;						// Shift amount
	
	// Output ports
	output [`MANTISSA:0] Mmin ;						// The smaller mantissa
	
	// Internal Signal
	reg	  [`MANTISSA:0]		Lvl3;
	wire    [2*`MANTISSA+1:0]    Stage2;	
	integer           j;               // Loop variable
	
	assign Stage2 = {11'b0, MminP};

	always @(*) begin    // Rotate {0 | 1 | 2 | 3} bits
	  case (Shift[1:0])
			// Rotate by 0
			2'b00:  Lvl3 <= Stage2[`MANTISSA:0];   
			// Rotate by 1
			2'b01:  begin for (j=0; j<=`MANTISSA; j=j+1)  begin Lvl3[j] <= Stage2[j+1]; end /*Lvl3[`MANTISSA] <= 0; */end 
			// Rotate by 2
			2'b10:  begin for (j=0; j<=`MANTISSA; j=j+1)  begin Lvl3[j] <= Stage2[j+2]; end /*Lvl3[`MANTISSA:`MANTISSA-1] <= 0;*/ end 
			// Rotate by 3
			2'b11:  begin for (j=0; j<=`MANTISSA; j=j+1)  begin Lvl3[j] <= Stage2[j+3]; end /*Lvl3[`MANTISSA:`MANTISSA-2] <= 0;*/ end 	  
	  endcase
	end
	
	// Assign output
	assign Mmin = Lvl3;						// Take out smaller mantissa				

endmodule

// Description:	 Module that executes the addition or subtraction on mantissas.

module FPAddSub_ExecutionModule(
		Mmax,
		Mmin,
		Sa,
		Sb,
		MaxAB,
		OpMode,
		Sum,
		PSgn,
		Opr
    );

	// Input ports
	input [`MANTISSA-1:0] Mmax ;					// The larger mantissa
	input [`MANTISSA:0] Mmin ;					// The smaller mantissa
	input Sa ;								// Sign bit of larger number
	input Sb ;								// Sign bit of smaller number
	input MaxAB ;							// Indicates the larger number (0/A, 1/B)
	input OpMode ;							// Operation to be performed (0/Add, 1/Sub)
	
	// Output ports
	output [`DWIDTH:0] Sum ;					// The result of the operation
	output PSgn ;							// The sign for the result
	output Opr ;							// The effective (performed) operation

	assign Opr = (OpMode^Sa^Sb); 		// Resolve sign to determine operation

	// Perform effective operation
	assign Sum = (OpMode^Sa^Sb) ? ({1'b1, Mmax, 5'b00000} - {Mmin, 5'b00000}) : ({1'b1, Mmax, 5'b00000} + {Mmin, 5'b00000}) ;
	
	// Assign result sign
	assign PSgn = (MaxAB ? Sb : Sa) ;

endmodule

// Description:	 Determine the normalization shift amount and perform 16-shift

module FPAddSub_NormalizeModule(
		Sum,
		Mmin,
		Shift
    );

	// Input ports
	input [`DWIDTH:0] Sum ;					// Mantissa sum including hidden 1 and GRS
	
	// Output ports
	output [`DWIDTH:0] Mmin ;					// Mantissa after 16|0 shift
	output [4:0] Shift ;					// Shift amount
	
	// Determine normalization shift amount by finding leading nought
	assign Shift =  ( 
		Sum[16] ? 5'b00000 :	 
		Sum[15] ? 5'b00001 : 
		Sum[14] ? 5'b00010 : 
		Sum[13] ? 5'b00011 : 
		Sum[12] ? 5'b00100 : 
		Sum[11] ? 5'b00101 : 
		Sum[10] ? 5'b00110 : 
		Sum[9] ? 5'b00111 :
		Sum[8] ? 5'b01000 :
		Sum[7] ? 5'b01001 :
		Sum[6] ? 5'b01010 :
		Sum[5] ? 5'b01011 :
		Sum[4] ? 5'b01100 : 5'b01101
	//	Sum[19] ? 5'b01101 :
	//	Sum[18] ? 5'b01110 :
	//	Sum[17] ? 5'b01111 :
	//	Sum[16] ? 5'b10000 :
	//	Sum[15] ? 5'b10001 :
	//	Sum[14] ? 5'b10010 :
	//	Sum[13] ? 5'b10011 :
	//	Sum[12] ? 5'b10100 :
	//	Sum[11] ? 5'b10101 :
	//	Sum[10] ? 5'b10110 :
	//	Sum[9] ? 5'b10111 :
	//	Sum[8] ? 5'b11000 :
	//	Sum[7] ? 5'b11001 : 5'b11010
	);
	
	reg	  [`DWIDTH:0]		Lvl1;
	
	always @(*) begin
		// Rotate by 16?
		Lvl1 <= Shift[4] ? {Sum[8:0], 8'b00000000} : Sum; 
	end
	
	// Assign outputs
	assign Mmin = Lvl1;						// Take out smaller mantissa

endmodule

// Description:	 Normalization shift stage 1, performs 12|8|4|3|2|1|0 shift

module FPAddSub_NormalizeShift1(
		MminP,
		Shift,
		Mmin
	);
	
	// Input ports
	input [`DWIDTH:0] MminP ;						// Smaller mantissa after 16|12|8|4 shift
	input [3:0] Shift ;						// Shift amount
	
	// Output ports
	output [`DWIDTH:0] Mmin ;						// The smaller mantissa
	
	reg	  [`DWIDTH:0]		Lvl2;
	wire    [2*`DWIDTH+1:0]    Stage1;	
	reg	  [`DWIDTH:0]		Lvl3;
	wire    [2*`DWIDTH+1:0]    Stage2;	
	integer           i;               	// Loop variable
	
	assign Stage1 = {MminP, MminP};

	always @(*) begin    					// Rotate {0 | 4 | 8 | 12} bits
	  case (Shift[3:2])
			// Rotate by 0
			2'b00: //Lvl2 <= Stage1[`DWIDTH:0];       		
      begin Lvl2 = Stage1[`DWIDTH:0];  end
			// Rotate by 4
			2'b01: //begin for (i=2*`DWIDTH+1; i>=`DWIDTH+1; i=i-1) begin Lvl2[i-33] <= Stage1[i-4]; end Lvl2[3:0] <= 0; end
      begin Lvl2[`DWIDTH: (`DWIDTH-4)] = Stage1[3:0]; Lvl2[`DWIDTH-4-1:0] = Stage1[`DWIDTH-4]; end
			// Rotate by 8
			2'b10: //begin for (i=2*`DWIDTH+1; i>=`DWIDTH+1; i=i-1) begin Lvl2[i-33] <= Stage1[i-8]; end Lvl2[7:0] <= 0; end
      begin Lvl2[`DWIDTH: (`DWIDTH-8)] = Stage1[3:0]; Lvl2[`DWIDTH-8-1:0] = Stage1[`DWIDTH-8]; end
			// Rotate by 12
			2'b11: //begin for (i=2*`DWIDTH+1; i>=`DWIDTH+1; i=i-1) begin Lvl2[i-33] <= Stage1[i-12]; end Lvl2[11:0] <= 0; end
      begin Lvl2[`DWIDTH: (`DWIDTH-12)] = Stage1[3:0]; Lvl2[`DWIDTH-12-1:0] = Stage1[`DWIDTH-12]; end
	  endcase
	end
	
	assign Stage2 = {Lvl2, Lvl2};

	always @(*) begin   				 		// Rotate {0 | 1 | 2 | 3} bits
	  case (Shift[1:0])
			// Rotate by 0
			2'b00:  //Lvl3 <= Stage2[`DWIDTH:0];
      begin Lvl3 = Stage2[`DWIDTH:0]; end
			// Rotate by 1
			2'b01: //begin for (i=2*`DWIDTH+1; i>=`DWIDTH+1; i=i-1) begin Lvl3[i-`DWIDTH-1] <= Stage2[i-1]; end Lvl3[0] <= 0; end 
      begin Lvl3[`DWIDTH: (`DWIDTH-1)] = Stage2[3:0]; Lvl3[`DWIDTH-1-1:0] = Stage2[`DWIDTH-1]; end
			// Rotate by 2
			2'b10: //begin for (i=2*`DWIDTH+1; i>=`DWIDTH+1; i=i-1) begin Lvl3[i-`DWIDTH-1] <= Stage2[i-2]; end Lvl3[1:0] <= 0; end
      begin Lvl3[`DWIDTH: (`DWIDTH-2)] = Stage2[3:0]; Lvl3[`DWIDTH-2-1:0] = Stage2[`DWIDTH-2]; end
			// Rotate by 3
			2'b11: //begin for (i=2*`DWIDTH+1; i>=`DWIDTH+1; i=i-1) begin Lvl3[i-`DWIDTH-1] <= Stage2[i-3]; end Lvl3[2:0] <= 0; end
      begin Lvl3[`DWIDTH: (`DWIDTH-3)] = Stage2[3:0]; Lvl3[`DWIDTH-3-1:0] = Stage2[`DWIDTH-3]; end
	  endcase
	end
	
	// Assign outputs
	assign Mmin = Lvl3;						// Take out smaller mantissa			
	
endmodule

// Description:	 Normalization shift stage 2, calculates post-normalization
//						 mantissa and exponent, as well as the bits used in rounding		

module FPAddSub_NormalizeShift2(
		PSSum,
		CExp,
		Shift,
		NormM,
		NormE,
		ZeroSum,
		NegE,
		R,
		S,
		FG
	);
	
	// Input ports
	input [`DWIDTH:0] PSSum ;					// The Pre-Shift-Sum
	input [`EXPONENT-1:0] CExp ;
	input [4:0] Shift ;					// Amount to be shifted

	// Output ports
	output [`MANTISSA-1:0] NormM ;				// Normalized mantissa
	output [`EXPONENT:0] NormE ;					// Adjusted exponent
	output ZeroSum ;						// Zero flag
	output NegE ;							// Flag indicating negative exponent
	output R ;								// Round bit
	output S ;								// Final sticky bit
	output FG ;

	// Internal signals
	wire MSBShift ;						// Flag indicating that a second shift is needed
	wire [`EXPONENT:0] ExpOF ;					// MSB set in sum indicates overflow
	wire [`EXPONENT:0] ExpOK ;					// MSB not set, no adjustment
	
	// Calculate normalized exponent and mantissa, check for all-zero sum
	assign MSBShift = PSSum[`DWIDTH] ;		// Check MSB in unnormalized sum
	assign ZeroSum = ~|PSSum ;			// Check for all zero sum
	assign ExpOK = CExp - Shift ;		// Adjust exponent for new normalized mantissa
	assign NegE = ExpOK[`EXPONENT] ;			// Check for exponent overflow
	assign ExpOF = CExp - Shift + 1'b1 ;		// If MSB set, add one to exponent(x2)
	assign NormE = MSBShift ? ExpOF : ExpOK ;			// Check for exponent overflow
	assign NormM = PSSum[`DWIDTH-1:`EXPONENT+1] ;		// The new, normalized mantissa
	
	// Also need to compute sticky and round bits for the rounding stage
	assign FG = PSSum[`EXPONENT] ; 
	assign R = PSSum[`EXPONENT-1] ;
	assign S = |PSSum[`EXPONENT-2:0] ;
	
endmodule

// Description:	 Performs 'Round to nearest, tie to even'-rounding on the
//						 normalized mantissa according to the G, R, S bits. Calculates
//						 final result and checks for exponent overflow.

module FPAddSub_RoundModule(
		ZeroSum,
		NormE,
		NormM,
		R,
		S,
		G,
		Sa,
		Sb,
		Ctrl,
		MaxAB,
		Z,
		EOF
    );

	// Input ports
	input ZeroSum ;					// Sum is zero
	input [`EXPONENT:0] NormE ;				// Normalized exponent
	input [`MANTISSA-1:0] NormM ;				// Normalized mantissa
	input R ;							// Round bit
	input S ;							// Sticky bit
	input G ;
	input Sa ;							// A's sign bit
	input Sb ;							// B's sign bit
	input Ctrl ;						// Control bit (operation)
	input MaxAB ;
	
	// Output ports
	output [`DWIDTH-1:0] Z ;					// Final result
	output EOF ;
	
	// Internal signals
	wire [`MANTISSA:0] RoundUpM ;			// Rounded up sum with room for overflow
	wire [`MANTISSA-1:0] RoundM ;				// The final rounded sum
	wire [`EXPONENT:0] RoundE ;				// Rounded exponent (note extra bit due to poential overflow	)
	wire RoundUp ;						// Flag indicating that the sum should be rounded up
        wire FSgn;
	wire ExpAdd ;						// May have to add 1 to compensate for overflow 
	wire RoundOF ;						// Rounding overflow
	
	// The cases where we need to round upwards (= adding one) in Round to nearest, tie to even
	assign RoundUp = (G & ((R | S) | NormM[0])) ;
	
	// Note that in the other cases (rounding down), the sum is already 'rounded'
	assign RoundUpM = (NormM + 1) ;								// The sum, rounded up by 1
	assign RoundM = (RoundUp ? RoundUpM[`MANTISSA-1:0] : NormM) ; 	// Compute final mantissa	
	assign RoundOF = RoundUp & RoundUpM[`MANTISSA] ; 				// Check for overflow when rounding up

	// Calculate post-rounding exponent
	assign ExpAdd = (RoundOF ? 1'b1 : 1'b0) ; 				// Add 1 to exponent to compensate for overflow
	assign RoundE = ZeroSum ? 5'b00000 : (NormE + ExpAdd) ; 							// Final exponent

	// If zero, need to determine sign according to rounding
	assign FSgn = (ZeroSum & (Sa ^ Sb)) | (ZeroSum ? (Sa & Sb & ~Ctrl) : ((~MaxAB & Sa) | ((Ctrl ^ Sb) & (MaxAB | Sa)))) ;

	// Assign final result
	assign Z = {FSgn, RoundE[`EXPONENT-1:0], RoundM[`MANTISSA-1:0]} ;
	
	// Indicate exponent overflow
	assign EOF = RoundE[`EXPONENT];
	
endmodule

// Description:	 Check the final result for exception conditions and set
//						 flags accordingly.

module FPAddSub_ExceptionModule(
		Z,
		NegE,
		R,
		S,
		InputExc,
		EOF,
		P,
		Flags
    );
	 
	// Input ports
	input [`DWIDTH-1:0] Z	;					// Final product
	input NegE ;						// Negative exponent?
	input R ;							// Round bit
	input S ;							// Sticky bit
	input [4:0] InputExc ;			// Exceptions in inputs A and B
	input EOF ;
	
	// Output ports
	output [`DWIDTH-1:0] P ;					// Final result
	output [4:0] Flags ;				// Exception flags
	
	// Internal signals
	wire Overflow ;					// Overflow flag
	wire Underflow ;					// Underflow flag
	wire DivideByZero ;				// Divide-by-Zero flag (always 0 in Add/Sub)
	wire Invalid ;						// Invalid inputs or result
	wire Inexact ;						// Result is inexact because of rounding
	
	// Exception flags
	
	// Result is too big to be represented
	assign Overflow = EOF | InputExc[1] | InputExc[0] ;
	
	// Result is too small to be represented
	assign Underflow = NegE & (R | S);
	
	// Infinite result computed exactly from finite operands
	assign DivideByZero = &(Z[`MANTISSA+`EXPONENT-1:`MANTISSA]) & ~|(Z[`MANTISSA+`EXPONENT-1:`MANTISSA]) & ~InputExc[1] & ~InputExc[0];
	
	// Invalid inputs or operation
	assign Invalid = |(InputExc[4:2]) ;
	
	// Inexact answer due to rounding, overflow or underflow
	assign Inexact = (R | S) | Overflow | Underflow;
	
	// Put pieces together to form final result
	assign P = Z ;
	
	// Collect exception flags	
	assign Flags = {Overflow, Underflow, DivideByZero, Invalid, Inexact} ; 	
	
endmodule
`endif

