
module dense_latency_ap_fixed_ap_fixed_config14_0_0_0_0_0_0 (
        ap_clk,
        ap_rst,
        data_0_V_read,
        data_1_V_read,
        data_2_V_read,
        data_3_V_read,
        data_4_V_read,
        data_5_V_read,
        data_6_V_read,
        data_7_V_read,
        data_8_V_read,
        data_9_V_read,
        data_10_V_read,
        data_11_V_read,
        data_12_V_read,
        data_13_V_read,
        data_14_V_read,
        data_15_V_read,
        data_16_V_read,
        data_17_V_read,
        data_18_V_read,
        data_19_V_read,
        data_20_V_read,
        data_21_V_read,
        data_22_V_read,
        data_23_V_read,
        data_24_V_read,
        data_25_V_read,
        data_26_V_read,
        data_27_V_read,
        data_28_V_read,
        data_29_V_read,
        data_30_V_read,
        data_31_V_read,
        ap_return_0,
        ap_return_1,
        ap_return_2,
        ap_return_3,
        ap_return_4,
        ap_ce
);


input   ap_clk;
input   ap_rst;
input  [15:0] data_0_V_read;
input  [15:0] data_1_V_read;
input  [15:0] data_2_V_read;
input  [15:0] data_3_V_read;
input  [15:0] data_4_V_read;
input  [15:0] data_5_V_read;
input  [15:0] data_6_V_read;
input  [15:0] data_7_V_read;
input  [15:0] data_8_V_read;
input  [15:0] data_9_V_read;
input  [15:0] data_10_V_read;
input  [15:0] data_11_V_read;
input  [15:0] data_12_V_read;
input  [15:0] data_13_V_read;
input  [15:0] data_14_V_read;
input  [15:0] data_15_V_read;
input  [15:0] data_16_V_read;
input  [15:0] data_17_V_read;
input  [15:0] data_18_V_read;
input  [15:0] data_19_V_read;
input  [15:0] data_20_V_read;
input  [15:0] data_21_V_read;
input  [15:0] data_22_V_read;
input  [15:0] data_23_V_read;
input  [15:0] data_24_V_read;
input  [15:0] data_25_V_read;
input  [15:0] data_26_V_read;
input  [15:0] data_27_V_read;
input  [15:0] data_28_V_read;
input  [15:0] data_29_V_read;
input  [15:0] data_30_V_read;
input  [15:0] data_31_V_read;
output  [15:0] ap_return_0;
output  [15:0] ap_return_1;
output  [15:0] ap_return_2;
output  [15:0] ap_return_3;
output  [15:0] ap_return_4;
input   ap_ce;

reg[15:0] ap_return_0;
reg[15:0] ap_return_1;
reg[15:0] ap_return_2;
reg[15:0] ap_return_3;
reg[15:0] ap_return_4;

reg   [15:0] data_31_V_read32_reg_989;
wire    ap_block_state1_pp0_stage0_iter0;
wire    ap_block_state2_pp0_stage0_iter1;
wire    ap_block_state3_pp0_stage0_iter2;
wire    ap_block_state4_pp0_stage0_iter3;
wire    ap_block_state5_pp0_stage0_iter4;
wire    ap_block_state6_pp0_stage0_iter5;
wire    ap_block_state7_pp0_stage0_iter6;
wire    ap_block_state8_pp0_stage0_iter7;
wire    ap_block_pp0_stage0_11001;
reg   [15:0] data_31_V_read32_reg_989_pp0_iter1_reg;
reg   [15:0] data_31_V_read32_reg_989_pp0_iter2_reg;
reg   [15:0] data_31_V_read32_reg_989_pp0_iter3_reg;
reg   [15:0] data_31_V_read32_reg_989_pp0_iter4_reg;
reg   [15:0] data_31_V_read32_reg_989_pp0_iter5_reg;
reg   [15:0] data_31_V_read32_reg_989_pp0_iter6_reg;
reg   [15:0] data_30_V_read31_reg_998;
reg   [15:0] data_30_V_read31_reg_998_pp0_iter1_reg;
reg   [15:0] data_30_V_read31_reg_998_pp0_iter2_reg;
reg   [15:0] data_30_V_read31_reg_998_pp0_iter3_reg;
reg   [15:0] data_30_V_read31_reg_998_pp0_iter4_reg;
reg   [15:0] data_30_V_read31_reg_998_pp0_iter5_reg;
reg   [15:0] data_30_V_read31_reg_998_pp0_iter6_reg;
reg   [15:0] data_29_V_read_6_reg_1006;
reg   [15:0] data_29_V_read_6_reg_1006_pp0_iter1_reg;
reg   [15:0] data_29_V_read_6_reg_1006_pp0_iter2_reg;
reg   [15:0] data_29_V_read_6_reg_1006_pp0_iter3_reg;
reg   [15:0] data_29_V_read_6_reg_1006_pp0_iter4_reg;
reg   [15:0] data_29_V_read_6_reg_1006_pp0_iter5_reg;
reg   [15:0] data_29_V_read_6_reg_1006_pp0_iter6_reg;
reg   [15:0] data_28_V_read_6_reg_1014;
reg   [15:0] data_28_V_read_6_reg_1014_pp0_iter1_reg;
reg   [15:0] data_28_V_read_6_reg_1014_pp0_iter2_reg;
reg   [15:0] data_28_V_read_6_reg_1014_pp0_iter3_reg;
reg   [15:0] data_28_V_read_6_reg_1014_pp0_iter4_reg;
reg   [15:0] data_28_V_read_6_reg_1014_pp0_iter5_reg;
reg   [15:0] data_28_V_read_6_reg_1014_pp0_iter6_reg;
reg   [15:0] data_27_V_read_7_reg_1023;
reg   [15:0] data_27_V_read_7_reg_1023_pp0_iter1_reg;
reg   [15:0] data_27_V_read_7_reg_1023_pp0_iter2_reg;
reg   [15:0] data_27_V_read_7_reg_1023_pp0_iter3_reg;
reg   [15:0] data_27_V_read_7_reg_1023_pp0_iter4_reg;
reg   [15:0] data_27_V_read_7_reg_1023_pp0_iter5_reg;
reg   [15:0] data_26_V_read_7_reg_1032;
reg   [15:0] data_26_V_read_7_reg_1032_pp0_iter1_reg;
reg   [15:0] data_26_V_read_7_reg_1032_pp0_iter2_reg;
reg   [15:0] data_26_V_read_7_reg_1032_pp0_iter3_reg;
reg   [15:0] data_26_V_read_7_reg_1032_pp0_iter4_reg;
reg   [15:0] data_26_V_read_7_reg_1032_pp0_iter5_reg;
reg   [15:0] data_25_V_read26_reg_1041;
reg   [15:0] data_25_V_read26_reg_1041_pp0_iter1_reg;
reg   [15:0] data_25_V_read26_reg_1041_pp0_iter2_reg;
reg   [15:0] data_25_V_read26_reg_1041_pp0_iter3_reg;
reg   [15:0] data_25_V_read26_reg_1041_pp0_iter4_reg;
reg   [15:0] data_25_V_read26_reg_1041_pp0_iter5_reg;
reg   [15:0] data_24_V_read25_reg_1050;
reg   [15:0] data_24_V_read25_reg_1050_pp0_iter1_reg;
reg   [15:0] data_24_V_read25_reg_1050_pp0_iter2_reg;
reg   [15:0] data_24_V_read25_reg_1050_pp0_iter3_reg;
reg   [15:0] data_24_V_read25_reg_1050_pp0_iter4_reg;
reg   [15:0] data_24_V_read25_reg_1050_pp0_iter5_reg;
reg   [15:0] data_23_V_read24_reg_1059;
reg   [15:0] data_23_V_read24_reg_1059_pp0_iter1_reg;
reg   [15:0] data_23_V_read24_reg_1059_pp0_iter2_reg;
reg   [15:0] data_23_V_read24_reg_1059_pp0_iter3_reg;
reg   [15:0] data_23_V_read24_reg_1059_pp0_iter4_reg;
reg   [15:0] data_22_V_read23_reg_1068;
reg   [15:0] data_22_V_read23_reg_1068_pp0_iter1_reg;
reg   [15:0] data_22_V_read23_reg_1068_pp0_iter2_reg;
reg   [15:0] data_22_V_read23_reg_1068_pp0_iter3_reg;
reg   [15:0] data_22_V_read23_reg_1068_pp0_iter4_reg;
reg   [15:0] data_22_V_read23_reg_1068_pp0_iter5_reg;
reg   [15:0] data_21_V_read22_reg_1077;
reg   [15:0] data_21_V_read22_reg_1077_pp0_iter1_reg;
reg   [15:0] data_21_V_read22_reg_1077_pp0_iter2_reg;
reg   [15:0] data_21_V_read22_reg_1077_pp0_iter3_reg;
reg   [15:0] data_21_V_read22_reg_1077_pp0_iter4_reg;
reg   [15:0] data_20_V_read21_reg_1086;
reg   [15:0] data_20_V_read21_reg_1086_pp0_iter1_reg;
reg   [15:0] data_20_V_read21_reg_1086_pp0_iter2_reg;
reg   [15:0] data_20_V_read21_reg_1086_pp0_iter3_reg;
reg   [15:0] data_20_V_read21_reg_1086_pp0_iter4_reg;
reg   [15:0] data_19_V_read_6_reg_1095;
reg   [15:0] data_19_V_read_6_reg_1095_pp0_iter1_reg;
reg   [15:0] data_19_V_read_6_reg_1095_pp0_iter2_reg;
reg   [15:0] data_19_V_read_6_reg_1095_pp0_iter3_reg;
reg   [15:0] data_19_V_read_6_reg_1095_pp0_iter4_reg;
reg   [15:0] data_18_V_read_6_reg_1103;
reg   [15:0] data_18_V_read_6_reg_1103_pp0_iter1_reg;
reg   [15:0] data_18_V_read_6_reg_1103_pp0_iter2_reg;
reg   [15:0] data_18_V_read_6_reg_1103_pp0_iter3_reg;
reg   [15:0] data_18_V_read_6_reg_1103_pp0_iter4_reg;
reg   [15:0] data_17_V_read_7_reg_1111;
reg   [15:0] data_17_V_read_7_reg_1111_pp0_iter1_reg;
reg   [15:0] data_17_V_read_7_reg_1111_pp0_iter2_reg;
reg   [15:0] data_17_V_read_7_reg_1111_pp0_iter3_reg;
reg   [15:0] data_16_V_read_7_reg_1120;
reg   [15:0] data_16_V_read_7_reg_1120_pp0_iter1_reg;
reg   [15:0] data_16_V_read_7_reg_1120_pp0_iter2_reg;
reg   [15:0] data_16_V_read_7_reg_1120_pp0_iter3_reg;
reg   [15:0] data_15_V_read16_reg_1129;
reg   [15:0] data_15_V_read16_reg_1129_pp0_iter1_reg;
reg   [15:0] data_15_V_read16_reg_1129_pp0_iter2_reg;
reg   [15:0] data_15_V_read16_reg_1129_pp0_iter3_reg;
reg   [15:0] data_14_V_read15_reg_1138;
reg   [15:0] data_14_V_read15_reg_1138_pp0_iter1_reg;
reg   [15:0] data_14_V_read15_reg_1138_pp0_iter2_reg;
reg   [15:0] data_14_V_read15_reg_1138_pp0_iter3_reg;
reg   [15:0] data_13_V_read14_reg_1147;
reg   [15:0] data_13_V_read14_reg_1147_pp0_iter1_reg;
reg   [15:0] data_13_V_read14_reg_1147_pp0_iter2_reg;
reg   [15:0] data_12_V_read13_reg_1156;
reg   [15:0] data_12_V_read13_reg_1156_pp0_iter1_reg;
reg   [15:0] data_12_V_read13_reg_1156_pp0_iter2_reg;
reg   [15:0] data_11_V_read12_reg_1165;
reg   [15:0] data_11_V_read12_reg_1165_pp0_iter1_reg;
reg   [15:0] data_11_V_read12_reg_1165_pp0_iter2_reg;
reg   [15:0] data_10_V_read11_reg_1174;
reg   [15:0] data_10_V_read11_reg_1174_pp0_iter1_reg;
reg   [15:0] data_10_V_read11_reg_1174_pp0_iter2_reg;
reg   [15:0] data_9_V_read_6_reg_1183;
reg   [15:0] data_9_V_read_6_reg_1183_pp0_iter1_reg;
reg   [15:0] data_8_V_read_6_reg_1192;
reg   [15:0] data_8_V_read_6_reg_1192_pp0_iter1_reg;
reg   [15:0] data_7_V_read_7_reg_1201;
reg   [15:0] data_7_V_read_7_reg_1201_pp0_iter1_reg;
reg   [15:0] data_6_V_read_7_reg_1208;
reg   [15:0] data_5_V_read_7_reg_1215;
reg   [15:0] data_5_V_read_7_reg_1215_pp0_iter1_reg;
reg   [15:0] data_4_V_read_8_reg_1224;
reg   [15:0] data_3_V_read_8_reg_1232;
reg   [15:0] data_2_V_read_8_reg_1240;
wire   [15:0] add_ln703_fu_280_p2;
reg   [15:0] add_ln703_reg_1246;
wire   [15:0] sub_ln703_1_fu_286_p2;
reg   [15:0] sub_ln703_1_reg_1252;
wire   [15:0] sub_ln703_5_fu_319_p2;
reg   [15:0] sub_ln703_5_reg_1258;
wire   [15:0] sub_ln703_6_fu_324_p2;
reg   [15:0] sub_ln703_6_reg_1263;
wire   [15:0] add_ln703_136_fu_347_p2;
reg   [15:0] add_ln703_136_reg_1268;
wire   [15:0] sub_ln703_9_fu_353_p2;
reg   [15:0] sub_ln703_9_reg_1273;
wire   [15:0] add_ln703_138_fu_363_p2;
reg   [15:0] add_ln703_138_reg_1278;
wire   [15:0] add_ln703_139_fu_367_p2;
reg   [15:0] add_ln703_139_reg_1284;
wire   [15:0] add_ln703_145_fu_433_p2;
reg   [15:0] add_ln703_145_reg_1289;
wire   [15:0] sub_ln703_18_fu_443_p2;
reg   [15:0] sub_ln703_18_reg_1294;
wire   [15:0] add_ln703_146_fu_453_p2;
reg   [15:0] add_ln703_146_reg_1299;
wire   [15:0] add_ln703_147_fu_458_p2;
reg   [15:0] add_ln703_147_reg_1304;
wire   [15:0] add_ln703_148_fu_463_p2;
reg   [15:0] add_ln703_148_reg_1309;
wire   [15:0] add_ln703_149_fu_468_p2;
reg   [15:0] add_ln703_149_reg_1314;
wire   [15:0] sub_ln703_25_fu_517_p2;
reg   [15:0] sub_ln703_25_reg_1319;
wire   [15:0] sub_ln703_26_fu_527_p2;
reg   [15:0] sub_ln703_26_reg_1324;
wire   [15:0] sub_ln703_28_fu_537_p2;
reg   [15:0] sub_ln703_28_reg_1329;
wire   [15:0] sub_ln703_30_fu_542_p2;
reg   [15:0] sub_ln703_30_reg_1334;
wire   [15:0] sub_ln703_33_fu_562_p2;
reg   [15:0] sub_ln703_33_reg_1339;
wire   [15:0] add_ln703_166_fu_567_p2;
reg   [15:0] add_ln703_166_reg_1344;
wire   [15:0] add_ln703_163_fu_621_p2;
reg   [15:0] add_ln703_163_reg_1350;
wire   [15:0] sub_ln703_38_fu_626_p2;
reg   [15:0] sub_ln703_38_reg_1355;
wire   [15:0] add_ln703_167_fu_641_p2;
reg   [15:0] add_ln703_167_reg_1360;
wire   [15:0] sub_ln703_41_fu_646_p2;
reg   [15:0] sub_ln703_41_reg_1365;
wire   [15:0] add_ln703_176_fu_660_p2;
reg   [15:0] add_ln703_176_reg_1370;
reg   [15:0] add_ln703_176_reg_1370_pp0_iter5_reg;
wire   [15:0] sub_ln703_46_fu_697_p2;
reg   [15:0] sub_ln703_46_reg_1375;
wire   [15:0] add_ln703_173_fu_732_p2;
reg   [15:0] add_ln703_173_reg_1380;
wire   [15:0] sub_ln703_49_fu_737_p2;
reg   [15:0] sub_ln703_49_reg_1385;
wire   [15:0] sub_ln703_50_fu_742_p2;
reg   [15:0] sub_ln703_50_reg_1390;
wire   [15:0] add_ln703_180_fu_760_p2;
reg   [15:0] add_ln703_180_reg_1395;
wire   [15:0] add_ln703_184_fu_770_p2;
reg   [15:0] add_ln703_184_reg_1400;
wire   [15:0] sub_ln703_61_fu_840_p2;
reg   [15:0] sub_ln703_61_reg_1405;
wire   [15:0] add_ln703_189_fu_855_p2;
reg   [15:0] add_ln703_189_reg_1410;
wire   [15:0] sub_ln703_62_fu_860_p2;
reg   [15:0] sub_ln703_62_reg_1415;
wire   [15:0] sub_ln703_64_fu_865_p2;
reg   [15:0] sub_ln703_64_reg_1420;
wire   [15:0] add_ln703_192_fu_870_p2;
reg   [15:0] add_ln703_192_reg_1425;
wire   [15:0] add_ln703_194_fu_874_p2;
reg   [15:0] add_ln703_194_reg_1431;
wire    ap_block_pp0_stage0;
wire   [15:0] sub_ln703_fu_274_p2;
wire   [15:0] add_ln703_130_fu_300_p2;
wire   [15:0] sub_ln703_2_fu_292_p2;
wire   [15:0] sub_ln703_3_fu_296_p2;
wire   [15:0] add_ln703_131_fu_304_p2;
wire   [15:0] sub_ln703_4_fu_309_p2;
wire   [15:0] add_ln703_132_fu_314_p2;
wire   [15:0] add_ln703_134_fu_338_p2;
wire   [15:0] add_ln703_135_fu_342_p2;
wire   [15:0] add_ln703_133_fu_334_p2;
wire   [15:0] sub_ln703_8_fu_329_p2;
wire   [15:0] add_ln703_137_fu_358_p2;
wire   [15:0] sub_ln703_7_fu_373_p2;
wire   [15:0] add_ln703_141_fu_386_p2;
wire   [15:0] sub_ln703_10_fu_377_p2;
wire   [15:0] add_ln703_140_fu_381_p2;
wire   [15:0] add_ln703_142_fu_390_p2;
wire   [15:0] add_ln703_143_fu_395_p2;
wire   [15:0] add_ln703_144_fu_399_p2;
wire   [15:0] sub_ln703_11_fu_404_p2;
wire   [15:0] sub_ln703_13_fu_413_p2;
wire   [15:0] sub_ln703_14_fu_418_p2;
wire   [15:0] sub_ln703_15_fu_423_p2;
wire   [15:0] sub_ln703_16_fu_428_p2;
wire   [15:0] sub_ln703_17_fu_438_p2;
wire   [15:0] sub_ln703_19_fu_448_p2;
wire   [15:0] sub_ln703_12_fu_408_p2;
wire   [15:0] sub_ln703_20_fu_472_p2;
wire   [15:0] add_ln703_151_fu_489_p2;
wire   [15:0] add_ln703_150_fu_476_p2;
wire   [15:0] sub_ln703_21_fu_480_p2;
wire   [15:0] sub_ln703_22_fu_485_p2;
wire   [15:0] add_ln703_152_fu_493_p2;
wire   [15:0] sub_ln703_24_fu_502_p2;
wire   [15:0] add_ln703_153_fu_507_p2;
wire   [15:0] add_ln703_154_fu_512_p2;
wire   [15:0] add_ln703_155_fu_522_p2;
wire   [15:0] sub_ln703_27_fu_532_p2;
wire   [15:0] sub_ln703_23_fu_498_p2;
wire   [15:0] add_ln703_158_fu_552_p2;
wire   [15:0] add_ln703_157_fu_547_p2;
wire   [15:0] add_ln703_159_fu_556_p2;
wire   [15:0] add_ln703_156_fu_571_p2;
wire   [15:0] sub_ln703_29_fu_575_p2;
wire   [15:0] sub_ln703_32_fu_584_p2;
wire   [15:0] add_ln703_160_fu_588_p2;
wire   [15:0] add_ln703_161_fu_593_p2;
wire   [15:0] sub_ln703_34_fu_597_p2;
wire   [15:0] sub_ln703_35_fu_602_p2;
wire   [15:0] add_ln703_162_fu_616_p2;
wire   [15:0] add_ln703_164_fu_631_p2;
wire   [15:0] sub_ln703_36_fu_607_p2;
wire   [15:0] sub_ln703_37_fu_612_p2;
wire   [15:0] add_ln703_165_fu_635_p2;
wire   [15:0] sub_ln703_31_fu_579_p2;
wire   [15:0] add_ln703_175_fu_656_p2;
wire   [15:0] add_ln703_174_fu_651_p2;
wire   [15:0] sub_ln703_39_fu_666_p2;
wire   [15:0] add_ln703_168_fu_674_p2;
wire   [15:0] sub_ln703_42_fu_679_p2;
wire   [15:0] sub_ln703_43_fu_683_p2;
wire   [15:0] sub_ln703_44_fu_688_p2;
wire   [15:0] sub_ln703_45_fu_692_p2;
wire   [15:0] sub_ln703_40_fu_670_p2;
wire   [15:0] add_ln703_171_fu_717_p2;
wire   [15:0] add_ln703_170_fu_712_p2;
wire   [15:0] add_ln703_169_fu_702_p2;
wire   [15:0] sub_ln703_47_fu_707_p2;
wire   [15:0] add_ln703_172_fu_721_p2;
wire   [15:0] sub_ln703_48_fu_727_p2;
wire   [15:0] add_ln703_178_fu_751_p2;
wire   [15:0] add_ln703_179_fu_755_p2;
wire   [15:0] add_ln703_177_fu_747_p2;
wire   [15:0] add_ln703_183_fu_766_p2;
wire   [15:0] add_ln703_181_fu_775_p2;
wire   [15:0] sub_ln703_51_fu_779_p2;
wire   [15:0] sub_ln703_52_fu_783_p2;
wire   [15:0] add_ln703_182_fu_806_p2;
wire   [15:0] sub_ln703_53_fu_787_p2;
wire   [15:0] sub_ln703_54_fu_791_p2;
wire   [15:0] sub_ln703_56_fu_801_p2;
wire   [15:0] add_ln703_185_fu_810_p2;
wire   [15:0] add_ln703_186_fu_815_p2;
wire   [15:0] sub_ln703_57_fu_820_p2;
wire   [15:0] add_ln703_187_fu_845_p2;
wire   [15:0] sub_ln703_55_fu_796_p2;
wire   [15:0] sub_ln703_59_fu_830_p2;
wire   [15:0] sub_ln703_60_fu_835_p2;
wire   [15:0] add_ln703_188_fu_849_p2;
wire   [15:0] sub_ln703_58_fu_825_p2;
wire   [15:0] sub_ln703_63_fu_879_p2;
wire   [15:0] sub_ln703_65_fu_883_p2;
wire   [15:0] add_ln703_190_fu_887_p2;
wire   [15:0] sub_ln703_66_fu_891_p2;
wire   [15:0] add_ln703_195_fu_915_p2;
wire   [15:0] add_ln703_191_fu_896_p2;
wire   [15:0] sub_ln703_68_fu_906_p2;
wire   [15:0] add_ln703_193_fu_911_p2;
wire   [15:0] add_ln703_196_fu_919_p2;
wire   [15:0] sub_ln703_69_fu_924_p2;
wire   [15:0] add_ln703_198_fu_949_p2;
wire   [15:0] sub_ln703_67_fu_901_p2;
wire   [15:0] sub_ln703_70_fu_929_p2;
wire   [15:0] acc_1_V_fu_934_p2;
wire   [15:0] acc_2_V_fu_939_p2;
wire   [15:0] acc_3_V_fu_944_p2;
wire   [15:0] acc_4_V_fu_953_p2;
reg    ap_ce_reg;
reg   [15:0] data_0_V_read_int_reg;
reg   [15:0] data_1_V_read_int_reg;
reg   [15:0] data_2_V_read_int_reg;
reg   [15:0] data_3_V_read_int_reg;
reg   [15:0] data_4_V_read_int_reg;
reg   [15:0] data_5_V_read_int_reg;
reg   [15:0] data_6_V_read_int_reg;
reg   [15:0] data_7_V_read_int_reg;
reg   [15:0] data_8_V_read_int_reg;
reg   [15:0] data_9_V_read_int_reg;
reg   [15:0] data_10_V_read_int_reg;
reg   [15:0] data_11_V_read_int_reg;
reg   [15:0] data_12_V_read_int_reg;
reg   [15:0] data_13_V_read_int_reg;
reg   [15:0] data_14_V_read_int_reg;
reg   [15:0] data_15_V_read_int_reg;
reg   [15:0] data_16_V_read_int_reg;
reg   [15:0] data_17_V_read_int_reg;
reg   [15:0] data_18_V_read_int_reg;
reg   [15:0] data_19_V_read_int_reg;
reg   [15:0] data_20_V_read_int_reg;
reg   [15:0] data_21_V_read_int_reg;
reg   [15:0] data_22_V_read_int_reg;
reg   [15:0] data_23_V_read_int_reg;
reg   [15:0] data_24_V_read_int_reg;
reg   [15:0] data_25_V_read_int_reg;
reg   [15:0] data_26_V_read_int_reg;
reg   [15:0] data_27_V_read_int_reg;
reg   [15:0] data_28_V_read_int_reg;
reg   [15:0] data_29_V_read_int_reg;
reg   [15:0] data_30_V_read_int_reg;
reg   [15:0] data_31_V_read_int_reg;
reg   [15:0] ap_return_0_int_reg;
reg   [15:0] ap_return_1_int_reg;
reg   [15:0] ap_return_2_int_reg;
reg   [15:0] ap_return_3_int_reg;
reg   [15:0] ap_return_4_int_reg;

always @ (posedge ap_clk) begin
    ap_ce_reg <= ap_ce;
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_ce_reg) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        add_ln703_136_reg_1268 <= add_ln703_136_fu_347_p2;
        add_ln703_138_reg_1278 <= add_ln703_138_fu_363_p2;
        add_ln703_139_reg_1284 <= add_ln703_139_fu_367_p2;
        add_ln703_145_reg_1289 <= add_ln703_145_fu_433_p2;
        add_ln703_146_reg_1299 <= add_ln703_146_fu_453_p2;
        add_ln703_147_reg_1304 <= add_ln703_147_fu_458_p2;
        add_ln703_148_reg_1309 <= add_ln703_148_fu_463_p2;
        add_ln703_149_reg_1314 <= add_ln703_149_fu_468_p2;
        add_ln703_163_reg_1350 <= add_ln703_163_fu_621_p2;
        add_ln703_166_reg_1344 <= add_ln703_166_fu_567_p2;
        add_ln703_167_reg_1360 <= add_ln703_167_fu_641_p2;
        add_ln703_173_reg_1380 <= add_ln703_173_fu_732_p2;
        add_ln703_176_reg_1370 <= add_ln703_176_fu_660_p2;
        add_ln703_176_reg_1370_pp0_iter5_reg <= add_ln703_176_reg_1370;
        add_ln703_180_reg_1395 <= add_ln703_180_fu_760_p2;
        add_ln703_184_reg_1400 <= add_ln703_184_fu_770_p2;
        add_ln703_189_reg_1410 <= add_ln703_189_fu_855_p2;
        add_ln703_192_reg_1425 <= add_ln703_192_fu_870_p2;
        add_ln703_194_reg_1431 <= add_ln703_194_fu_874_p2;
        add_ln703_reg_1246 <= add_ln703_fu_280_p2;
        data_10_V_read11_reg_1174 <= data_10_V_read_int_reg;
        data_10_V_read11_reg_1174_pp0_iter1_reg <= data_10_V_read11_reg_1174;
        data_10_V_read11_reg_1174_pp0_iter2_reg <= data_10_V_read11_reg_1174_pp0_iter1_reg;
        data_11_V_read12_reg_1165 <= data_11_V_read_int_reg;
        data_11_V_read12_reg_1165_pp0_iter1_reg <= data_11_V_read12_reg_1165;
        data_11_V_read12_reg_1165_pp0_iter2_reg <= data_11_V_read12_reg_1165_pp0_iter1_reg;
        data_12_V_read13_reg_1156 <= data_12_V_read_int_reg;
        data_12_V_read13_reg_1156_pp0_iter1_reg <= data_12_V_read13_reg_1156;
        data_12_V_read13_reg_1156_pp0_iter2_reg <= data_12_V_read13_reg_1156_pp0_iter1_reg;
        data_13_V_read14_reg_1147 <= data_13_V_read_int_reg;
        data_13_V_read14_reg_1147_pp0_iter1_reg <= data_13_V_read14_reg_1147;
        data_13_V_read14_reg_1147_pp0_iter2_reg <= data_13_V_read14_reg_1147_pp0_iter1_reg;
        data_14_V_read15_reg_1138 <= data_14_V_read_int_reg;
        data_14_V_read15_reg_1138_pp0_iter1_reg <= data_14_V_read15_reg_1138;
        data_14_V_read15_reg_1138_pp0_iter2_reg <= data_14_V_read15_reg_1138_pp0_iter1_reg;
        data_14_V_read15_reg_1138_pp0_iter3_reg <= data_14_V_read15_reg_1138_pp0_iter2_reg;
        data_15_V_read16_reg_1129 <= data_15_V_read_int_reg;
        data_15_V_read16_reg_1129_pp0_iter1_reg <= data_15_V_read16_reg_1129;
        data_15_V_read16_reg_1129_pp0_iter2_reg <= data_15_V_read16_reg_1129_pp0_iter1_reg;
        data_15_V_read16_reg_1129_pp0_iter3_reg <= data_15_V_read16_reg_1129_pp0_iter2_reg;
        data_16_V_read_7_reg_1120 <= data_16_V_read_int_reg;
        data_16_V_read_7_reg_1120_pp0_iter1_reg <= data_16_V_read_7_reg_1120;
        data_16_V_read_7_reg_1120_pp0_iter2_reg <= data_16_V_read_7_reg_1120_pp0_iter1_reg;
        data_16_V_read_7_reg_1120_pp0_iter3_reg <= data_16_V_read_7_reg_1120_pp0_iter2_reg;
        data_17_V_read_7_reg_1111 <= data_17_V_read_int_reg;
        data_17_V_read_7_reg_1111_pp0_iter1_reg <= data_17_V_read_7_reg_1111;
        data_17_V_read_7_reg_1111_pp0_iter2_reg <= data_17_V_read_7_reg_1111_pp0_iter1_reg;
        data_17_V_read_7_reg_1111_pp0_iter3_reg <= data_17_V_read_7_reg_1111_pp0_iter2_reg;
        data_18_V_read_6_reg_1103 <= data_18_V_read_int_reg;
        data_18_V_read_6_reg_1103_pp0_iter1_reg <= data_18_V_read_6_reg_1103;
        data_18_V_read_6_reg_1103_pp0_iter2_reg <= data_18_V_read_6_reg_1103_pp0_iter1_reg;
        data_18_V_read_6_reg_1103_pp0_iter3_reg <= data_18_V_read_6_reg_1103_pp0_iter2_reg;
        data_18_V_read_6_reg_1103_pp0_iter4_reg <= data_18_V_read_6_reg_1103_pp0_iter3_reg;
        data_19_V_read_6_reg_1095 <= data_19_V_read_int_reg;
        data_19_V_read_6_reg_1095_pp0_iter1_reg <= data_19_V_read_6_reg_1095;
        data_19_V_read_6_reg_1095_pp0_iter2_reg <= data_19_V_read_6_reg_1095_pp0_iter1_reg;
        data_19_V_read_6_reg_1095_pp0_iter3_reg <= data_19_V_read_6_reg_1095_pp0_iter2_reg;
        data_19_V_read_6_reg_1095_pp0_iter4_reg <= data_19_V_read_6_reg_1095_pp0_iter3_reg;
        data_20_V_read21_reg_1086 <= data_20_V_read_int_reg;
        data_20_V_read21_reg_1086_pp0_iter1_reg <= data_20_V_read21_reg_1086;
        data_20_V_read21_reg_1086_pp0_iter2_reg <= data_20_V_read21_reg_1086_pp0_iter1_reg;
        data_20_V_read21_reg_1086_pp0_iter3_reg <= data_20_V_read21_reg_1086_pp0_iter2_reg;
        data_20_V_read21_reg_1086_pp0_iter4_reg <= data_20_V_read21_reg_1086_pp0_iter3_reg;
        data_21_V_read22_reg_1077 <= data_21_V_read_int_reg;
        data_21_V_read22_reg_1077_pp0_iter1_reg <= data_21_V_read22_reg_1077;
        data_21_V_read22_reg_1077_pp0_iter2_reg <= data_21_V_read22_reg_1077_pp0_iter1_reg;
        data_21_V_read22_reg_1077_pp0_iter3_reg <= data_21_V_read22_reg_1077_pp0_iter2_reg;
        data_21_V_read22_reg_1077_pp0_iter4_reg <= data_21_V_read22_reg_1077_pp0_iter3_reg;
        data_22_V_read23_reg_1068 <= data_22_V_read_int_reg;
        data_22_V_read23_reg_1068_pp0_iter1_reg <= data_22_V_read23_reg_1068;
        data_22_V_read23_reg_1068_pp0_iter2_reg <= data_22_V_read23_reg_1068_pp0_iter1_reg;
        data_22_V_read23_reg_1068_pp0_iter3_reg <= data_22_V_read23_reg_1068_pp0_iter2_reg;
        data_22_V_read23_reg_1068_pp0_iter4_reg <= data_22_V_read23_reg_1068_pp0_iter3_reg;
        data_22_V_read23_reg_1068_pp0_iter5_reg <= data_22_V_read23_reg_1068_pp0_iter4_reg;
        data_23_V_read24_reg_1059 <= data_23_V_read_int_reg;
        data_23_V_read24_reg_1059_pp0_iter1_reg <= data_23_V_read24_reg_1059;
        data_23_V_read24_reg_1059_pp0_iter2_reg <= data_23_V_read24_reg_1059_pp0_iter1_reg;
        data_23_V_read24_reg_1059_pp0_iter3_reg <= data_23_V_read24_reg_1059_pp0_iter2_reg;
        data_23_V_read24_reg_1059_pp0_iter4_reg <= data_23_V_read24_reg_1059_pp0_iter3_reg;
        data_24_V_read25_reg_1050 <= data_24_V_read_int_reg;
        data_24_V_read25_reg_1050_pp0_iter1_reg <= data_24_V_read25_reg_1050;
        data_24_V_read25_reg_1050_pp0_iter2_reg <= data_24_V_read25_reg_1050_pp0_iter1_reg;
        data_24_V_read25_reg_1050_pp0_iter3_reg <= data_24_V_read25_reg_1050_pp0_iter2_reg;
        data_24_V_read25_reg_1050_pp0_iter4_reg <= data_24_V_read25_reg_1050_pp0_iter3_reg;
        data_24_V_read25_reg_1050_pp0_iter5_reg <= data_24_V_read25_reg_1050_pp0_iter4_reg;
        data_25_V_read26_reg_1041 <= data_25_V_read_int_reg;
        data_25_V_read26_reg_1041_pp0_iter1_reg <= data_25_V_read26_reg_1041;
        data_25_V_read26_reg_1041_pp0_iter2_reg <= data_25_V_read26_reg_1041_pp0_iter1_reg;
        data_25_V_read26_reg_1041_pp0_iter3_reg <= data_25_V_read26_reg_1041_pp0_iter2_reg;
        data_25_V_read26_reg_1041_pp0_iter4_reg <= data_25_V_read26_reg_1041_pp0_iter3_reg;
        data_25_V_read26_reg_1041_pp0_iter5_reg <= data_25_V_read26_reg_1041_pp0_iter4_reg;
        data_26_V_read_7_reg_1032 <= data_26_V_read_int_reg;
        data_26_V_read_7_reg_1032_pp0_iter1_reg <= data_26_V_read_7_reg_1032;
        data_26_V_read_7_reg_1032_pp0_iter2_reg <= data_26_V_read_7_reg_1032_pp0_iter1_reg;
        data_26_V_read_7_reg_1032_pp0_iter3_reg <= data_26_V_read_7_reg_1032_pp0_iter2_reg;
        data_26_V_read_7_reg_1032_pp0_iter4_reg <= data_26_V_read_7_reg_1032_pp0_iter3_reg;
        data_26_V_read_7_reg_1032_pp0_iter5_reg <= data_26_V_read_7_reg_1032_pp0_iter4_reg;
        data_27_V_read_7_reg_1023 <= data_27_V_read_int_reg;
        data_27_V_read_7_reg_1023_pp0_iter1_reg <= data_27_V_read_7_reg_1023;
        data_27_V_read_7_reg_1023_pp0_iter2_reg <= data_27_V_read_7_reg_1023_pp0_iter1_reg;
        data_27_V_read_7_reg_1023_pp0_iter3_reg <= data_27_V_read_7_reg_1023_pp0_iter2_reg;
        data_27_V_read_7_reg_1023_pp0_iter4_reg <= data_27_V_read_7_reg_1023_pp0_iter3_reg;
        data_27_V_read_7_reg_1023_pp0_iter5_reg <= data_27_V_read_7_reg_1023_pp0_iter4_reg;
        data_28_V_read_6_reg_1014 <= data_28_V_read_int_reg;
        data_28_V_read_6_reg_1014_pp0_iter1_reg <= data_28_V_read_6_reg_1014;
        data_28_V_read_6_reg_1014_pp0_iter2_reg <= data_28_V_read_6_reg_1014_pp0_iter1_reg;
        data_28_V_read_6_reg_1014_pp0_iter3_reg <= data_28_V_read_6_reg_1014_pp0_iter2_reg;
        data_28_V_read_6_reg_1014_pp0_iter4_reg <= data_28_V_read_6_reg_1014_pp0_iter3_reg;
        data_28_V_read_6_reg_1014_pp0_iter5_reg <= data_28_V_read_6_reg_1014_pp0_iter4_reg;
        data_28_V_read_6_reg_1014_pp0_iter6_reg <= data_28_V_read_6_reg_1014_pp0_iter5_reg;
        data_29_V_read_6_reg_1006 <= data_29_V_read_int_reg;
        data_29_V_read_6_reg_1006_pp0_iter1_reg <= data_29_V_read_6_reg_1006;
        data_29_V_read_6_reg_1006_pp0_iter2_reg <= data_29_V_read_6_reg_1006_pp0_iter1_reg;
        data_29_V_read_6_reg_1006_pp0_iter3_reg <= data_29_V_read_6_reg_1006_pp0_iter2_reg;
        data_29_V_read_6_reg_1006_pp0_iter4_reg <= data_29_V_read_6_reg_1006_pp0_iter3_reg;
        data_29_V_read_6_reg_1006_pp0_iter5_reg <= data_29_V_read_6_reg_1006_pp0_iter4_reg;
        data_29_V_read_6_reg_1006_pp0_iter6_reg <= data_29_V_read_6_reg_1006_pp0_iter5_reg;
        data_2_V_read_8_reg_1240 <= data_2_V_read_int_reg;
        data_30_V_read31_reg_998 <= data_30_V_read_int_reg;
        data_30_V_read31_reg_998_pp0_iter1_reg <= data_30_V_read31_reg_998;
        data_30_V_read31_reg_998_pp0_iter2_reg <= data_30_V_read31_reg_998_pp0_iter1_reg;
        data_30_V_read31_reg_998_pp0_iter3_reg <= data_30_V_read31_reg_998_pp0_iter2_reg;
        data_30_V_read31_reg_998_pp0_iter4_reg <= data_30_V_read31_reg_998_pp0_iter3_reg;
        data_30_V_read31_reg_998_pp0_iter5_reg <= data_30_V_read31_reg_998_pp0_iter4_reg;
        data_30_V_read31_reg_998_pp0_iter6_reg <= data_30_V_read31_reg_998_pp0_iter5_reg;
        data_31_V_read32_reg_989 <= data_31_V_read_int_reg;
        data_31_V_read32_reg_989_pp0_iter1_reg <= data_31_V_read32_reg_989;
        data_31_V_read32_reg_989_pp0_iter2_reg <= data_31_V_read32_reg_989_pp0_iter1_reg;
        data_31_V_read32_reg_989_pp0_iter3_reg <= data_31_V_read32_reg_989_pp0_iter2_reg;
        data_31_V_read32_reg_989_pp0_iter4_reg <= data_31_V_read32_reg_989_pp0_iter3_reg;
        data_31_V_read32_reg_989_pp0_iter5_reg <= data_31_V_read32_reg_989_pp0_iter4_reg;
        data_31_V_read32_reg_989_pp0_iter6_reg <= data_31_V_read32_reg_989_pp0_iter5_reg;
        data_3_V_read_8_reg_1232 <= data_3_V_read_int_reg;
        data_4_V_read_8_reg_1224 <= data_4_V_read_int_reg;
        data_5_V_read_7_reg_1215 <= data_5_V_read_int_reg;
        data_5_V_read_7_reg_1215_pp0_iter1_reg <= data_5_V_read_7_reg_1215;
        data_6_V_read_7_reg_1208 <= data_6_V_read_int_reg;
        data_7_V_read_7_reg_1201 <= data_7_V_read_int_reg;
        data_7_V_read_7_reg_1201_pp0_iter1_reg <= data_7_V_read_7_reg_1201;
        data_8_V_read_6_reg_1192 <= data_8_V_read_int_reg;
        data_8_V_read_6_reg_1192_pp0_iter1_reg <= data_8_V_read_6_reg_1192;
        data_9_V_read_6_reg_1183 <= data_9_V_read_int_reg;
        data_9_V_read_6_reg_1183_pp0_iter1_reg <= data_9_V_read_6_reg_1183;
        sub_ln703_18_reg_1294 <= sub_ln703_18_fu_443_p2;
        sub_ln703_1_reg_1252 <= sub_ln703_1_fu_286_p2;
        sub_ln703_25_reg_1319 <= sub_ln703_25_fu_517_p2;
        sub_ln703_26_reg_1324 <= sub_ln703_26_fu_527_p2;
        sub_ln703_28_reg_1329 <= sub_ln703_28_fu_537_p2;
        sub_ln703_30_reg_1334 <= sub_ln703_30_fu_542_p2;
        sub_ln703_33_reg_1339 <= sub_ln703_33_fu_562_p2;
        sub_ln703_38_reg_1355 <= sub_ln703_38_fu_626_p2;
        sub_ln703_41_reg_1365 <= sub_ln703_41_fu_646_p2;
        sub_ln703_46_reg_1375 <= sub_ln703_46_fu_697_p2;
        sub_ln703_49_reg_1385 <= sub_ln703_49_fu_737_p2;
        sub_ln703_50_reg_1390 <= sub_ln703_50_fu_742_p2;
        sub_ln703_5_reg_1258 <= sub_ln703_5_fu_319_p2;
        sub_ln703_61_reg_1405 <= sub_ln703_61_fu_840_p2;
        sub_ln703_62_reg_1415 <= sub_ln703_62_fu_860_p2;
        sub_ln703_64_reg_1420 <= sub_ln703_64_fu_865_p2;
        sub_ln703_6_reg_1263 <= sub_ln703_6_fu_324_p2;
        sub_ln703_9_reg_1273 <= sub_ln703_9_fu_353_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_ce_reg)) begin
        ap_return_0_int_reg <= sub_ln703_70_fu_929_p2;
        ap_return_1_int_reg <= acc_1_V_fu_934_p2;
        ap_return_2_int_reg <= acc_2_V_fu_939_p2;
        ap_return_3_int_reg <= acc_3_V_fu_944_p2;
        ap_return_4_int_reg <= acc_4_V_fu_953_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_ce)) begin
        data_0_V_read_int_reg <= data_0_V_read;
        data_10_V_read_int_reg <= data_10_V_read;
        data_11_V_read_int_reg <= data_11_V_read;
        data_12_V_read_int_reg <= data_12_V_read;
        data_13_V_read_int_reg <= data_13_V_read;
        data_14_V_read_int_reg <= data_14_V_read;
        data_15_V_read_int_reg <= data_15_V_read;
        data_16_V_read_int_reg <= data_16_V_read;
        data_17_V_read_int_reg <= data_17_V_read;
        data_18_V_read_int_reg <= data_18_V_read;
        data_19_V_read_int_reg <= data_19_V_read;
        data_1_V_read_int_reg <= data_1_V_read;
        data_20_V_read_int_reg <= data_20_V_read;
        data_21_V_read_int_reg <= data_21_V_read;
        data_22_V_read_int_reg <= data_22_V_read;
        data_23_V_read_int_reg <= data_23_V_read;
        data_24_V_read_int_reg <= data_24_V_read;
        data_25_V_read_int_reg <= data_25_V_read;
        data_26_V_read_int_reg <= data_26_V_read;
        data_27_V_read_int_reg <= data_27_V_read;
        data_28_V_read_int_reg <= data_28_V_read;
        data_29_V_read_int_reg <= data_29_V_read;
        data_2_V_read_int_reg <= data_2_V_read;
        data_30_V_read_int_reg <= data_30_V_read;
        data_31_V_read_int_reg <= data_31_V_read;
        data_3_V_read_int_reg <= data_3_V_read;
        data_4_V_read_int_reg <= data_4_V_read;
        data_5_V_read_int_reg <= data_5_V_read;
        data_6_V_read_int_reg <= data_6_V_read;
        data_7_V_read_int_reg <= data_7_V_read;
        data_8_V_read_int_reg <= data_8_V_read;
        data_9_V_read_int_reg <= data_9_V_read;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_0 = ap_return_0_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_0 = sub_ln703_70_fu_929_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_1 = ap_return_1_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_1 = acc_1_V_fu_934_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_2 = ap_return_2_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_2 = acc_2_V_fu_939_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_3 = ap_return_3_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_3 = acc_3_V_fu_944_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_4 = ap_return_4_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_4 = acc_4_V_fu_953_p2;
    end
end

assign acc_1_V_fu_934_p2 = (add_ln703_193_fu_911_p2 - data_31_V_read32_reg_989_pp0_iter6_reg);

assign acc_2_V_fu_939_p2 = (add_ln703_196_fu_919_p2 - data_31_V_read32_reg_989_pp0_iter6_reg);

assign acc_3_V_fu_944_p2 = (sub_ln703_69_fu_924_p2 + data_31_V_read32_reg_989_pp0_iter6_reg);

assign acc_4_V_fu_953_p2 = (add_ln703_198_fu_949_p2 + sub_ln703_67_fu_901_p2);

assign add_ln703_130_fu_300_p2 = (data_2_V_read_8_reg_1240 + data_3_V_read_8_reg_1232);

assign add_ln703_131_fu_304_p2 = (add_ln703_130_fu_300_p2 + add_ln703_reg_1246);

assign add_ln703_132_fu_314_p2 = (sub_ln703_3_fu_296_p2 + data_4_V_read_8_reg_1224);

assign add_ln703_133_fu_334_p2 = (sub_ln703_1_reg_1252 + data_3_V_read_8_reg_1232);

assign add_ln703_134_fu_338_p2 = (data_5_V_read_7_reg_1215 + data_6_V_read_7_reg_1208);

assign add_ln703_135_fu_342_p2 = (add_ln703_134_fu_338_p2 + data_4_V_read_8_reg_1224);

assign add_ln703_136_fu_347_p2 = (add_ln703_135_fu_342_p2 + add_ln703_133_fu_334_p2);

assign add_ln703_137_fu_358_p2 = (add_ln703_132_fu_314_p2 + data_5_V_read_7_reg_1215);

assign add_ln703_138_fu_363_p2 = (data_6_V_read_7_reg_1208 + data_7_V_read_7_reg_1201);

assign add_ln703_139_fu_367_p2 = (add_ln703_138_fu_363_p2 + add_ln703_137_fu_358_p2);

assign add_ln703_140_fu_381_p2 = (add_ln703_138_reg_1278 + sub_ln703_7_fu_373_p2);

assign add_ln703_141_fu_386_p2 = (sub_ln703_6_reg_1263 + data_5_V_read_7_reg_1215_pp0_iter1_reg);

assign add_ln703_142_fu_390_p2 = (add_ln703_138_reg_1278 + add_ln703_141_fu_386_p2);

assign add_ln703_143_fu_395_p2 = (sub_ln703_9_reg_1273 + data_7_V_read_7_reg_1201_pp0_iter1_reg);

assign add_ln703_144_fu_399_p2 = (sub_ln703_10_fu_377_p2 + data_8_V_read_6_reg_1192_pp0_iter1_reg);

assign add_ln703_145_fu_433_p2 = (sub_ln703_13_fu_413_p2 + data_9_V_read_6_reg_1183_pp0_iter1_reg);

assign add_ln703_146_fu_453_p2 = (sub_ln703_17_fu_438_p2 + data_10_V_read11_reg_1174_pp0_iter1_reg);

assign add_ln703_147_fu_458_p2 = (sub_ln703_19_fu_448_p2 + data_11_V_read12_reg_1165_pp0_iter1_reg);

assign add_ln703_148_fu_463_p2 = (sub_ln703_12_fu_408_p2 + data_9_V_read_6_reg_1183_pp0_iter1_reg);

assign add_ln703_149_fu_468_p2 = (data_10_V_read11_reg_1174_pp0_iter1_reg + data_11_V_read12_reg_1165_pp0_iter1_reg);

assign add_ln703_150_fu_476_p2 = (add_ln703_149_reg_1314 + add_ln703_148_reg_1309);

assign add_ln703_151_fu_489_p2 = (data_11_V_read12_reg_1165_pp0_iter2_reg + data_12_V_read13_reg_1156_pp0_iter2_reg);

assign add_ln703_152_fu_493_p2 = (add_ln703_151_fu_489_p2 + sub_ln703_18_reg_1294);

assign add_ln703_153_fu_507_p2 = (sub_ln703_21_fu_480_p2 + data_12_V_read13_reg_1156_pp0_iter2_reg);

assign add_ln703_154_fu_512_p2 = (sub_ln703_22_fu_485_p2 + data_12_V_read13_reg_1156_pp0_iter2_reg);

assign add_ln703_155_fu_522_p2 = (sub_ln703_24_fu_502_p2 + data_13_V_read14_reg_1147_pp0_iter2_reg);

assign add_ln703_156_fu_571_p2 = (sub_ln703_25_reg_1319 + data_14_V_read15_reg_1138_pp0_iter3_reg);

assign add_ln703_157_fu_547_p2 = (sub_ln703_23_fu_498_p2 + data_13_V_read14_reg_1147_pp0_iter2_reg);

assign add_ln703_158_fu_552_p2 = (data_14_V_read15_reg_1138_pp0_iter2_reg + data_15_V_read16_reg_1129_pp0_iter2_reg);

assign add_ln703_159_fu_556_p2 = (add_ln703_158_fu_552_p2 + add_ln703_157_fu_547_p2);

assign add_ln703_160_fu_588_p2 = (sub_ln703_29_fu_575_p2 + data_15_V_read16_reg_1129_pp0_iter3_reg);

assign add_ln703_161_fu_593_p2 = (sub_ln703_30_reg_1334 + data_15_V_read16_reg_1129_pp0_iter3_reg);

assign add_ln703_162_fu_616_p2 = (sub_ln703_34_fu_597_p2 + data_17_V_read_7_reg_1111_pp0_iter3_reg);

assign add_ln703_163_fu_621_p2 = (sub_ln703_35_fu_602_p2 + data_17_V_read_7_reg_1111_pp0_iter3_reg);

assign add_ln703_164_fu_631_p2 = (data_17_V_read_7_reg_1111_pp0_iter3_reg + data_18_V_read_6_reg_1103_pp0_iter3_reg);

assign add_ln703_165_fu_635_p2 = (add_ln703_164_fu_631_p2 + sub_ln703_36_fu_607_p2);

assign add_ln703_166_fu_567_p2 = (data_18_V_read_6_reg_1103_pp0_iter2_reg + data_19_V_read_6_reg_1095_pp0_iter2_reg);

assign add_ln703_167_fu_641_p2 = (add_ln703_166_reg_1344 + sub_ln703_37_fu_612_p2);

assign add_ln703_168_fu_674_p2 = (sub_ln703_39_fu_666_p2 + data_19_V_read_6_reg_1095_pp0_iter4_reg);

assign add_ln703_169_fu_702_p2 = (sub_ln703_44_fu_688_p2 + data_21_V_read22_reg_1077_pp0_iter4_reg);

assign add_ln703_170_fu_712_p2 = (sub_ln703_40_fu_670_p2 + data_20_V_read21_reg_1086_pp0_iter4_reg);

assign add_ln703_171_fu_717_p2 = (data_21_V_read22_reg_1077_pp0_iter4_reg + data_22_V_read23_reg_1068_pp0_iter4_reg);

assign add_ln703_172_fu_721_p2 = (add_ln703_171_fu_717_p2 + add_ln703_170_fu_712_p2);

assign add_ln703_173_fu_732_p2 = (sub_ln703_47_fu_707_p2 + data_23_V_read24_reg_1059_pp0_iter4_reg);

assign add_ln703_174_fu_651_p2 = (sub_ln703_31_fu_579_p2 + data_16_V_read_7_reg_1120_pp0_iter3_reg);

assign add_ln703_175_fu_656_p2 = (add_ln703_166_reg_1344 + data_17_V_read_7_reg_1111_pp0_iter3_reg);

assign add_ln703_176_fu_660_p2 = (add_ln703_175_fu_656_p2 + add_ln703_174_fu_651_p2);

assign add_ln703_177_fu_747_p2 = (data_20_V_read21_reg_1086_pp0_iter4_reg + data_21_V_read22_reg_1077_pp0_iter4_reg);

assign add_ln703_178_fu_751_p2 = (data_23_V_read24_reg_1059_pp0_iter4_reg + data_24_V_read25_reg_1050_pp0_iter4_reg);

assign add_ln703_179_fu_755_p2 = (add_ln703_178_fu_751_p2 + data_22_V_read23_reg_1068_pp0_iter4_reg);

assign add_ln703_180_fu_760_p2 = (add_ln703_179_fu_755_p2 + add_ln703_177_fu_747_p2);

assign add_ln703_181_fu_775_p2 = (add_ln703_180_reg_1395 + add_ln703_176_reg_1370_pp0_iter5_reg);

assign add_ln703_182_fu_806_p2 = (sub_ln703_46_reg_1375 + data_22_V_read23_reg_1068_pp0_iter5_reg);

assign add_ln703_183_fu_766_p2 = (data_24_V_read25_reg_1050_pp0_iter4_reg + data_25_V_read26_reg_1041_pp0_iter4_reg);

assign add_ln703_184_fu_770_p2 = (add_ln703_183_fu_766_p2 + data_23_V_read24_reg_1059_pp0_iter4_reg);

assign add_ln703_185_fu_810_p2 = (add_ln703_184_reg_1400 + add_ln703_182_fu_806_p2);

assign add_ln703_186_fu_815_p2 = (sub_ln703_53_fu_787_p2 + data_25_V_read26_reg_1041_pp0_iter5_reg);

assign add_ln703_187_fu_845_p2 = (data_26_V_read_7_reg_1032_pp0_iter5_reg + data_27_V_read_7_reg_1023_pp0_iter5_reg);

assign add_ln703_188_fu_849_p2 = (add_ln703_187_fu_845_p2 + sub_ln703_55_fu_796_p2);

assign add_ln703_189_fu_855_p2 = (sub_ln703_59_fu_830_p2 + data_27_V_read_7_reg_1023_pp0_iter5_reg);

assign add_ln703_190_fu_887_p2 = (sub_ln703_62_reg_1415 + data_28_V_read_6_reg_1014_pp0_iter6_reg);

assign add_ln703_191_fu_896_p2 = (sub_ln703_65_fu_883_p2 + data_29_V_read_6_reg_1006_pp0_iter6_reg);

assign add_ln703_192_fu_870_p2 = (data_29_V_read_6_reg_1006_pp0_iter5_reg + data_30_V_read31_reg_998_pp0_iter5_reg);

assign add_ln703_193_fu_911_p2 = (add_ln703_192_reg_1425 + sub_ln703_64_reg_1420);

assign add_ln703_194_fu_874_p2 = (sub_ln703_58_fu_825_p2 + data_27_V_read_7_reg_1023_pp0_iter5_reg);

assign add_ln703_195_fu_915_p2 = (add_ln703_192_reg_1425 + data_28_V_read_6_reg_1014_pp0_iter6_reg);

assign add_ln703_196_fu_919_p2 = (add_ln703_195_fu_915_p2 + add_ln703_194_reg_1431);

assign add_ln703_198_fu_949_p2 = (data_30_V_read31_reg_998_pp0_iter6_reg + data_31_V_read32_reg_989_pp0_iter6_reg);

assign add_ln703_fu_280_p2 = (data_0_V_read_int_reg + data_1_V_read_int_reg);

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_state1_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter4 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter5 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage0_iter6 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage0_iter7 = ~(1'b1 == 1'b1);

assign sub_ln703_10_fu_377_p2 = (add_ln703_136_reg_1268 - data_7_V_read_7_reg_1201_pp0_iter1_reg);

assign sub_ln703_11_fu_404_p2 = (add_ln703_139_reg_1284 - data_8_V_read_6_reg_1192_pp0_iter1_reg);

assign sub_ln703_12_fu_408_p2 = (add_ln703_140_fu_381_p2 - data_8_V_read_6_reg_1192_pp0_iter1_reg);

assign sub_ln703_13_fu_413_p2 = (add_ln703_142_fu_390_p2 - data_8_V_read_6_reg_1192_pp0_iter1_reg);

assign sub_ln703_14_fu_418_p2 = (add_ln703_143_fu_395_p2 - data_8_V_read_6_reg_1192_pp0_iter1_reg);

assign sub_ln703_15_fu_423_p2 = (add_ln703_144_fu_399_p2 - data_9_V_read_6_reg_1183_pp0_iter1_reg);

assign sub_ln703_16_fu_428_p2 = (sub_ln703_11_fu_404_p2 - data_9_V_read_6_reg_1183_pp0_iter1_reg);

assign sub_ln703_17_fu_438_p2 = (sub_ln703_14_fu_418_p2 - data_9_V_read_6_reg_1183_pp0_iter1_reg);

assign sub_ln703_18_fu_443_p2 = (sub_ln703_15_fu_423_p2 - data_10_V_read11_reg_1174_pp0_iter1_reg);

assign sub_ln703_19_fu_448_p2 = (sub_ln703_16_fu_428_p2 - data_10_V_read11_reg_1174_pp0_iter1_reg);

assign sub_ln703_1_fu_286_p2 = (sub_ln703_fu_274_p2 - data_2_V_read_int_reg);

assign sub_ln703_20_fu_472_p2 = (add_ln703_145_reg_1289 - data_10_V_read11_reg_1174_pp0_iter2_reg);

assign sub_ln703_21_fu_480_p2 = (sub_ln703_20_fu_472_p2 - data_11_V_read12_reg_1165_pp0_iter2_reg);

assign sub_ln703_22_fu_485_p2 = (add_ln703_146_reg_1299 - data_11_V_read12_reg_1165_pp0_iter2_reg);

assign sub_ln703_23_fu_498_p2 = (add_ln703_147_reg_1304 - data_12_V_read13_reg_1156_pp0_iter2_reg);

assign sub_ln703_24_fu_502_p2 = (add_ln703_150_fu_476_p2 - data_12_V_read13_reg_1156_pp0_iter2_reg);

assign sub_ln703_25_fu_517_p2 = (add_ln703_152_fu_493_p2 - data_13_V_read14_reg_1147_pp0_iter2_reg);

assign sub_ln703_26_fu_527_p2 = (add_ln703_153_fu_507_p2 - data_13_V_read14_reg_1147_pp0_iter2_reg);

assign sub_ln703_27_fu_532_p2 = (add_ln703_154_fu_512_p2 - data_13_V_read14_reg_1147_pp0_iter2_reg);

assign sub_ln703_28_fu_537_p2 = (add_ln703_155_fu_522_p2 - data_14_V_read15_reg_1138_pp0_iter2_reg);

assign sub_ln703_29_fu_575_p2 = (sub_ln703_26_reg_1324 - data_14_V_read15_reg_1138_pp0_iter3_reg);

assign sub_ln703_2_fu_292_p2 = (data_2_V_read_8_reg_1240 - add_ln703_reg_1246);

assign sub_ln703_30_fu_542_p2 = (sub_ln703_27_fu_532_p2 - data_14_V_read15_reg_1138_pp0_iter2_reg);

assign sub_ln703_31_fu_579_p2 = (add_ln703_156_fu_571_p2 - data_15_V_read16_reg_1129_pp0_iter3_reg);

assign sub_ln703_32_fu_584_p2 = (sub_ln703_28_reg_1329 - data_15_V_read16_reg_1129_pp0_iter3_reg);

assign sub_ln703_33_fu_562_p2 = (add_ln703_159_fu_556_p2 - data_16_V_read_7_reg_1120_pp0_iter2_reg);

assign sub_ln703_34_fu_597_p2 = (sub_ln703_32_fu_584_p2 - data_16_V_read_7_reg_1120_pp0_iter3_reg);

assign sub_ln703_35_fu_602_p2 = (add_ln703_160_fu_588_p2 - data_16_V_read_7_reg_1120_pp0_iter3_reg);

assign sub_ln703_36_fu_607_p2 = (add_ln703_161_fu_593_p2 - data_16_V_read_7_reg_1120_pp0_iter3_reg);

assign sub_ln703_37_fu_612_p2 = (sub_ln703_33_reg_1339 - data_17_V_read_7_reg_1111_pp0_iter3_reg);

assign sub_ln703_38_fu_626_p2 = (add_ln703_162_fu_616_p2 - data_18_V_read_6_reg_1103_pp0_iter3_reg);

assign sub_ln703_39_fu_666_p2 = (add_ln703_163_reg_1350 - data_18_V_read_6_reg_1103_pp0_iter4_reg);

assign sub_ln703_3_fu_296_p2 = (sub_ln703_1_reg_1252 - data_3_V_read_8_reg_1232);

assign sub_ln703_40_fu_670_p2 = (sub_ln703_38_reg_1355 - data_19_V_read_6_reg_1095_pp0_iter4_reg);

assign sub_ln703_41_fu_646_p2 = (add_ln703_165_fu_635_p2 - data_19_V_read_6_reg_1095_pp0_iter3_reg);

assign sub_ln703_42_fu_679_p2 = (add_ln703_167_reg_1360 - data_20_V_read21_reg_1086_pp0_iter4_reg);

assign sub_ln703_43_fu_683_p2 = (add_ln703_168_fu_674_p2 - data_20_V_read21_reg_1086_pp0_iter4_reg);

assign sub_ln703_44_fu_688_p2 = (sub_ln703_41_reg_1365 - data_20_V_read21_reg_1086_pp0_iter4_reg);

assign sub_ln703_45_fu_692_p2 = (sub_ln703_42_fu_679_p2 - data_21_V_read22_reg_1077_pp0_iter4_reg);

assign sub_ln703_46_fu_697_p2 = (sub_ln703_43_fu_683_p2 - data_21_V_read22_reg_1077_pp0_iter4_reg);

assign sub_ln703_47_fu_707_p2 = (sub_ln703_45_fu_692_p2 - data_22_V_read23_reg_1068_pp0_iter4_reg);

assign sub_ln703_48_fu_727_p2 = (add_ln703_169_fu_702_p2 - data_22_V_read23_reg_1068_pp0_iter4_reg);

assign sub_ln703_49_fu_737_p2 = (add_ln703_172_fu_721_p2 - data_23_V_read24_reg_1059_pp0_iter4_reg);

assign sub_ln703_4_fu_309_p2 = (sub_ln703_2_fu_292_p2 - data_3_V_read_8_reg_1232);

assign sub_ln703_50_fu_742_p2 = (sub_ln703_48_fu_727_p2 - data_23_V_read24_reg_1059_pp0_iter4_reg);

assign sub_ln703_51_fu_779_p2 = (add_ln703_173_reg_1380 - data_24_V_read25_reg_1050_pp0_iter5_reg);

assign sub_ln703_52_fu_783_p2 = (sub_ln703_49_reg_1385 - data_24_V_read25_reg_1050_pp0_iter5_reg);

assign sub_ln703_53_fu_787_p2 = (sub_ln703_50_reg_1390 - data_24_V_read25_reg_1050_pp0_iter5_reg);

assign sub_ln703_54_fu_791_p2 = (add_ln703_181_fu_775_p2 - data_25_V_read26_reg_1041_pp0_iter5_reg);

assign sub_ln703_55_fu_796_p2 = (sub_ln703_51_fu_779_p2 - data_25_V_read26_reg_1041_pp0_iter5_reg);

assign sub_ln703_56_fu_801_p2 = (sub_ln703_52_fu_783_p2 - data_25_V_read26_reg_1041_pp0_iter5_reg);

assign sub_ln703_57_fu_820_p2 = (sub_ln703_54_fu_791_p2 - data_26_V_read_7_reg_1032_pp0_iter5_reg);

assign sub_ln703_58_fu_825_p2 = (sub_ln703_56_fu_801_p2 - data_26_V_read_7_reg_1032_pp0_iter5_reg);

assign sub_ln703_59_fu_830_p2 = (add_ln703_185_fu_810_p2 - data_26_V_read_7_reg_1032_pp0_iter5_reg);

assign sub_ln703_5_fu_319_p2 = (add_ln703_131_fu_304_p2 - data_4_V_read_8_reg_1224);

assign sub_ln703_60_fu_835_p2 = (add_ln703_186_fu_815_p2 - data_26_V_read_7_reg_1032_pp0_iter5_reg);

assign sub_ln703_61_fu_840_p2 = (sub_ln703_57_fu_820_p2 - data_27_V_read_7_reg_1023_pp0_iter5_reg);

assign sub_ln703_62_fu_860_p2 = (sub_ln703_60_fu_835_p2 - data_27_V_read_7_reg_1023_pp0_iter5_reg);

assign sub_ln703_63_fu_879_p2 = (sub_ln703_61_reg_1405 - data_28_V_read_6_reg_1014_pp0_iter6_reg);

assign sub_ln703_64_fu_865_p2 = (add_ln703_188_fu_849_p2 - data_28_V_read_6_reg_1014_pp0_iter5_reg);

assign sub_ln703_65_fu_883_p2 = (add_ln703_189_reg_1410 - data_28_V_read_6_reg_1014_pp0_iter6_reg);

assign sub_ln703_66_fu_891_p2 = (sub_ln703_63_fu_879_p2 - data_29_V_read_6_reg_1006_pp0_iter6_reg);

assign sub_ln703_67_fu_901_p2 = (add_ln703_190_fu_887_p2 - data_29_V_read_6_reg_1006_pp0_iter6_reg);

assign sub_ln703_68_fu_906_p2 = (sub_ln703_66_fu_891_p2 - data_30_V_read31_reg_998_pp0_iter6_reg);

assign sub_ln703_69_fu_924_p2 = (add_ln703_191_fu_896_p2 - data_30_V_read31_reg_998_pp0_iter6_reg);

assign sub_ln703_6_fu_324_p2 = (sub_ln703_4_fu_309_p2 - data_4_V_read_8_reg_1224);

assign sub_ln703_70_fu_929_p2 = (sub_ln703_68_fu_906_p2 - data_31_V_read32_reg_989_pp0_iter6_reg);

assign sub_ln703_7_fu_373_p2 = (sub_ln703_5_reg_1258 - data_5_V_read_7_reg_1215_pp0_iter1_reg);

assign sub_ln703_8_fu_329_p2 = (add_ln703_132_fu_314_p2 - data_5_V_read_7_reg_1215);

assign sub_ln703_9_fu_353_p2 = (sub_ln703_8_fu_329_p2 - data_6_V_read_7_reg_1208);

assign sub_ln703_fu_274_p2 = (data_0_V_read_int_reg - data_1_V_read_int_reg);

endmodule //dense_latency_ap_fixed_ap_fixed_config14_0_0_0_0_0_0
