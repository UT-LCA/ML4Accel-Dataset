
module dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1 (
        ap_clk,
        ap_rst,
        data_V_read,
        ap_return_0,
        ap_return_1,
        ap_return_2,
        ap_return_3,
        ap_return_4,
        ap_return_5,
        ap_return_6,
        ap_return_7,
        ap_return_8,
        ap_return_9,
        ap_return_10,
        ap_return_11,
        ap_return_12,
        ap_return_13,
        ap_return_14,
        ap_return_15,
        ap_return_16,
        ap_return_17,
        ap_return_18,
        ap_return_19,
        ap_return_20,
        ap_return_21,
        ap_return_22,
        ap_return_23,
        ap_return_24,
        ap_return_25,
        ap_return_26,
        ap_return_27,
        ap_return_28,
        ap_return_29,
        ap_return_30,
        ap_return_31,
        ap_return_32,
        ap_return_33,
        ap_return_34,
        ap_return_35,
        ap_return_36,
        ap_return_37,
        ap_return_38,
        ap_return_39,
        ap_return_40,
        ap_return_41,
        ap_return_42,
        ap_return_43,
        ap_return_44,
        ap_return_45,
        ap_return_46,
        ap_return_47,
        ap_return_48,
        ap_return_49,
        ap_return_50,
        ap_return_51,
        ap_return_52,
        ap_return_53,
        ap_return_54,
        ap_return_55,
        ap_return_56,
        ap_return_57,
        ap_return_58,
        ap_return_59,
        ap_return_60,
        ap_return_61,
        ap_return_62,
        ap_return_63,
        ap_ce
);


input   ap_clk;
input   ap_rst;
input  [255:0] data_V_read;
output  [15:0] ap_return_0;
output  [15:0] ap_return_1;
output  [15:0] ap_return_2;
output  [15:0] ap_return_3;
output  [15:0] ap_return_4;
output  [15:0] ap_return_5;
output  [15:0] ap_return_6;
output  [15:0] ap_return_7;
output  [15:0] ap_return_8;
output  [15:0] ap_return_9;
output  [15:0] ap_return_10;
output  [15:0] ap_return_11;
output  [15:0] ap_return_12;
output  [15:0] ap_return_13;
output  [15:0] ap_return_14;
output  [15:0] ap_return_15;
output  [15:0] ap_return_16;
output  [15:0] ap_return_17;
output  [15:0] ap_return_18;
output  [15:0] ap_return_19;
output  [15:0] ap_return_20;
output  [15:0] ap_return_21;
output  [15:0] ap_return_22;
output  [15:0] ap_return_23;
output  [15:0] ap_return_24;
output  [15:0] ap_return_25;
output  [15:0] ap_return_26;
output  [15:0] ap_return_27;
output  [15:0] ap_return_28;
output  [15:0] ap_return_29;
output  [15:0] ap_return_30;
output  [15:0] ap_return_31;
output  [15:0] ap_return_32;
output  [15:0] ap_return_33;
output  [15:0] ap_return_34;
output  [15:0] ap_return_35;
output  [15:0] ap_return_36;
output  [15:0] ap_return_37;
output  [15:0] ap_return_38;
output  [15:0] ap_return_39;
output  [15:0] ap_return_40;
output  [15:0] ap_return_41;
output  [15:0] ap_return_42;
output  [15:0] ap_return_43;
output  [15:0] ap_return_44;
output  [15:0] ap_return_45;
output  [15:0] ap_return_46;
output  [15:0] ap_return_47;
output  [15:0] ap_return_48;
output  [15:0] ap_return_49;
output  [15:0] ap_return_50;
output  [15:0] ap_return_51;
output  [15:0] ap_return_52;
output  [15:0] ap_return_53;
output  [15:0] ap_return_54;
output  [15:0] ap_return_55;
output  [15:0] ap_return_56;
output  [15:0] ap_return_57;
output  [15:0] ap_return_58;
output  [15:0] ap_return_59;
output  [15:0] ap_return_60;
output  [15:0] ap_return_61;
output  [15:0] ap_return_62;
output  [15:0] ap_return_63;
input   ap_ce;

reg[15:0] ap_return_0;
reg[15:0] ap_return_1;
reg[15:0] ap_return_2;
reg[15:0] ap_return_3;
reg[15:0] ap_return_4;
reg[15:0] ap_return_5;
reg[15:0] ap_return_6;
reg[15:0] ap_return_7;
reg[15:0] ap_return_8;
reg[15:0] ap_return_9;
reg[15:0] ap_return_10;
reg[15:0] ap_return_11;
reg[15:0] ap_return_12;
reg[15:0] ap_return_13;
reg[15:0] ap_return_14;
reg[15:0] ap_return_15;
reg[15:0] ap_return_16;
reg[15:0] ap_return_17;
reg[15:0] ap_return_18;
reg[15:0] ap_return_19;
reg[15:0] ap_return_20;
reg[15:0] ap_return_21;
reg[15:0] ap_return_22;
reg[15:0] ap_return_23;
reg[15:0] ap_return_24;
reg[15:0] ap_return_25;
reg[15:0] ap_return_26;
reg[15:0] ap_return_27;
reg[15:0] ap_return_28;
reg[15:0] ap_return_29;
reg[15:0] ap_return_30;
reg[15:0] ap_return_31;
reg[15:0] ap_return_32;
reg[15:0] ap_return_33;
reg[15:0] ap_return_34;
reg[15:0] ap_return_35;
reg[15:0] ap_return_36;
reg[15:0] ap_return_37;
reg[15:0] ap_return_38;
reg[15:0] ap_return_39;
reg[15:0] ap_return_40;
reg[15:0] ap_return_41;
reg[15:0] ap_return_42;
reg[15:0] ap_return_43;
reg[15:0] ap_return_44;
reg[15:0] ap_return_45;
reg[15:0] ap_return_46;
reg[15:0] ap_return_47;
reg[15:0] ap_return_48;
reg[15:0] ap_return_49;
reg[15:0] ap_return_50;
reg[15:0] ap_return_51;
reg[15:0] ap_return_52;
reg[15:0] ap_return_53;
reg[15:0] ap_return_54;
reg[15:0] ap_return_55;
reg[15:0] ap_return_56;
reg[15:0] ap_return_57;
reg[15:0] ap_return_58;
reg[15:0] ap_return_59;
reg[15:0] ap_return_60;
reg[15:0] ap_return_61;
reg[15:0] ap_return_62;
reg[15:0] ap_return_63;

wire   [15:0] trunc_ln203_fu_88_p1;
reg   [15:0] trunc_ln203_reg_3431;
wire    ap_block_state1_pp0_stage0_iter0;
wire    ap_block_state2_pp0_stage0_iter1;
wire    ap_block_state3_pp0_stage0_iter2;
wire    ap_block_state4_pp0_stage0_iter3;
wire    ap_block_state5_pp0_stage0_iter4;
wire    ap_block_state6_pp0_stage0_iter5;
wire    ap_block_state7_pp0_stage0_iter6;
wire    ap_block_state8_pp0_stage0_iter7;
wire    ap_block_state9_pp0_stage0_iter8;
wire    ap_block_pp0_stage0_11001;
wire   [15:0] tmp_2_fu_92_p4;
reg   [15:0] tmp_2_reg_3437;
reg   [15:0] tmp_3_reg_3443;
reg   [15:0] tmp_3_reg_3443_pp0_iter1_reg;
reg   [15:0] tmp_3_reg_3443_pp0_iter2_reg;
reg   [15:0] tmp_4_reg_3454;
reg   [15:0] tmp_4_reg_3454_pp0_iter1_reg;
reg   [15:0] tmp_4_reg_3454_pp0_iter2_reg;
reg   [15:0] tmp_4_reg_3454_pp0_iter3_reg;
reg   [15:0] tmp_4_reg_3454_pp0_iter4_reg;
reg   [15:0] mult_307_V_reg_3472;
reg   [15:0] mult_307_V_reg_3472_pp0_iter1_reg;
reg   [15:0] mult_307_V_reg_3472_pp0_iter2_reg;
reg   [15:0] mult_307_V_reg_3472_pp0_iter3_reg;
reg   [15:0] mult_307_V_reg_3472_pp0_iter4_reg;
reg   [15:0] mult_307_V_reg_3472_pp0_iter5_reg;
reg   [15:0] mult_320_V_reg_3500;
reg   [15:0] mult_320_V_reg_3500_pp0_iter1_reg;
reg   [15:0] mult_320_V_reg_3500_pp0_iter2_reg;
reg   [15:0] mult_320_V_reg_3500_pp0_iter3_reg;
reg   [15:0] mult_320_V_reg_3500_pp0_iter4_reg;
reg   [15:0] mult_320_V_reg_3500_pp0_iter5_reg;
reg   [15:0] mult_386_V_reg_3539;
reg   [15:0] mult_386_V_reg_3539_pp0_iter1_reg;
reg   [15:0] mult_386_V_reg_3539_pp0_iter2_reg;
reg   [15:0] mult_386_V_reg_3539_pp0_iter3_reg;
reg   [15:0] mult_386_V_reg_3539_pp0_iter4_reg;
reg   [15:0] mult_386_V_reg_3539_pp0_iter5_reg;
reg   [15:0] mult_386_V_reg_3539_pp0_iter6_reg;
reg   [15:0] mult_449_V_reg_3582;
reg   [15:0] mult_449_V_reg_3582_pp0_iter1_reg;
reg   [15:0] mult_449_V_reg_3582_pp0_iter2_reg;
reg   [15:0] mult_449_V_reg_3582_pp0_iter3_reg;
reg   [15:0] mult_449_V_reg_3582_pp0_iter4_reg;
reg   [15:0] mult_449_V_reg_3582_pp0_iter5_reg;
reg   [15:0] mult_449_V_reg_3582_pp0_iter6_reg;
reg   [15:0] mult_512_V_reg_3629;
reg   [15:0] mult_512_V_reg_3629_pp0_iter1_reg;
reg   [15:0] mult_512_V_reg_3629_pp0_iter2_reg;
reg   [15:0] mult_512_V_reg_3629_pp0_iter3_reg;
reg   [15:0] mult_512_V_reg_3629_pp0_iter4_reg;
reg   [15:0] mult_512_V_reg_3629_pp0_iter5_reg;
reg   [15:0] mult_512_V_reg_3629_pp0_iter6_reg;
reg   [15:0] mult_576_V_reg_3674;
reg   [15:0] mult_576_V_reg_3674_pp0_iter1_reg;
reg   [15:0] mult_576_V_reg_3674_pp0_iter2_reg;
reg   [15:0] mult_576_V_reg_3674_pp0_iter3_reg;
reg   [15:0] mult_576_V_reg_3674_pp0_iter4_reg;
reg   [15:0] mult_576_V_reg_3674_pp0_iter5_reg;
reg   [15:0] mult_576_V_reg_3674_pp0_iter6_reg;
reg   [15:0] mult_640_V_reg_3716;
reg   [15:0] mult_640_V_reg_3716_pp0_iter1_reg;
reg   [15:0] mult_640_V_reg_3716_pp0_iter2_reg;
reg   [15:0] mult_640_V_reg_3716_pp0_iter3_reg;
reg   [15:0] mult_640_V_reg_3716_pp0_iter4_reg;
reg   [15:0] mult_640_V_reg_3716_pp0_iter5_reg;
reg   [15:0] mult_640_V_reg_3716_pp0_iter6_reg;
reg   [15:0] mult_704_V_reg_3765;
reg   [15:0] mult_704_V_reg_3765_pp0_iter1_reg;
reg   [15:0] mult_704_V_reg_3765_pp0_iter2_reg;
reg   [15:0] mult_704_V_reg_3765_pp0_iter3_reg;
reg   [15:0] mult_704_V_reg_3765_pp0_iter4_reg;
reg   [15:0] mult_704_V_reg_3765_pp0_iter5_reg;
reg   [15:0] mult_704_V_reg_3765_pp0_iter6_reg;
reg   [15:0] mult_704_V_reg_3765_pp0_iter7_reg;
reg   [15:0] mult_770_V_reg_3814;
reg   [15:0] mult_770_V_reg_3814_pp0_iter1_reg;
reg   [15:0] mult_770_V_reg_3814_pp0_iter2_reg;
reg   [15:0] mult_770_V_reg_3814_pp0_iter3_reg;
reg   [15:0] mult_770_V_reg_3814_pp0_iter4_reg;
reg   [15:0] mult_770_V_reg_3814_pp0_iter5_reg;
reg   [15:0] mult_770_V_reg_3814_pp0_iter6_reg;
reg   [15:0] mult_770_V_reg_3814_pp0_iter7_reg;
reg   [15:0] mult_832_V_reg_3861;
reg   [15:0] mult_832_V_reg_3861_pp0_iter1_reg;
reg   [15:0] mult_832_V_reg_3861_pp0_iter2_reg;
reg   [15:0] mult_832_V_reg_3861_pp0_iter3_reg;
reg   [15:0] mult_832_V_reg_3861_pp0_iter4_reg;
reg   [15:0] mult_832_V_reg_3861_pp0_iter5_reg;
reg   [15:0] mult_832_V_reg_3861_pp0_iter6_reg;
reg   [15:0] mult_832_V_reg_3861_pp0_iter7_reg;
reg   [15:0] mult_896_V_reg_3909;
reg   [15:0] mult_896_V_reg_3909_pp0_iter1_reg;
reg   [15:0] mult_896_V_reg_3909_pp0_iter2_reg;
reg   [15:0] mult_896_V_reg_3909_pp0_iter3_reg;
reg   [15:0] mult_896_V_reg_3909_pp0_iter4_reg;
reg   [15:0] mult_896_V_reg_3909_pp0_iter5_reg;
reg   [15:0] mult_896_V_reg_3909_pp0_iter6_reg;
reg   [15:0] mult_896_V_reg_3909_pp0_iter7_reg;
reg   [15:0] mult_960_V_reg_3958;
reg   [15:0] mult_960_V_reg_3958_pp0_iter1_reg;
reg   [15:0] mult_960_V_reg_3958_pp0_iter2_reg;
reg   [15:0] mult_960_V_reg_3958_pp0_iter3_reg;
reg   [15:0] mult_960_V_reg_3958_pp0_iter4_reg;
reg   [15:0] mult_960_V_reg_3958_pp0_iter5_reg;
reg   [15:0] mult_960_V_reg_3958_pp0_iter6_reg;
reg   [15:0] mult_960_V_reg_3958_pp0_iter7_reg;
wire   [15:0] add_ln703_fu_242_p2;
reg   [15:0] add_ln703_reg_4010;
reg   [15:0] add_ln703_reg_4010_pp0_iter1_reg;
reg   [15:0] add_ln703_reg_4010_pp0_iter2_reg;
wire   [15:0] sub_ln703_fu_248_p2;
reg   [15:0] sub_ln703_reg_4017;
reg   [15:0] sub_ln703_reg_4017_pp0_iter2_reg;
wire   [15:0] sub_ln703_531_fu_252_p2;
reg   [15:0] sub_ln703_531_reg_4023;
reg   [15:0] sub_ln703_531_reg_4023_pp0_iter2_reg;
wire   [15:0] sub_ln703_534_fu_256_p2;
reg   [15:0] sub_ln703_534_reg_4029;
reg   [15:0] sub_ln703_534_reg_4029_pp0_iter2_reg;
reg   [15:0] sub_ln703_534_reg_4029_pp0_iter3_reg;
reg   [15:0] sub_ln703_534_reg_4029_pp0_iter4_reg;
wire   [15:0] add_ln703_539_fu_260_p2;
reg   [15:0] add_ln703_539_reg_4035;
reg   [15:0] add_ln703_539_reg_4035_pp0_iter2_reg;
reg   [15:0] add_ln703_539_reg_4035_pp0_iter3_reg;
wire   [15:0] sub_ln703_533_fu_264_p2;
reg   [15:0] sub_ln703_533_reg_4042;
reg   [15:0] sub_ln703_533_reg_4042_pp0_iter3_reg;
reg   [15:0] sub_ln703_533_reg_4042_pp0_iter4_reg;
wire   [15:0] sub_ln703_538_fu_268_p2;
reg   [15:0] sub_ln703_538_reg_4048;
reg   [15:0] sub_ln703_538_reg_4048_pp0_iter3_reg;
reg   [15:0] sub_ln703_538_reg_4048_pp0_iter4_reg;
reg   [15:0] sub_ln703_538_reg_4048_pp0_iter5_reg;
wire   [15:0] add_ln703_543_fu_272_p2;
reg   [15:0] add_ln703_543_reg_4054;
reg   [15:0] add_ln703_543_reg_4054_pp0_iter3_reg;
reg   [15:0] add_ln703_543_reg_4054_pp0_iter4_reg;
wire   [15:0] sub_ln703_532_fu_276_p2;
reg   [15:0] sub_ln703_532_reg_4061;
reg   [15:0] sub_ln703_532_reg_4061_pp0_iter4_reg;
wire   [15:0] add_ln703_538_fu_280_p2;
reg   [15:0] add_ln703_538_reg_4067;
reg   [15:0] add_ln703_538_reg_4067_pp0_iter4_reg;
wire   [15:0] sub_ln703_535_fu_284_p2;
reg   [15:0] sub_ln703_535_reg_4073;
reg   [15:0] sub_ln703_535_reg_4073_pp0_iter4_reg;
wire   [15:0] add_ln703_540_fu_288_p2;
reg   [15:0] add_ln703_540_reg_4079;
reg   [15:0] add_ln703_540_reg_4079_pp0_iter4_reg;
wire   [15:0] sub_ln703_537_fu_292_p2;
reg   [15:0] sub_ln703_537_reg_4085;
reg   [15:0] sub_ln703_537_reg_4085_pp0_iter4_reg;
reg   [15:0] sub_ln703_537_reg_4085_pp0_iter5_reg;
wire   [15:0] sub_ln703_543_fu_296_p2;
reg   [15:0] sub_ln703_543_reg_4091;
reg   [15:0] sub_ln703_543_reg_4091_pp0_iter4_reg;
wire   [15:0] sub_ln703_545_fu_300_p2;
reg   [15:0] sub_ln703_545_reg_4097;
reg   [15:0] sub_ln703_545_reg_4097_pp0_iter4_reg;
reg   [15:0] sub_ln703_545_reg_4097_pp0_iter5_reg;
wire   [15:0] add_ln703_549_fu_304_p2;
reg   [15:0] add_ln703_549_reg_4103;
reg   [15:0] add_ln703_549_reg_4103_pp0_iter4_reg;
reg   [15:0] add_ln703_549_reg_4103_pp0_iter5_reg;
wire   [15:0] sub_ln703_540_fu_308_p2;
reg   [15:0] sub_ln703_540_reg_4110;
reg   [15:0] sub_ln703_540_reg_4110_pp0_iter5_reg;
wire   [15:0] add_ln703_544_fu_312_p2;
reg   [15:0] add_ln703_544_reg_4116;
reg   [15:0] add_ln703_544_reg_4116_pp0_iter5_reg;
wire   [15:0] sub_ln703_544_fu_316_p2;
reg   [15:0] sub_ln703_544_reg_4122;
reg   [15:0] sub_ln703_544_reg_4122_pp0_iter5_reg;
wire   [15:0] add_ln703_547_fu_320_p2;
reg   [15:0] add_ln703_547_reg_4128;
wire   [15:0] add_ln703_554_fu_324_p2;
reg   [15:0] add_ln703_554_reg_4134;
reg   [15:0] add_ln703_554_reg_4134_pp0_iter5_reg;
wire   [15:0] sub_ln703_558_fu_328_p2;
reg   [15:0] sub_ln703_558_reg_4140;
reg   [15:0] sub_ln703_558_reg_4140_pp0_iter5_reg;
wire   [15:0] add_ln703_559_fu_332_p2;
reg   [15:0] add_ln703_559_reg_4146;
reg   [15:0] add_ln703_559_reg_4146_pp0_iter5_reg;
wire   [15:0] add_ln703_560_fu_336_p2;
reg   [15:0] add_ln703_560_reg_4153;
reg   [15:0] add_ln703_560_reg_4153_pp0_iter5_reg;
wire   [15:0] sub_ln703_536_fu_340_p2;
reg   [15:0] sub_ln703_536_reg_4159;
wire   [15:0] sub_ln703_539_fu_344_p2;
reg   [15:0] sub_ln703_539_reg_4165;
wire   [15:0] add_ln703_541_fu_348_p2;
reg   [15:0] add_ln703_541_reg_4171;
wire   [15:0] add_ln703_542_fu_352_p2;
reg   [15:0] add_ln703_542_reg_4177;
wire   [15:0] add_ln703_545_fu_364_p2;
reg   [15:0] add_ln703_545_reg_4183;
wire   [15:0] add_ln703_548_fu_368_p2;
reg   [15:0] add_ln703_548_reg_4188;
wire   [15:0] sub_ln703_549_fu_372_p2;
reg   [15:0] sub_ln703_549_reg_4194;
wire   [15:0] sub_ln703_550_fu_376_p2;
reg   [15:0] sub_ln703_550_reg_4200;
wire   [15:0] sub_ln703_551_fu_380_p2;
reg   [15:0] sub_ln703_551_reg_4205;
wire   [15:0] add_ln703_550_fu_384_p2;
reg   [15:0] add_ln703_550_reg_4211;
wire   [15:0] sub_ln703_552_fu_388_p2;
reg   [15:0] sub_ln703_552_reg_4217;
wire   [15:0] add_ln703_551_fu_393_p2;
reg   [15:0] add_ln703_551_reg_4222;
wire   [15:0] sub_ln703_554_fu_398_p2;
reg   [15:0] sub_ln703_554_reg_4228;
wire   [15:0] sub_ln703_557_fu_402_p2;
reg   [15:0] sub_ln703_557_reg_4234;
wire   [15:0] add_ln703_564_fu_406_p2;
reg   [15:0] add_ln703_564_reg_4240;
wire   [15:0] sub_ln703_570_fu_410_p2;
reg   [15:0] sub_ln703_570_reg_4246;
wire   [15:0] sub_ln703_576_fu_414_p2;
reg   [15:0] sub_ln703_576_reg_4252;
reg   [15:0] sub_ln703_576_reg_4252_pp0_iter6_reg;
wire   [15:0] add_ln703_566_fu_418_p2;
reg   [15:0] add_ln703_566_reg_4258;
reg   [15:0] add_ln703_566_reg_4258_pp0_iter6_reg;
wire   [15:0] sub_ln703_584_fu_422_p2;
reg   [15:0] sub_ln703_584_reg_4264;
reg   [15:0] sub_ln703_584_reg_4264_pp0_iter6_reg;
wire   [15:0] add_ln703_568_fu_426_p2;
reg   [15:0] add_ln703_568_reg_4270;
wire   [15:0] sub_ln703_591_fu_430_p2;
reg   [15:0] sub_ln703_591_reg_4277;
wire   [15:0] add_ln703_597_fu_434_p2;
reg   [15:0] add_ln703_597_reg_4282;
reg   [15:0] add_ln703_597_reg_4282_pp0_iter6_reg;
wire   [15:0] add_ln703_557_fu_488_p2;
reg   [15:0] add_ln703_557_reg_4293;
wire   [15:0] add_ln703_558_fu_498_p2;
reg   [15:0] add_ln703_558_reg_4298;
wire   [15:0] sub_ln703_567_fu_540_p2;
reg   [15:0] sub_ln703_567_reg_4303;
wire   [15:0] sub_ln703_572_fu_563_p2;
reg   [15:0] sub_ln703_572_reg_4309;
wire   [15:0] sub_ln703_574_fu_572_p2;
reg   [15:0] sub_ln703_574_reg_4314;
wire   [15:0] sub_ln703_578_fu_585_p2;
reg   [15:0] sub_ln703_578_reg_4319;
wire   [15:0] sub_ln703_579_fu_590_p2;
reg   [15:0] sub_ln703_579_reg_4324;
wire   [15:0] sub_ln703_582_fu_599_p2;
reg   [15:0] sub_ln703_582_reg_4329;
wire   [15:0] sub_ln703_585_fu_609_p2;
reg   [15:0] sub_ln703_585_reg_4334;
wire   [15:0] sub_ln703_586_fu_614_p2;
reg   [15:0] sub_ln703_586_reg_4340;
wire   [15:0] sub_ln703_587_fu_619_p2;
reg   [15:0] sub_ln703_587_reg_4345;
wire   [15:0] sub_ln703_588_fu_624_p2;
reg   [15:0] sub_ln703_588_reg_4350;
wire   [15:0] sub_ln703_589_fu_638_p2;
reg   [15:0] sub_ln703_589_reg_4355;
wire   [15:0] sub_ln703_590_fu_643_p2;
reg   [15:0] sub_ln703_590_reg_4361;
wire   [15:0] sub_ln703_592_fu_653_p2;
reg   [15:0] sub_ln703_592_reg_4366;
wire   [15:0] add_ln703_571_fu_657_p2;
reg   [15:0] add_ln703_571_reg_4372;
wire   [15:0] sub_ln703_594_fu_666_p2;
reg   [15:0] sub_ln703_594_reg_4377;
wire   [15:0] add_ln703_572_fu_670_p2;
reg   [15:0] add_ln703_572_reg_4382;
wire   [15:0] add_ln703_573_fu_675_p2;
reg   [15:0] add_ln703_573_reg_4387;
wire   [15:0] add_ln703_574_fu_679_p2;
reg   [15:0] add_ln703_574_reg_4393;
wire   [15:0] sub_ln703_596_fu_683_p2;
reg   [15:0] sub_ln703_596_reg_4398;
wire   [15:0] sub_ln703_599_fu_693_p2;
reg   [15:0] sub_ln703_599_reg_4403;
wire   [15:0] add_ln703_576_fu_702_p2;
reg   [15:0] add_ln703_576_reg_4408;
wire   [15:0] add_ln703_577_fu_707_p2;
reg   [15:0] add_ln703_577_reg_4413;
wire   [15:0] add_ln703_579_fu_716_p2;
reg   [15:0] add_ln703_579_reg_4418;
wire   [15:0] sub_ln703_605_fu_720_p2;
reg   [15:0] sub_ln703_605_reg_4423;
wire   [15:0] sub_ln703_608_fu_725_p2;
reg   [15:0] sub_ln703_608_reg_4428;
wire   [15:0] add_ln703_580_fu_730_p2;
reg   [15:0] add_ln703_580_reg_4433;
wire   [15:0] sub_ln703_610_fu_734_p2;
reg   [15:0] sub_ln703_610_reg_4439;
wire   [15:0] sub_ln703_611_fu_739_p2;
reg   [15:0] sub_ln703_611_reg_4444;
wire   [15:0] add_ln703_583_fu_754_p2;
reg   [15:0] add_ln703_583_reg_4450;
wire   [15:0] sub_ln703_613_fu_758_p2;
reg   [15:0] sub_ln703_613_reg_4455;
wire   [15:0] sub_ln703_617_fu_763_p2;
reg   [15:0] sub_ln703_617_reg_4460;
wire   [15:0] sub_ln703_620_fu_772_p2;
reg   [15:0] sub_ln703_620_reg_4466;
wire   [15:0] add_ln703_587_fu_786_p2;
reg   [15:0] add_ln703_587_reg_4471;
wire   [15:0] add_ln703_588_fu_792_p2;
reg   [15:0] add_ln703_588_reg_4476;
wire   [15:0] add_ln703_590_fu_801_p2;
reg   [15:0] add_ln703_590_reg_4481;
wire   [15:0] sub_ln703_627_fu_807_p2;
reg   [15:0] sub_ln703_627_reg_4486;
wire   [15:0] sub_ln703_632_fu_818_p2;
reg   [15:0] sub_ln703_632_reg_4491;
wire   [15:0] sub_ln703_641_fu_838_p2;
reg   [15:0] sub_ln703_641_reg_4496;
wire   [15:0] sub_ln703_645_fu_843_p2;
reg   [15:0] sub_ln703_645_reg_4501;
wire   [15:0] sub_ln703_660_fu_872_p2;
reg   [15:0] sub_ln703_660_reg_4506;
wire   [15:0] sub_ln703_661_fu_877_p2;
reg   [15:0] sub_ln703_661_reg_4511;
wire   [15:0] sub_ln703_662_fu_882_p2;
reg   [15:0] sub_ln703_662_reg_4516;
wire   [15:0] add_ln703_611_fu_887_p2;
reg   [15:0] add_ln703_611_reg_4521;
wire   [15:0] add_ln703_620_fu_891_p2;
reg   [15:0] add_ln703_620_reg_4537;
wire   [15:0] sub_ln703_671_fu_896_p2;
reg   [15:0] sub_ln703_671_reg_4543;
wire   [15:0] sub_ln703_676_fu_901_p2;
reg   [15:0] sub_ln703_676_reg_4548;
wire   [15:0] add_ln703_637_fu_906_p2;
reg   [15:0] add_ln703_637_reg_4553;
wire   [15:0] add_ln703_655_fu_910_p2;
reg   [15:0] add_ln703_655_reg_4558;
wire   [15:0] add_ln703_659_fu_914_p2;
reg   [15:0] add_ln703_659_reg_4568;
wire   [15:0] add_ln703_692_fu_920_p2;
reg   [15:0] add_ln703_692_reg_4573;
reg   [15:0] add_ln703_692_reg_4573_pp0_iter7_reg;
wire   [15:0] add_ln703_631_fu_1397_p2;
reg   [15:0] add_ln703_631_reg_4588;
wire   [15:0] add_ln703_634_fu_1416_p2;
reg   [15:0] add_ln703_634_reg_4593;
wire   [15:0] sub_ln703_692_fu_1433_p2;
reg   [15:0] sub_ln703_692_reg_4598;
wire   [15:0] sub_ln703_693_fu_1438_p2;
reg   [15:0] sub_ln703_693_reg_4603;
wire   [15:0] add_ln703_639_fu_1459_p2;
reg   [15:0] add_ln703_639_reg_4608;
wire   [15:0] sub_ln703_695_fu_1464_p2;
reg   [15:0] sub_ln703_695_reg_4613;
wire   [15:0] sub_ln703_699_fu_1495_p2;
reg   [15:0] sub_ln703_699_reg_4618;
wire   [15:0] sub_ln703_700_fu_1500_p2;
reg   [15:0] sub_ln703_700_reg_4623;
wire   [15:0] add_ln703_642_fu_1505_p2;
reg   [15:0] add_ln703_642_reg_4628;
wire   [15:0] sub_ln703_701_fu_1509_p2;
reg   [15:0] sub_ln703_701_reg_4633;
wire   [15:0] sub_ln703_702_fu_1514_p2;
reg   [15:0] sub_ln703_702_reg_4638;
wire   [15:0] sub_ln703_704_fu_1524_p2;
reg   [15:0] sub_ln703_704_reg_4643;
wire   [15:0] add_ln703_645_fu_1538_p2;
reg   [15:0] add_ln703_645_reg_4648;
wire   [15:0] sub_ln703_706_fu_1548_p2;
reg   [15:0] sub_ln703_706_reg_4653;
wire   [15:0] add_ln703_646_fu_1553_p2;
reg   [15:0] add_ln703_646_reg_4658;
wire   [15:0] sub_ln703_707_fu_1559_p2;
reg   [15:0] sub_ln703_707_reg_4663;
wire   [15:0] sub_ln703_708_fu_1564_p2;
reg   [15:0] sub_ln703_708_reg_4668;
wire   [15:0] sub_ln703_709_fu_1569_p2;
reg   [15:0] sub_ln703_709_reg_4673;
wire   [15:0] sub_ln703_710_fu_1606_p2;
reg   [15:0] sub_ln703_710_reg_4678;
wire   [15:0] sub_ln703_711_fu_1611_p2;
reg   [15:0] sub_ln703_711_reg_4683;
wire   [15:0] sub_ln703_712_fu_1616_p2;
reg   [15:0] sub_ln703_712_reg_4688;
wire   [15:0] sub_ln703_714_fu_1626_p2;
reg   [15:0] sub_ln703_714_reg_4693;
wire   [15:0] sub_ln703_715_fu_1631_p2;
reg   [15:0] sub_ln703_715_reg_4698;
wire   [15:0] sub_ln703_716_fu_1636_p2;
reg   [15:0] sub_ln703_716_reg_4703;
wire   [15:0] sub_ln703_718_fu_1646_p2;
reg   [15:0] sub_ln703_718_reg_4708;
wire   [15:0] sub_ln703_720_fu_1676_p2;
reg   [15:0] sub_ln703_720_reg_4713;
wire   [15:0] sub_ln703_722_fu_1681_p2;
reg   [15:0] sub_ln703_722_reg_4718;
wire   [15:0] sub_ln703_724_fu_1686_p2;
reg   [15:0] sub_ln703_724_reg_4723;
wire   [15:0] sub_ln703_725_fu_1691_p2;
reg   [15:0] sub_ln703_725_reg_4728;
wire   [15:0] add_ln703_658_fu_1696_p2;
reg   [15:0] add_ln703_658_reg_4733;
wire   [15:0] sub_ln703_727_fu_1701_p2;
reg   [15:0] sub_ln703_727_reg_4738;
wire   [15:0] add_ln703_661_fu_1710_p2;
reg   [15:0] add_ln703_661_reg_4744;
wire   [15:0] sub_ln703_729_fu_1715_p2;
reg   [15:0] sub_ln703_729_reg_4749;
wire   [15:0] sub_ln703_730_fu_1720_p2;
reg   [15:0] sub_ln703_730_reg_4754;
wire   [15:0] sub_ln703_731_fu_1725_p2;
reg   [15:0] sub_ln703_731_reg_4759;
wire   [15:0] add_ln703_663_fu_1735_p2;
reg   [15:0] add_ln703_663_reg_4764;
wire   [15:0] sub_ln703_732_fu_1741_p2;
reg   [15:0] sub_ln703_732_reg_4769;
wire   [15:0] sub_ln703_738_fu_1757_p2;
reg   [15:0] sub_ln703_738_reg_4774;
wire   [15:0] sub_ln703_742_fu_1762_p2;
reg   [15:0] sub_ln703_742_reg_4779;
wire   [15:0] add_ln703_667_fu_1767_p2;
reg   [15:0] add_ln703_667_reg_4784;
wire   [15:0] sub_ln703_743_fu_1772_p2;
reg   [15:0] sub_ln703_743_reg_4789;
wire   [15:0] sub_ln703_744_fu_1777_p2;
reg   [15:0] sub_ln703_744_reg_4794;
wire   [15:0] sub_ln703_745_fu_1782_p2;
reg   [15:0] sub_ln703_745_reg_4799;
wire   [15:0] add_ln703_669_fu_1787_p2;
reg   [15:0] add_ln703_669_reg_4804;
wire   [15:0] sub_ln703_748_fu_1792_p2;
reg   [15:0] sub_ln703_748_reg_4809;
wire   [15:0] sub_ln703_751_fu_1797_p2;
reg   [15:0] sub_ln703_751_reg_4814;
wire   [15:0] add_ln703_670_fu_1802_p2;
reg   [15:0] add_ln703_670_reg_4819;
wire   [15:0] sub_ln703_752_fu_1807_p2;
reg   [15:0] sub_ln703_752_reg_4824;
wire   [15:0] add_ln703_672_fu_1812_p2;
reg   [15:0] add_ln703_672_reg_4829;
wire   [15:0] sub_ln703_753_fu_1817_p2;
reg   [15:0] sub_ln703_753_reg_4834;
wire   [15:0] add_ln703_674_fu_1822_p2;
reg   [15:0] add_ln703_674_reg_4839;
wire   [15:0] add_ln703_679_fu_1826_p2;
reg   [15:0] add_ln703_679_reg_4847;
wire   [15:0] sub_ln703_765_fu_1832_p2;
reg   [15:0] sub_ln703_765_reg_4852;
wire   [15:0] add_ln703_687_fu_1847_p2;
reg   [15:0] add_ln703_687_reg_4857;
wire   [15:0] add_ln703_688_fu_1853_p2;
reg   [15:0] add_ln703_688_reg_4862;
wire   [15:0] add_ln703_707_fu_1877_p2;
reg   [15:0] add_ln703_707_reg_4867;
wire   [15:0] add_ln703_711_fu_1887_p2;
reg   [15:0] add_ln703_711_reg_4872;
wire   [15:0] add_ln703_716_fu_1902_p2;
reg   [15:0] add_ln703_716_reg_4877;
wire   [15:0] add_ln703_722_fu_1913_p2;
reg   [15:0] add_ln703_722_reg_4882;
wire   [15:0] add_ln703_724_fu_1923_p2;
reg   [15:0] add_ln703_724_reg_4887;
wire   [15:0] add_ln703_727_fu_1934_p2;
reg   [15:0] add_ln703_727_reg_4892;
wire   [15:0] add_ln703_729_fu_1945_p2;
reg   [15:0] add_ln703_729_reg_4897;
wire   [15:0] add_ln703_732_fu_1956_p2;
reg   [15:0] add_ln703_732_reg_4902;
wire   [15:0] add_ln703_737_fu_1962_p2;
reg   [15:0] add_ln703_737_reg_4907;
wire   [15:0] add_ln703_739_fu_1966_p2;
reg   [15:0] add_ln703_739_reg_4915;
wire   [15:0] add_ln703_751_fu_1971_p2;
reg   [15:0] add_ln703_751_reg_4920;
wire    ap_block_pp0_stage0;
wire   [15:0] sub_ln703_541_fu_356_p2;
wire   [15:0] sub_ln703_542_fu_360_p2;
wire   [15:0] add_ln703_546_fu_438_p2;
wire   [15:0] sub_ln703_546_fu_442_p2;
wire   [15:0] sub_ln703_547_fu_446_p2;
wire   [15:0] sub_ln703_548_fu_450_p2;
wire   [15:0] add_ln703_552_fu_454_p2;
wire   [15:0] add_ln703_553_fu_458_p2;
wire   [15:0] sub_ln703_553_fu_462_p2;
wire   [15:0] add_ln703_555_fu_466_p2;
wire   [15:0] sub_ln703_555_fu_470_p2;
wire   [15:0] sub_ln703_556_fu_474_p2;
wire   [15:0] add_ln703_556_fu_478_p2;
wire   [15:0] sub_ln703_559_fu_483_p2;
wire   [15:0] sub_ln703_560_fu_493_p2;
wire   [15:0] sub_ln703_561_fu_502_p2;
wire   [15:0] sub_ln703_562_fu_506_p2;
wire   [15:0] add_ln703_561_fu_510_p2;
wire   [15:0] add_ln703_562_fu_522_p2;
wire   [15:0] add_ln703_567_fu_629_p2;
wire   [15:0] add_ln703_563_fu_526_p2;
wire   [15:0] sub_ln703_565_fu_530_p2;
wire   [15:0] sub_ln703_566_fu_535_p2;
wire   [15:0] sub_ln703_568_fu_545_p2;
wire   [15:0] sub_ln703_569_fu_549_p2;
wire   [15:0] add_ln703_565_fu_554_p2;
wire   [15:0] sub_ln703_571_fu_558_p2;
wire   [15:0] sub_ln703_573_fu_567_p2;
wire   [15:0] sub_ln703_575_fu_577_p2;
wire   [15:0] sub_ln703_577_fu_581_p2;
wire   [15:0] sub_ln703_580_fu_594_p2;
wire   [15:0] sub_ln703_583_fu_604_p2;
wire   [15:0] sub_ln703_564_fu_518_p2;
wire   [15:0] add_ln703_581_fu_744_p2;
wire   [15:0] add_ln703_569_fu_633_p2;
wire   [15:0] add_ln703_570_fu_648_p2;
wire   [15:0] sub_ln703_593_fu_661_p2;
wire   [15:0] add_ln703_585_fu_777_p2;
wire   [15:0] add_ln703_586_fu_781_p2;
wire   [15:0] sub_ln703_597_fu_688_p2;
wire   [15:0] add_ln703_589_fu_797_p2;
wire   [15:0] add_ln703_575_fu_698_p2;
wire   [15:0] sub_ln703_602_fu_712_p2;
wire   [15:0] add_ln703_595_fu_828_p2;
wire   [15:0] add_ln703_582_fu_748_p2;
wire   [15:0] sub_ln703_618_fu_768_p2;
wire   [15:0] add_ln703_600_fu_848_p2;
wire   [15:0] add_ln703_601_fu_852_p2;
wire   [15:0] add_ln703_605_fu_862_p2;
wire   [15:0] add_ln703_593_fu_812_p2;
wire   [15:0] add_ln703_594_fu_823_p2;
wire   [15:0] add_ln703_596_fu_832_p2;
wire   [15:0] add_ln703_602_fu_856_p2;
wire   [15:0] add_ln703_606_fu_866_p2;
wire   [15:0] sub_ln703_563_fu_514_p2;
wire   [15:0] sub_ln703_581_fu_924_p2;
wire   [15:0] sub_ln703_595_fu_928_p2;
wire   [15:0] sub_ln703_600_fu_936_p2;
wire   [15:0] add_ln703_578_fu_944_p2;
wire   [15:0] sub_ln703_607_fu_961_p2;
wire   [15:0] sub_ln703_609_fu_965_p2;
wire   [15:0] sub_ln703_612_fu_969_p2;
wire   [15:0] add_ln703_584_fu_985_p2;
wire   [15:0] sub_ln703_621_fu_993_p2;
wire   [15:0] sub_ln703_623_fu_1002_p2;
wire   [15:0] sub_ln703_624_fu_1006_p2;
wire   [15:0] sub_ln703_625_fu_1010_p2;
wire   [15:0] sub_ln703_598_fu_932_p2;
wire   [15:0] add_ln703_591_fu_1027_p2;
wire   [15:0] add_ln703_592_fu_1031_p2;
wire   [15:0] sub_ln703_630_fu_1035_p2;
wire   [15:0] sub_ln703_631_fu_1039_p2;
wire   [15:0] add_ln703_598_fu_1052_p2;
wire   [15:0] sub_ln703_604_fu_952_p2;
wire   [15:0] sub_ln703_635_fu_1056_p2;
wire   [15:0] sub_ln703_637_fu_1065_p2;
wire   [15:0] sub_ln703_638_fu_1069_p2;
wire   [15:0] add_ln703_599_fu_1073_p2;
wire   [15:0] sub_ln703_639_fu_1078_p2;
wire   [15:0] sub_ln703_643_fu_1091_p2;
wire   [15:0] sub_ln703_644_fu_1095_p2;
wire   [15:0] sub_ln703_615_fu_977_p2;
wire   [15:0] sub_ln703_616_fu_981_p2;
wire   [15:0] sub_ln703_646_fu_1099_p2;
wire   [15:0] sub_ln703_636_fu_1060_p2;
wire   [15:0] sub_ln703_647_fu_1104_p2;
wire   [15:0] sub_ln703_648_fu_1108_p2;
wire   [15:0] sub_ln703_649_fu_1113_p2;
wire   [15:0] sub_ln703_651_fu_1122_p2;
wire   [15:0] sub_ln703_652_fu_1127_p2;
wire   [15:0] add_ln703_603_fu_1132_p2;
wire   [15:0] sub_ln703_653_fu_1136_p2;
wire   [15:0] add_ln703_604_fu_1140_p2;
wire   [15:0] sub_ln703_655_fu_1149_p2;
wire   [15:0] sub_ln703_629_fu_1022_p2;
wire   [15:0] sub_ln703_656_fu_1153_p2;
wire   [15:0] add_ln703_626_fu_1321_p2;
wire   [15:0] sub_ln703_657_fu_1158_p2;
wire   [15:0] add_ln703_607_fu_1163_p2;
wire   [15:0] sub_ln703_658_fu_1167_p2;
wire   [15:0] sub_ln703_659_fu_1171_p2;
wire   [15:0] sub_ln703_601_fu_940_p2;
wire   [15:0] add_ln703_628_fu_1350_p2;
wire   [15:0] add_ln703_608_fu_1176_p2;
wire   [15:0] add_ln703_609_fu_1181_p2;
wire   [15:0] add_ln703_610_fu_1185_p2;
wire   [15:0] sub_ln703_634_fu_1048_p2;
wire   [15:0] sub_ln703_663_fu_1189_p2;
wire   [15:0] add_ln703_612_fu_1194_p2;
wire   [15:0] sub_ln703_664_fu_1199_p2;
wire   [15:0] sub_ln703_606_fu_956_p2;
wire   [15:0] add_ln703_632_fu_1407_p2;
wire   [15:0] add_ln703_633_fu_1412_p2;
wire   [15:0] sub_ln703_665_fu_1204_p2;
wire   [15:0] add_ln703_613_fu_1209_p2;
wire   [15:0] sub_ln703_666_fu_1214_p2;
wire   [15:0] add_ln703_614_fu_1219_p2;
wire   [15:0] sub_ln703_640_fu_1082_p2;
wire   [15:0] add_ln703_638_fu_1454_p2;
wire   [15:0] sub_ln703_667_fu_1224_p2;
wire   [15:0] sub_ln703_642_fu_1086_p2;
wire   [15:0] add_ln703_615_fu_1228_p2;
wire   [15:0] sub_ln703_668_fu_1233_p2;
wire   [15:0] add_ln703_616_fu_1238_p2;
wire   [15:0] add_ln703_617_fu_1243_p2;
wire   [15:0] add_ln703_618_fu_1248_p2;
wire   [15:0] add_ln703_619_fu_1252_p2;
wire   [15:0] add_ln703_621_fu_1256_p2;
wire   [15:0] sub_ln703_669_fu_1261_p2;
wire   [15:0] sub_ln703_670_fu_1266_p2;
wire   [15:0] add_ln703_622_fu_1271_p2;
wire   [15:0] add_ln703_643_fu_1529_p2;
wire   [15:0] add_ln703_644_fu_1533_p2;
wire   [15:0] add_ln703_623_fu_1276_p2;
wire   [15:0] sub_ln703_650_fu_1118_p2;
wire   [15:0] sub_ln703_672_fu_1281_p2;
wire   [15:0] add_ln703_624_fu_1286_p2;
wire   [15:0] sub_ln703_674_fu_1296_p2;
wire   [15:0] sub_ln703_626_fu_1014_p2;
wire   [15:0] add_ln703_648_fu_1579_p2;
wire   [15:0] sub_ln703_677_fu_1306_p2;
wire   [15:0] sub_ln703_628_fu_1018_p2;
wire   [15:0] add_ln703_651_fu_1595_p2;
wire   [15:0] add_ln703_625_fu_1311_p2;
wire   [15:0] sub_ln703_678_fu_1316_p2;
wire   [15:0] add_ln703_627_fu_1325_p2;
wire   [15:0] sub_ln703_681_fu_1340_p2;
wire   [15:0] sub_ln703_682_fu_1345_p2;
wire   [15:0] add_ln703_629_fu_1355_p2;
wire   [15:0] sub_ln703_683_fu_1360_p2;
wire   [15:0] sub_ln703_684_fu_1365_p2;
wire   [15:0] sub_ln703_686_fu_1374_p2;
wire   [15:0] sub_ln703_687_fu_1378_p2;
wire   [15:0] add_ln703_630_fu_1387_p2;
wire   [15:0] sub_ln703_603_fu_948_p2;
wire   [15:0] add_ln703_654_fu_1661_p2;
wire   [15:0] add_ln703_656_fu_1666_p2;
wire   [15:0] sub_ln703_689_fu_1392_p2;
wire   [15:0] sub_ln703_690_fu_1402_p2;
wire   [15:0] add_ln703_635_fu_1422_p2;
wire   [15:0] sub_ln703_691_fu_1428_p2;
wire   [15:0] sub_ln703_694_fu_1443_p2;
wire   [15:0] add_ln703_636_fu_1448_p2;
wire   [15:0] add_ln703_660_fu_1706_p2;
wire   [15:0] add_ln703_640_fu_1469_p2;
wire   [15:0] sub_ln703_696_fu_1475_p2;
wire   [15:0] add_ln703_641_fu_1480_p2;
wire   [15:0] sub_ln703_614_fu_973_p2;
wire   [15:0] add_ln703_662_fu_1730_p2;
wire   [15:0] sub_ln703_697_fu_1485_p2;
wire   [15:0] sub_ln703_619_fu_989_p2;
wire   [15:0] add_ln703_665_fu_1746_p2;
wire   [15:0] sub_ln703_705_fu_1544_p2;
wire   [15:0] add_ln703_647_fu_1574_p2;
wire   [15:0] sub_ln703_675_fu_1301_p2;
wire   [15:0] add_ln703_649_fu_1584_p2;
wire   [15:0] add_ln703_650_fu_1590_p2;
wire   [15:0] add_ln703_652_fu_1600_p2;
wire   [15:0] sub_ln703_680_fu_1335_p2;
wire   [15:0] sub_ln703_713_fu_1621_p2;
wire   [15:0] sub_ln703_717_fu_1641_p2;
wire   [15:0] sub_ln703_685_fu_1370_p2;
wire   [15:0] add_ln703_653_fu_1651_p2;
wire   [15:0] sub_ln703_719_fu_1656_p2;
wire   [15:0] add_ln703_657_fu_1670_p2;
wire   [15:0] sub_ln703_698_fu_1490_p2;
wire   [15:0] add_ln703_666_fu_1751_p2;
wire   [15:0] sub_ln703_654_fu_1145_p2;
wire   [15:0] add_ln703_685_fu_1837_p2;
wire   [15:0] add_ln703_686_fu_1842_p2;
wire   [15:0] sub_ln703_679_fu_1330_p2;
wire   [15:0] add_ln703_703_fu_1858_p2;
wire   [15:0] add_ln703_705_fu_1867_p2;
wire   [15:0] add_ln703_704_fu_1862_p2;
wire   [15:0] add_ln703_706_fu_1871_p2;
wire   [15:0] add_ln703_710_fu_1883_p2;
wire   [15:0] sub_ln703_622_fu_997_p2;
wire   [15:0] add_ln703_714_fu_1893_p2;
wire   [15:0] add_ln703_715_fu_1898_p2;
wire   [15:0] sub_ln703_673_fu_1291_p2;
wire   [15:0] add_ln703_721_fu_1908_p2;
wire   [15:0] add_ln703_723_fu_1919_p2;
wire   [15:0] add_ln703_726_fu_1929_p2;
wire   [15:0] sub_ln703_633_fu_1043_p2;
wire   [15:0] add_ln703_728_fu_1940_p2;
wire   [15:0] sub_ln703_688_fu_1382_p2;
wire   [15:0] add_ln703_731_fu_1951_p2;
wire   [15:0] sub_ln703_703_fu_1519_p2;
wire   [15:0] sub_ln703_723_fu_1979_p2;
wire   [15:0] sub_ln703_726_fu_1983_p2;
wire   [15:0] add_ln703_664_fu_1991_p2;
wire   [15:0] sub_ln703_736_fu_2007_p2;
wire   [15:0] sub_ln703_739_fu_2015_p2;
wire   [15:0] sub_ln703_740_fu_2019_p2;
wire   [15:0] sub_ln703_741_fu_2023_p2;
wire   [15:0] sub_ln703_746_fu_2027_p2;
wire   [15:0] sub_ln703_747_fu_2031_p2;
wire   [15:0] add_ln703_668_fu_2035_p2;
wire   [15:0] sub_ln703_749_fu_2039_p2;
wire   [15:0] sub_ln703_750_fu_2043_p2;
wire   [15:0] add_ln703_671_fu_2047_p2;
wire   [15:0] sub_ln703_754_fu_2051_p2;
wire   [15:0] sub_ln703_721_fu_1975_p2;
wire   [15:0] sub_ln703_755_fu_2055_p2;
wire   [15:0] sub_ln703_757_fu_2064_p2;
wire   [15:0] add_ln703_673_fu_2068_p2;
wire   [15:0] add_ln703_675_fu_2072_p2;
wire   [15:0] sub_ln703_758_fu_2076_p2;
wire   [15:0] sub_ln703_759_fu_2081_p2;
wire   [15:0] sub_ln703_728_fu_1987_p2;
wire   [15:0] sub_ln703_761_fu_2089_p2;
wire   [15:0] add_ln703_676_fu_2093_p2;
wire   [15:0] sub_ln703_762_fu_2097_p2;
wire   [15:0] add_ln703_677_fu_2101_p2;
wire   [15:0] sub_ln703_763_fu_2105_p2;
wire   [15:0] add_ln703_678_fu_2109_p2;
wire   [15:0] sub_ln703_733_fu_1995_p2;
wire   [15:0] sub_ln703_734_fu_1999_p2;
wire   [15:0] sub_ln703_735_fu_2003_p2;
wire   [15:0] add_ln703_680_fu_2118_p2;
wire   [15:0] add_ln703_708_fu_2323_p2;
wire   [15:0] sub_ln703_737_fu_2011_p2;
wire   [15:0] sub_ln703_766_fu_2123_p2;
wire   [15:0] add_ln703_717_fu_2342_p2;
wire   [15:0] add_ln703_681_fu_2132_p2;
wire   [15:0] add_ln703_682_fu_2136_p2;
wire   [15:0] add_ln703_719_fu_2361_p2;
wire   [15:0] add_ln703_683_fu_2146_p2;
wire   [15:0] sub_ln703_769_fu_2150_p2;
wire   [15:0] add_ln703_684_fu_2154_p2;
wire   [15:0] sub_ln703_770_fu_2158_p2;
wire   [15:0] sub_ln703_771_fu_2162_p2;
wire   [15:0] add_ln703_689_fu_2181_p2;
wire   [15:0] sub_ln703_775_fu_2185_p2;
wire   [15:0] add_ln703_690_fu_2189_p2;
wire   [15:0] add_ln703_691_fu_2193_p2;
wire   [15:0] sub_ln703_778_fu_2207_p2;
wire   [15:0] sub_ln703_779_fu_2211_p2;
wire   [15:0] sub_ln703_780_fu_2215_p2;
wire   [15:0] sub_ln703_781_fu_2220_p2;
wire   [15:0] sub_ln703_782_fu_2224_p2;
wire   [15:0] add_ln703_693_fu_2229_p2;
wire   [15:0] add_ln703_694_fu_2234_p2;
wire   [15:0] add_ln703_695_fu_2239_p2;
wire   [15:0] sub_ln703_783_fu_2244_p2;
wire   [15:0] sub_ln703_784_fu_2249_p2;
wire   [15:0] sub_ln703_786_fu_2259_p2;
wire   [15:0] add_ln703_696_fu_2264_p2;
wire   [15:0] add_ln703_697_fu_2269_p2;
wire   [15:0] sub_ln703_787_fu_2274_p2;
wire   [15:0] add_ln703_698_fu_2279_p2;
wire   [15:0] sub_ln703_788_fu_2284_p2;
wire   [15:0] add_ln703_699_fu_2289_p2;
wire   [15:0] sub_ln703_789_fu_2294_p2;
wire   [15:0] add_ln703_700_fu_2303_p2;
wire   [15:0] add_ln703_701_fu_2308_p2;
wire   [15:0] add_ln703_702_fu_2313_p2;
wire   [15:0] add_ln703_740_fu_2532_p2;
wire   [15:0] add_ln703_709_fu_2327_p2;
wire   [15:0] add_ln703_712_fu_2332_p2;
wire   [15:0] add_ln703_713_fu_2337_p2;
wire   [15:0] add_ln703_718_fu_2346_p2;
wire   [15:0] sub_ln703_792_fu_2351_p2;
wire   [15:0] add_ln703_720_fu_2365_p2;
wire   [15:0] sub_ln703_768_fu_2141_p2;
wire   [15:0] sub_ln703_794_fu_2370_p2;
wire   [15:0] sub_ln703_795_fu_2375_p2;
wire   [15:0] sub_ln703_796_fu_2380_p2;
wire   [15:0] add_ln703_725_fu_2389_p2;
wire   [15:0] sub_ln703_798_fu_2394_p2;
wire   [15:0] sub_ln703_799_fu_2399_p2;
wire   [15:0] sub_ln703_800_fu_2404_p2;
wire   [15:0] sub_ln703_801_fu_2409_p2;
wire   [15:0] sub_ln703_802_fu_2414_p2;
wire   [15:0] sub_ln703_776_fu_2197_p2;
wire   [15:0] sub_ln703_803_fu_2419_p2;
wire   [15:0] add_ln703_730_fu_2424_p2;
wire   [15:0] add_ln703_733_fu_2434_p2;
wire   [15:0] add_ln703_750_fu_2669_p2;
wire   [15:0] sub_ln703_805_fu_2439_p2;
wire   [15:0] sub_ln703_806_fu_2444_p2;
wire   [15:0] sub_ln703_807_fu_2449_p2;
wire   [15:0] sub_ln703_756_fu_2059_p2;
wire   [15:0] add_ln703_754_fu_2693_p2;
wire   [15:0] sub_ln703_808_fu_2454_p2;
wire   [15:0] sub_ln703_809_fu_2459_p2;
wire   [15:0] sub_ln703_810_fu_2464_p2;
wire   [15:0] sub_ln703_785_fu_2254_p2;
wire   [15:0] add_ln703_734_fu_2469_p2;
wire   [15:0] sub_ln703_760_fu_2085_p2;
wire   [15:0] add_ln703_758_fu_2728_p2;
wire   [15:0] sub_ln703_811_fu_2474_p2;
wire   [15:0] sub_ln703_812_fu_2479_p2;
wire   [15:0] add_ln703_735_fu_2484_p2;
wire   [15:0] sub_ln703_813_fu_2489_p2;
wire   [15:0] sub_ln703_814_fu_2494_p2;
wire   [15:0] add_ln703_761_fu_2763_p2;
wire   [15:0] add_ln703_762_fu_2767_p2;
wire   [15:0] sub_ln703_815_fu_2499_p2;
wire   [15:0] add_ln703_736_fu_2504_p2;
wire   [15:0] sub_ln703_790_fu_2299_p2;
wire   [15:0] sub_ln703_764_fu_2113_p2;
wire   [15:0] add_ln703_765_fu_2792_p2;
wire   [15:0] sub_ln703_816_fu_2509_p2;
wire   [15:0] sub_ln703_817_fu_2514_p2;
wire   [15:0] sub_ln703_818_fu_2519_p2;
wire   [15:0] sub_ln703_819_fu_2524_p2;
wire   [15:0] sub_ln703_791_fu_2318_p2;
wire   [15:0] add_ln703_738_fu_2528_p2;
wire   [15:0] add_ln703_741_fu_2536_p2;
wire   [15:0] sub_ln703_820_fu_2541_p2;
wire   [15:0] sub_ln703_821_fu_2546_p2;
wire   [15:0] sub_ln703_822_fu_2550_p2;
wire   [15:0] sub_ln703_823_fu_2555_p2;
wire   [15:0] sub_ln703_824_fu_2560_p2;
wire   [15:0] sub_ln703_825_fu_2564_p2;
wire   [15:0] sub_ln703_767_fu_2127_p2;
wire   [15:0] add_ln703_770_fu_2867_p2;
wire   [15:0] add_ln703_742_fu_2569_p2;
wire   [15:0] sub_ln703_793_fu_2356_p2;
wire   [15:0] sub_ln703_826_fu_2574_p2;
wire   [15:0] sub_ln703_827_fu_2579_p2;
wire   [15:0] add_ln703_743_fu_2583_p2;
wire   [15:0] sub_ln703_828_fu_2588_p2;
wire   [15:0] sub_ln703_829_fu_2593_p2;
wire   [15:0] sub_ln703_830_fu_2598_p2;
wire   [15:0] sub_ln703_831_fu_2602_p2;
wire   [15:0] sub_ln703_797_fu_2385_p2;
wire   [15:0] sub_ln703_832_fu_2607_p2;
wire   [15:0] add_ln703_744_fu_2612_p2;
wire   [15:0] sub_ln703_772_fu_2166_p2;
wire   [15:0] add_ln703_776_fu_2937_p2;
wire   [15:0] sub_ln703_773_fu_2171_p2;
wire   [15:0] add_ln703_778_fu_2947_p2;
wire   [15:0] sub_ln703_774_fu_2176_p2;
wire   [15:0] add_ln703_780_fu_2957_p2;
wire   [15:0] add_ln703_745_fu_2617_p2;
wire   [15:0] add_ln703_746_fu_2622_p2;
wire   [15:0] add_ln703_747_fu_2627_p2;
wire   [15:0] add_ln703_748_fu_2632_p2;
wire   [15:0] add_ln703_749_fu_2637_p2;
wire   [15:0] sub_ln703_777_fu_2202_p2;
wire   [15:0] add_ln703_782_fu_2992_p2;
wire   [15:0] sub_ln703_833_fu_2642_p2;
wire   [15:0] sub_ln703_834_fu_2646_p2;
wire   [15:0] sub_ln703_835_fu_2651_p2;
wire   [15:0] sub_ln703_836_fu_2655_p2;
wire   [15:0] sub_ln703_804_fu_2429_p2;
wire   [15:0] add_ln703_786_fu_3027_p2;
wire   [15:0] sub_ln703_837_fu_2660_p2;
wire   [15:0] sub_ln703_838_fu_2664_p2;
wire   [15:0] add_ln703_752_fu_2673_p2;
wire   [15:0] acc_1_V_fu_2678_p2;
wire   [15:0] acc_2_V_fu_2683_p2;
wire   [15:0] acc_3_V_fu_2688_p2;
wire   [15:0] acc_4_V_fu_2698_p2;
wire   [15:0] acc_5_V_fu_2703_p2;
wire   [15:0] acc_6_V_fu_2708_p2;
wire   [15:0] acc_7_V_fu_2713_p2;
wire   [15:0] acc_8_V_fu_2718_p2;
wire   [15:0] acc_9_V_fu_2723_p2;
wire   [15:0] acc_10_V_fu_2733_p2;
wire   [15:0] acc_11_V_fu_2738_p2;
wire   [15:0] acc_12_V_fu_2743_p2;
wire   [15:0] acc_13_V_fu_2748_p2;
wire   [15:0] acc_14_V_fu_2753_p2;
wire   [15:0] acc_15_V_fu_2758_p2;
wire   [15:0] acc_16_V_fu_2771_p2;
wire   [15:0] acc_17_V_fu_2777_p2;
wire   [15:0] acc_18_V_fu_2782_p2;
wire   [15:0] acc_19_V_fu_2787_p2;
wire   [15:0] acc_20_V_fu_2797_p2;
wire   [15:0] acc_21_V_fu_2802_p2;
wire   [15:0] acc_22_V_fu_2807_p2;
wire   [15:0] acc_23_V_fu_2812_p2;
wire   [15:0] acc_24_V_fu_2817_p2;
wire   [15:0] acc_25_V_fu_2822_p2;
wire   [15:0] acc_26_V_fu_2827_p2;
wire   [15:0] acc_27_V_fu_2832_p2;
wire   [15:0] acc_28_V_fu_2837_p2;
wire   [15:0] acc_29_V_fu_2842_p2;
wire   [15:0] acc_30_V_fu_2847_p2;
wire   [15:0] acc_31_V_fu_2852_p2;
wire   [15:0] acc_32_V_fu_2857_p2;
wire   [15:0] acc_33_V_fu_2862_p2;
wire   [15:0] acc_34_V_fu_2872_p2;
wire   [15:0] acc_35_V_fu_2877_p2;
wire   [15:0] acc_36_V_fu_2882_p2;
wire   [15:0] acc_37_V_fu_2887_p2;
wire   [15:0] acc_38_V_fu_2892_p2;
wire   [15:0] acc_39_V_fu_2897_p2;
wire   [15:0] acc_40_V_fu_2902_p2;
wire   [15:0] acc_41_V_fu_2907_p2;
wire   [15:0] acc_42_V_fu_2912_p2;
wire   [15:0] acc_43_V_fu_2917_p2;
wire   [15:0] acc_44_V_fu_2922_p2;
wire   [15:0] acc_45_V_fu_2927_p2;
wire   [15:0] acc_46_V_fu_2932_p2;
wire   [15:0] acc_47_V_fu_2942_p2;
wire   [15:0] acc_48_V_fu_2952_p2;
wire   [15:0] acc_49_V_fu_2962_p2;
wire   [15:0] acc_50_V_fu_2967_p2;
wire   [15:0] acc_51_V_fu_2972_p2;
wire   [15:0] acc_52_V_fu_2977_p2;
wire   [15:0] acc_53_V_fu_2982_p2;
wire   [15:0] acc_54_V_fu_2987_p2;
wire   [15:0] acc_55_V_fu_2997_p2;
wire   [15:0] acc_56_V_fu_3002_p2;
wire   [15:0] acc_57_V_fu_3007_p2;
wire   [15:0] acc_58_V_fu_3012_p2;
wire   [15:0] acc_59_V_fu_3017_p2;
wire   [15:0] acc_60_V_fu_3022_p2;
wire   [15:0] acc_61_V_fu_3031_p2;
wire   [15:0] acc_62_V_fu_3037_p2;
wire   [15:0] acc_63_V_fu_3042_p2;
reg    ap_ce_reg;
reg   [255:0] data_V_read_int_reg;
reg   [15:0] ap_return_0_int_reg;
reg   [15:0] ap_return_1_int_reg;
reg   [15:0] ap_return_2_int_reg;
reg   [15:0] ap_return_3_int_reg;
reg   [15:0] ap_return_4_int_reg;
reg   [15:0] ap_return_5_int_reg;
reg   [15:0] ap_return_6_int_reg;
reg   [15:0] ap_return_7_int_reg;
reg   [15:0] ap_return_8_int_reg;
reg   [15:0] ap_return_9_int_reg;
reg   [15:0] ap_return_10_int_reg;
reg   [15:0] ap_return_11_int_reg;
reg   [15:0] ap_return_12_int_reg;
reg   [15:0] ap_return_13_int_reg;
reg   [15:0] ap_return_14_int_reg;
reg   [15:0] ap_return_15_int_reg;
reg   [15:0] ap_return_16_int_reg;
reg   [15:0] ap_return_17_int_reg;
reg   [15:0] ap_return_18_int_reg;
reg   [15:0] ap_return_19_int_reg;
reg   [15:0] ap_return_20_int_reg;
reg   [15:0] ap_return_21_int_reg;
reg   [15:0] ap_return_22_int_reg;
reg   [15:0] ap_return_23_int_reg;
reg   [15:0] ap_return_24_int_reg;
reg   [15:0] ap_return_25_int_reg;
reg   [15:0] ap_return_26_int_reg;
reg   [15:0] ap_return_27_int_reg;
reg   [15:0] ap_return_28_int_reg;
reg   [15:0] ap_return_29_int_reg;
reg   [15:0] ap_return_30_int_reg;
reg   [15:0] ap_return_31_int_reg;
reg   [15:0] ap_return_32_int_reg;
reg   [15:0] ap_return_33_int_reg;
reg   [15:0] ap_return_34_int_reg;
reg   [15:0] ap_return_35_int_reg;
reg   [15:0] ap_return_36_int_reg;
reg   [15:0] ap_return_37_int_reg;
reg   [15:0] ap_return_38_int_reg;
reg   [15:0] ap_return_39_int_reg;
reg   [15:0] ap_return_40_int_reg;
reg   [15:0] ap_return_41_int_reg;
reg   [15:0] ap_return_42_int_reg;
reg   [15:0] ap_return_43_int_reg;
reg   [15:0] ap_return_44_int_reg;
reg   [15:0] ap_return_45_int_reg;
reg   [15:0] ap_return_46_int_reg;
reg   [15:0] ap_return_47_int_reg;
reg   [15:0] ap_return_48_int_reg;
reg   [15:0] ap_return_49_int_reg;
reg   [15:0] ap_return_50_int_reg;
reg   [15:0] ap_return_51_int_reg;
reg   [15:0] ap_return_52_int_reg;
reg   [15:0] ap_return_53_int_reg;
reg   [15:0] ap_return_54_int_reg;
reg   [15:0] ap_return_55_int_reg;
reg   [15:0] ap_return_56_int_reg;
reg   [15:0] ap_return_57_int_reg;
reg   [15:0] ap_return_58_int_reg;
reg   [15:0] ap_return_59_int_reg;
reg   [15:0] ap_return_60_int_reg;
reg   [15:0] ap_return_61_int_reg;
reg   [15:0] ap_return_62_int_reg;
reg   [15:0] ap_return_63_int_reg;

always @ (posedge ap_clk) begin
    ap_ce_reg <= ap_ce;
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        add_ln703_538_reg_4067 <= add_ln703_538_fu_280_p2;
        add_ln703_538_reg_4067_pp0_iter4_reg <= add_ln703_538_reg_4067;
        add_ln703_539_reg_4035 <= add_ln703_539_fu_260_p2;
        add_ln703_539_reg_4035_pp0_iter2_reg <= add_ln703_539_reg_4035;
        add_ln703_539_reg_4035_pp0_iter3_reg <= add_ln703_539_reg_4035_pp0_iter2_reg;
        add_ln703_540_reg_4079 <= add_ln703_540_fu_288_p2;
        add_ln703_540_reg_4079_pp0_iter4_reg <= add_ln703_540_reg_4079;
        add_ln703_541_reg_4171 <= add_ln703_541_fu_348_p2;
        add_ln703_542_reg_4177 <= add_ln703_542_fu_352_p2;
        add_ln703_543_reg_4054 <= add_ln703_543_fu_272_p2;
        add_ln703_543_reg_4054_pp0_iter3_reg <= add_ln703_543_reg_4054;
        add_ln703_543_reg_4054_pp0_iter4_reg <= add_ln703_543_reg_4054_pp0_iter3_reg;
        add_ln703_544_reg_4116 <= add_ln703_544_fu_312_p2;
        add_ln703_544_reg_4116_pp0_iter5_reg <= add_ln703_544_reg_4116;
        add_ln703_545_reg_4183 <= add_ln703_545_fu_364_p2;
        add_ln703_547_reg_4128 <= add_ln703_547_fu_320_p2;
        add_ln703_548_reg_4188 <= add_ln703_548_fu_368_p2;
        add_ln703_549_reg_4103 <= add_ln703_549_fu_304_p2;
        add_ln703_549_reg_4103_pp0_iter4_reg <= add_ln703_549_reg_4103;
        add_ln703_549_reg_4103_pp0_iter5_reg <= add_ln703_549_reg_4103_pp0_iter4_reg;
        add_ln703_550_reg_4211 <= add_ln703_550_fu_384_p2;
        add_ln703_551_reg_4222 <= add_ln703_551_fu_393_p2;
        add_ln703_554_reg_4134 <= add_ln703_554_fu_324_p2;
        add_ln703_554_reg_4134_pp0_iter5_reg <= add_ln703_554_reg_4134;
        add_ln703_557_reg_4293 <= add_ln703_557_fu_488_p2;
        add_ln703_558_reg_4298 <= add_ln703_558_fu_498_p2;
        add_ln703_559_reg_4146 <= add_ln703_559_fu_332_p2;
        add_ln703_559_reg_4146_pp0_iter5_reg <= add_ln703_559_reg_4146;
        add_ln703_560_reg_4153 <= add_ln703_560_fu_336_p2;
        add_ln703_560_reg_4153_pp0_iter5_reg <= add_ln703_560_reg_4153;
        add_ln703_564_reg_4240 <= add_ln703_564_fu_406_p2;
        add_ln703_566_reg_4258 <= add_ln703_566_fu_418_p2;
        add_ln703_566_reg_4258_pp0_iter6_reg <= add_ln703_566_reg_4258;
        add_ln703_568_reg_4270 <= add_ln703_568_fu_426_p2;
        add_ln703_571_reg_4372 <= add_ln703_571_fu_657_p2;
        add_ln703_572_reg_4382 <= add_ln703_572_fu_670_p2;
        add_ln703_573_reg_4387 <= add_ln703_573_fu_675_p2;
        add_ln703_574_reg_4393 <= add_ln703_574_fu_679_p2;
        add_ln703_576_reg_4408 <= add_ln703_576_fu_702_p2;
        add_ln703_577_reg_4413 <= add_ln703_577_fu_707_p2;
        add_ln703_579_reg_4418 <= add_ln703_579_fu_716_p2;
        add_ln703_580_reg_4433 <= add_ln703_580_fu_730_p2;
        add_ln703_583_reg_4450 <= add_ln703_583_fu_754_p2;
        add_ln703_587_reg_4471 <= add_ln703_587_fu_786_p2;
        add_ln703_588_reg_4476 <= add_ln703_588_fu_792_p2;
        add_ln703_590_reg_4481 <= add_ln703_590_fu_801_p2;
        add_ln703_597_reg_4282 <= add_ln703_597_fu_434_p2;
        add_ln703_597_reg_4282_pp0_iter6_reg <= add_ln703_597_reg_4282;
        add_ln703_611_reg_4521 <= add_ln703_611_fu_887_p2;
        add_ln703_620_reg_4537 <= add_ln703_620_fu_891_p2;
        add_ln703_631_reg_4588 <= add_ln703_631_fu_1397_p2;
        add_ln703_634_reg_4593 <= add_ln703_634_fu_1416_p2;
        add_ln703_637_reg_4553 <= add_ln703_637_fu_906_p2;
        add_ln703_639_reg_4608 <= add_ln703_639_fu_1459_p2;
        add_ln703_642_reg_4628 <= add_ln703_642_fu_1505_p2;
        add_ln703_645_reg_4648 <= add_ln703_645_fu_1538_p2;
        add_ln703_646_reg_4658 <= add_ln703_646_fu_1553_p2;
        add_ln703_655_reg_4558 <= add_ln703_655_fu_910_p2;
        add_ln703_658_reg_4733 <= add_ln703_658_fu_1696_p2;
        add_ln703_659_reg_4568 <= add_ln703_659_fu_914_p2;
        add_ln703_661_reg_4744 <= add_ln703_661_fu_1710_p2;
        add_ln703_663_reg_4764 <= add_ln703_663_fu_1735_p2;
        add_ln703_667_reg_4784 <= add_ln703_667_fu_1767_p2;
        add_ln703_669_reg_4804 <= add_ln703_669_fu_1787_p2;
        add_ln703_670_reg_4819 <= add_ln703_670_fu_1802_p2;
        add_ln703_672_reg_4829 <= add_ln703_672_fu_1812_p2;
        add_ln703_674_reg_4839 <= add_ln703_674_fu_1822_p2;
        add_ln703_679_reg_4847 <= add_ln703_679_fu_1826_p2;
        add_ln703_687_reg_4857 <= add_ln703_687_fu_1847_p2;
        add_ln703_688_reg_4862 <= add_ln703_688_fu_1853_p2;
        add_ln703_692_reg_4573 <= add_ln703_692_fu_920_p2;
        add_ln703_692_reg_4573_pp0_iter7_reg <= add_ln703_692_reg_4573;
        add_ln703_707_reg_4867 <= add_ln703_707_fu_1877_p2;
        add_ln703_711_reg_4872 <= add_ln703_711_fu_1887_p2;
        add_ln703_716_reg_4877 <= add_ln703_716_fu_1902_p2;
        add_ln703_722_reg_4882 <= add_ln703_722_fu_1913_p2;
        add_ln703_724_reg_4887 <= add_ln703_724_fu_1923_p2;
        add_ln703_727_reg_4892 <= add_ln703_727_fu_1934_p2;
        add_ln703_729_reg_4897 <= add_ln703_729_fu_1945_p2;
        add_ln703_732_reg_4902 <= add_ln703_732_fu_1956_p2;
        add_ln703_737_reg_4907 <= add_ln703_737_fu_1962_p2;
        add_ln703_739_reg_4915 <= add_ln703_739_fu_1966_p2;
        add_ln703_751_reg_4920 <= add_ln703_751_fu_1971_p2;
        add_ln703_reg_4010 <= add_ln703_fu_242_p2;
        add_ln703_reg_4010_pp0_iter1_reg <= add_ln703_reg_4010;
        add_ln703_reg_4010_pp0_iter2_reg <= add_ln703_reg_4010_pp0_iter1_reg;
        mult_307_V_reg_3472 <= {{data_V_read_int_reg[79:64]}};
        mult_307_V_reg_3472_pp0_iter1_reg <= mult_307_V_reg_3472;
        mult_307_V_reg_3472_pp0_iter2_reg <= mult_307_V_reg_3472_pp0_iter1_reg;
        mult_307_V_reg_3472_pp0_iter3_reg <= mult_307_V_reg_3472_pp0_iter2_reg;
        mult_307_V_reg_3472_pp0_iter4_reg <= mult_307_V_reg_3472_pp0_iter3_reg;
        mult_307_V_reg_3472_pp0_iter5_reg <= mult_307_V_reg_3472_pp0_iter4_reg;
        mult_320_V_reg_3500 <= {{data_V_read_int_reg[95:80]}};
        mult_320_V_reg_3500_pp0_iter1_reg <= mult_320_V_reg_3500;
        mult_320_V_reg_3500_pp0_iter2_reg <= mult_320_V_reg_3500_pp0_iter1_reg;
        mult_320_V_reg_3500_pp0_iter3_reg <= mult_320_V_reg_3500_pp0_iter2_reg;
        mult_320_V_reg_3500_pp0_iter4_reg <= mult_320_V_reg_3500_pp0_iter3_reg;
        mult_320_V_reg_3500_pp0_iter5_reg <= mult_320_V_reg_3500_pp0_iter4_reg;
        mult_386_V_reg_3539 <= {{data_V_read_int_reg[111:96]}};
        mult_386_V_reg_3539_pp0_iter1_reg <= mult_386_V_reg_3539;
        mult_386_V_reg_3539_pp0_iter2_reg <= mult_386_V_reg_3539_pp0_iter1_reg;
        mult_386_V_reg_3539_pp0_iter3_reg <= mult_386_V_reg_3539_pp0_iter2_reg;
        mult_386_V_reg_3539_pp0_iter4_reg <= mult_386_V_reg_3539_pp0_iter3_reg;
        mult_386_V_reg_3539_pp0_iter5_reg <= mult_386_V_reg_3539_pp0_iter4_reg;
        mult_386_V_reg_3539_pp0_iter6_reg <= mult_386_V_reg_3539_pp0_iter5_reg;
        mult_449_V_reg_3582 <= {{data_V_read_int_reg[127:112]}};
        mult_449_V_reg_3582_pp0_iter1_reg <= mult_449_V_reg_3582;
        mult_449_V_reg_3582_pp0_iter2_reg <= mult_449_V_reg_3582_pp0_iter1_reg;
        mult_449_V_reg_3582_pp0_iter3_reg <= mult_449_V_reg_3582_pp0_iter2_reg;
        mult_449_V_reg_3582_pp0_iter4_reg <= mult_449_V_reg_3582_pp0_iter3_reg;
        mult_449_V_reg_3582_pp0_iter5_reg <= mult_449_V_reg_3582_pp0_iter4_reg;
        mult_449_V_reg_3582_pp0_iter6_reg <= mult_449_V_reg_3582_pp0_iter5_reg;
        mult_512_V_reg_3629 <= {{data_V_read_int_reg[143:128]}};
        mult_512_V_reg_3629_pp0_iter1_reg <= mult_512_V_reg_3629;
        mult_512_V_reg_3629_pp0_iter2_reg <= mult_512_V_reg_3629_pp0_iter1_reg;
        mult_512_V_reg_3629_pp0_iter3_reg <= mult_512_V_reg_3629_pp0_iter2_reg;
        mult_512_V_reg_3629_pp0_iter4_reg <= mult_512_V_reg_3629_pp0_iter3_reg;
        mult_512_V_reg_3629_pp0_iter5_reg <= mult_512_V_reg_3629_pp0_iter4_reg;
        mult_512_V_reg_3629_pp0_iter6_reg <= mult_512_V_reg_3629_pp0_iter5_reg;
        mult_576_V_reg_3674 <= {{data_V_read_int_reg[159:144]}};
        mult_576_V_reg_3674_pp0_iter1_reg <= mult_576_V_reg_3674;
        mult_576_V_reg_3674_pp0_iter2_reg <= mult_576_V_reg_3674_pp0_iter1_reg;
        mult_576_V_reg_3674_pp0_iter3_reg <= mult_576_V_reg_3674_pp0_iter2_reg;
        mult_576_V_reg_3674_pp0_iter4_reg <= mult_576_V_reg_3674_pp0_iter3_reg;
        mult_576_V_reg_3674_pp0_iter5_reg <= mult_576_V_reg_3674_pp0_iter4_reg;
        mult_576_V_reg_3674_pp0_iter6_reg <= mult_576_V_reg_3674_pp0_iter5_reg;
        mult_640_V_reg_3716 <= {{data_V_read_int_reg[175:160]}};
        mult_640_V_reg_3716_pp0_iter1_reg <= mult_640_V_reg_3716;
        mult_640_V_reg_3716_pp0_iter2_reg <= mult_640_V_reg_3716_pp0_iter1_reg;
        mult_640_V_reg_3716_pp0_iter3_reg <= mult_640_V_reg_3716_pp0_iter2_reg;
        mult_640_V_reg_3716_pp0_iter4_reg <= mult_640_V_reg_3716_pp0_iter3_reg;
        mult_640_V_reg_3716_pp0_iter5_reg <= mult_640_V_reg_3716_pp0_iter4_reg;
        mult_640_V_reg_3716_pp0_iter6_reg <= mult_640_V_reg_3716_pp0_iter5_reg;
        mult_704_V_reg_3765 <= {{data_V_read_int_reg[191:176]}};
        mult_704_V_reg_3765_pp0_iter1_reg <= mult_704_V_reg_3765;
        mult_704_V_reg_3765_pp0_iter2_reg <= mult_704_V_reg_3765_pp0_iter1_reg;
        mult_704_V_reg_3765_pp0_iter3_reg <= mult_704_V_reg_3765_pp0_iter2_reg;
        mult_704_V_reg_3765_pp0_iter4_reg <= mult_704_V_reg_3765_pp0_iter3_reg;
        mult_704_V_reg_3765_pp0_iter5_reg <= mult_704_V_reg_3765_pp0_iter4_reg;
        mult_704_V_reg_3765_pp0_iter6_reg <= mult_704_V_reg_3765_pp0_iter5_reg;
        mult_704_V_reg_3765_pp0_iter7_reg <= mult_704_V_reg_3765_pp0_iter6_reg;
        mult_770_V_reg_3814 <= {{data_V_read_int_reg[207:192]}};
        mult_770_V_reg_3814_pp0_iter1_reg <= mult_770_V_reg_3814;
        mult_770_V_reg_3814_pp0_iter2_reg <= mult_770_V_reg_3814_pp0_iter1_reg;
        mult_770_V_reg_3814_pp0_iter3_reg <= mult_770_V_reg_3814_pp0_iter2_reg;
        mult_770_V_reg_3814_pp0_iter4_reg <= mult_770_V_reg_3814_pp0_iter3_reg;
        mult_770_V_reg_3814_pp0_iter5_reg <= mult_770_V_reg_3814_pp0_iter4_reg;
        mult_770_V_reg_3814_pp0_iter6_reg <= mult_770_V_reg_3814_pp0_iter5_reg;
        mult_770_V_reg_3814_pp0_iter7_reg <= mult_770_V_reg_3814_pp0_iter6_reg;
        mult_832_V_reg_3861 <= {{data_V_read_int_reg[223:208]}};
        mult_832_V_reg_3861_pp0_iter1_reg <= mult_832_V_reg_3861;
        mult_832_V_reg_3861_pp0_iter2_reg <= mult_832_V_reg_3861_pp0_iter1_reg;
        mult_832_V_reg_3861_pp0_iter3_reg <= mult_832_V_reg_3861_pp0_iter2_reg;
        mult_832_V_reg_3861_pp0_iter4_reg <= mult_832_V_reg_3861_pp0_iter3_reg;
        mult_832_V_reg_3861_pp0_iter5_reg <= mult_832_V_reg_3861_pp0_iter4_reg;
        mult_832_V_reg_3861_pp0_iter6_reg <= mult_832_V_reg_3861_pp0_iter5_reg;
        mult_832_V_reg_3861_pp0_iter7_reg <= mult_832_V_reg_3861_pp0_iter6_reg;
        mult_896_V_reg_3909 <= {{data_V_read_int_reg[239:224]}};
        mult_896_V_reg_3909_pp0_iter1_reg <= mult_896_V_reg_3909;
        mult_896_V_reg_3909_pp0_iter2_reg <= mult_896_V_reg_3909_pp0_iter1_reg;
        mult_896_V_reg_3909_pp0_iter3_reg <= mult_896_V_reg_3909_pp0_iter2_reg;
        mult_896_V_reg_3909_pp0_iter4_reg <= mult_896_V_reg_3909_pp0_iter3_reg;
        mult_896_V_reg_3909_pp0_iter5_reg <= mult_896_V_reg_3909_pp0_iter4_reg;
        mult_896_V_reg_3909_pp0_iter6_reg <= mult_896_V_reg_3909_pp0_iter5_reg;
        mult_896_V_reg_3909_pp0_iter7_reg <= mult_896_V_reg_3909_pp0_iter6_reg;
        mult_960_V_reg_3958 <= {{data_V_read_int_reg[255:240]}};
        mult_960_V_reg_3958_pp0_iter1_reg <= mult_960_V_reg_3958;
        mult_960_V_reg_3958_pp0_iter2_reg <= mult_960_V_reg_3958_pp0_iter1_reg;
        mult_960_V_reg_3958_pp0_iter3_reg <= mult_960_V_reg_3958_pp0_iter2_reg;
        mult_960_V_reg_3958_pp0_iter4_reg <= mult_960_V_reg_3958_pp0_iter3_reg;
        mult_960_V_reg_3958_pp0_iter5_reg <= mult_960_V_reg_3958_pp0_iter4_reg;
        mult_960_V_reg_3958_pp0_iter6_reg <= mult_960_V_reg_3958_pp0_iter5_reg;
        mult_960_V_reg_3958_pp0_iter7_reg <= mult_960_V_reg_3958_pp0_iter6_reg;
        sub_ln703_531_reg_4023 <= sub_ln703_531_fu_252_p2;
        sub_ln703_531_reg_4023_pp0_iter2_reg <= sub_ln703_531_reg_4023;
        sub_ln703_532_reg_4061 <= sub_ln703_532_fu_276_p2;
        sub_ln703_532_reg_4061_pp0_iter4_reg <= sub_ln703_532_reg_4061;
        sub_ln703_533_reg_4042 <= sub_ln703_533_fu_264_p2;
        sub_ln703_533_reg_4042_pp0_iter3_reg <= sub_ln703_533_reg_4042;
        sub_ln703_533_reg_4042_pp0_iter4_reg <= sub_ln703_533_reg_4042_pp0_iter3_reg;
        sub_ln703_534_reg_4029 <= sub_ln703_534_fu_256_p2;
        sub_ln703_534_reg_4029_pp0_iter2_reg <= sub_ln703_534_reg_4029;
        sub_ln703_534_reg_4029_pp0_iter3_reg <= sub_ln703_534_reg_4029_pp0_iter2_reg;
        sub_ln703_534_reg_4029_pp0_iter4_reg <= sub_ln703_534_reg_4029_pp0_iter3_reg;
        sub_ln703_535_reg_4073 <= sub_ln703_535_fu_284_p2;
        sub_ln703_535_reg_4073_pp0_iter4_reg <= sub_ln703_535_reg_4073;
        sub_ln703_536_reg_4159 <= sub_ln703_536_fu_340_p2;
        sub_ln703_537_reg_4085 <= sub_ln703_537_fu_292_p2;
        sub_ln703_537_reg_4085_pp0_iter4_reg <= sub_ln703_537_reg_4085;
        sub_ln703_537_reg_4085_pp0_iter5_reg <= sub_ln703_537_reg_4085_pp0_iter4_reg;
        sub_ln703_538_reg_4048 <= sub_ln703_538_fu_268_p2;
        sub_ln703_538_reg_4048_pp0_iter3_reg <= sub_ln703_538_reg_4048;
        sub_ln703_538_reg_4048_pp0_iter4_reg <= sub_ln703_538_reg_4048_pp0_iter3_reg;
        sub_ln703_538_reg_4048_pp0_iter5_reg <= sub_ln703_538_reg_4048_pp0_iter4_reg;
        sub_ln703_539_reg_4165 <= sub_ln703_539_fu_344_p2;
        sub_ln703_540_reg_4110 <= sub_ln703_540_fu_308_p2;
        sub_ln703_540_reg_4110_pp0_iter5_reg <= sub_ln703_540_reg_4110;
        sub_ln703_543_reg_4091 <= sub_ln703_543_fu_296_p2;
        sub_ln703_543_reg_4091_pp0_iter4_reg <= sub_ln703_543_reg_4091;
        sub_ln703_544_reg_4122 <= sub_ln703_544_fu_316_p2;
        sub_ln703_544_reg_4122_pp0_iter5_reg <= sub_ln703_544_reg_4122;
        sub_ln703_545_reg_4097 <= sub_ln703_545_fu_300_p2;
        sub_ln703_545_reg_4097_pp0_iter4_reg <= sub_ln703_545_reg_4097;
        sub_ln703_545_reg_4097_pp0_iter5_reg <= sub_ln703_545_reg_4097_pp0_iter4_reg;
        sub_ln703_549_reg_4194 <= sub_ln703_549_fu_372_p2;
        sub_ln703_550_reg_4200 <= sub_ln703_550_fu_376_p2;
        sub_ln703_551_reg_4205 <= sub_ln703_551_fu_380_p2;
        sub_ln703_552_reg_4217 <= sub_ln703_552_fu_388_p2;
        sub_ln703_554_reg_4228 <= sub_ln703_554_fu_398_p2;
        sub_ln703_557_reg_4234 <= sub_ln703_557_fu_402_p2;
        sub_ln703_558_reg_4140 <= sub_ln703_558_fu_328_p2;
        sub_ln703_558_reg_4140_pp0_iter5_reg <= sub_ln703_558_reg_4140;
        sub_ln703_567_reg_4303 <= sub_ln703_567_fu_540_p2;
        sub_ln703_570_reg_4246 <= sub_ln703_570_fu_410_p2;
        sub_ln703_572_reg_4309 <= sub_ln703_572_fu_563_p2;
        sub_ln703_574_reg_4314 <= sub_ln703_574_fu_572_p2;
        sub_ln703_576_reg_4252 <= sub_ln703_576_fu_414_p2;
        sub_ln703_576_reg_4252_pp0_iter6_reg <= sub_ln703_576_reg_4252;
        sub_ln703_578_reg_4319 <= sub_ln703_578_fu_585_p2;
        sub_ln703_579_reg_4324 <= sub_ln703_579_fu_590_p2;
        sub_ln703_582_reg_4329 <= sub_ln703_582_fu_599_p2;
        sub_ln703_584_reg_4264 <= sub_ln703_584_fu_422_p2;
        sub_ln703_584_reg_4264_pp0_iter6_reg <= sub_ln703_584_reg_4264;
        sub_ln703_585_reg_4334 <= sub_ln703_585_fu_609_p2;
        sub_ln703_586_reg_4340 <= sub_ln703_586_fu_614_p2;
        sub_ln703_587_reg_4345 <= sub_ln703_587_fu_619_p2;
        sub_ln703_588_reg_4350 <= sub_ln703_588_fu_624_p2;
        sub_ln703_589_reg_4355 <= sub_ln703_589_fu_638_p2;
        sub_ln703_590_reg_4361 <= sub_ln703_590_fu_643_p2;
        sub_ln703_591_reg_4277 <= sub_ln703_591_fu_430_p2;
        sub_ln703_592_reg_4366 <= sub_ln703_592_fu_653_p2;
        sub_ln703_594_reg_4377 <= sub_ln703_594_fu_666_p2;
        sub_ln703_596_reg_4398 <= sub_ln703_596_fu_683_p2;
        sub_ln703_599_reg_4403 <= sub_ln703_599_fu_693_p2;
        sub_ln703_605_reg_4423 <= sub_ln703_605_fu_720_p2;
        sub_ln703_608_reg_4428 <= sub_ln703_608_fu_725_p2;
        sub_ln703_610_reg_4439 <= sub_ln703_610_fu_734_p2;
        sub_ln703_611_reg_4444 <= sub_ln703_611_fu_739_p2;
        sub_ln703_613_reg_4455 <= sub_ln703_613_fu_758_p2;
        sub_ln703_617_reg_4460 <= sub_ln703_617_fu_763_p2;
        sub_ln703_620_reg_4466 <= sub_ln703_620_fu_772_p2;
        sub_ln703_627_reg_4486 <= sub_ln703_627_fu_807_p2;
        sub_ln703_632_reg_4491 <= sub_ln703_632_fu_818_p2;
        sub_ln703_641_reg_4496 <= sub_ln703_641_fu_838_p2;
        sub_ln703_645_reg_4501 <= sub_ln703_645_fu_843_p2;
        sub_ln703_660_reg_4506 <= sub_ln703_660_fu_872_p2;
        sub_ln703_661_reg_4511 <= sub_ln703_661_fu_877_p2;
        sub_ln703_662_reg_4516 <= sub_ln703_662_fu_882_p2;
        sub_ln703_671_reg_4543 <= sub_ln703_671_fu_896_p2;
        sub_ln703_676_reg_4548 <= sub_ln703_676_fu_901_p2;
        sub_ln703_692_reg_4598 <= sub_ln703_692_fu_1433_p2;
        sub_ln703_693_reg_4603 <= sub_ln703_693_fu_1438_p2;
        sub_ln703_695_reg_4613 <= sub_ln703_695_fu_1464_p2;
        sub_ln703_699_reg_4618 <= sub_ln703_699_fu_1495_p2;
        sub_ln703_700_reg_4623 <= sub_ln703_700_fu_1500_p2;
        sub_ln703_701_reg_4633 <= sub_ln703_701_fu_1509_p2;
        sub_ln703_702_reg_4638 <= sub_ln703_702_fu_1514_p2;
        sub_ln703_704_reg_4643 <= sub_ln703_704_fu_1524_p2;
        sub_ln703_706_reg_4653 <= sub_ln703_706_fu_1548_p2;
        sub_ln703_707_reg_4663 <= sub_ln703_707_fu_1559_p2;
        sub_ln703_708_reg_4668 <= sub_ln703_708_fu_1564_p2;
        sub_ln703_709_reg_4673 <= sub_ln703_709_fu_1569_p2;
        sub_ln703_710_reg_4678 <= sub_ln703_710_fu_1606_p2;
        sub_ln703_711_reg_4683 <= sub_ln703_711_fu_1611_p2;
        sub_ln703_712_reg_4688 <= sub_ln703_712_fu_1616_p2;
        sub_ln703_714_reg_4693 <= sub_ln703_714_fu_1626_p2;
        sub_ln703_715_reg_4698 <= sub_ln703_715_fu_1631_p2;
        sub_ln703_716_reg_4703 <= sub_ln703_716_fu_1636_p2;
        sub_ln703_718_reg_4708 <= sub_ln703_718_fu_1646_p2;
        sub_ln703_720_reg_4713 <= sub_ln703_720_fu_1676_p2;
        sub_ln703_722_reg_4718 <= sub_ln703_722_fu_1681_p2;
        sub_ln703_724_reg_4723 <= sub_ln703_724_fu_1686_p2;
        sub_ln703_725_reg_4728 <= sub_ln703_725_fu_1691_p2;
        sub_ln703_727_reg_4738 <= sub_ln703_727_fu_1701_p2;
        sub_ln703_729_reg_4749 <= sub_ln703_729_fu_1715_p2;
        sub_ln703_730_reg_4754 <= sub_ln703_730_fu_1720_p2;
        sub_ln703_731_reg_4759 <= sub_ln703_731_fu_1725_p2;
        sub_ln703_732_reg_4769 <= sub_ln703_732_fu_1741_p2;
        sub_ln703_738_reg_4774 <= sub_ln703_738_fu_1757_p2;
        sub_ln703_742_reg_4779 <= sub_ln703_742_fu_1762_p2;
        sub_ln703_743_reg_4789 <= sub_ln703_743_fu_1772_p2;
        sub_ln703_744_reg_4794 <= sub_ln703_744_fu_1777_p2;
        sub_ln703_745_reg_4799 <= sub_ln703_745_fu_1782_p2;
        sub_ln703_748_reg_4809 <= sub_ln703_748_fu_1792_p2;
        sub_ln703_751_reg_4814 <= sub_ln703_751_fu_1797_p2;
        sub_ln703_752_reg_4824 <= sub_ln703_752_fu_1807_p2;
        sub_ln703_753_reg_4834 <= sub_ln703_753_fu_1817_p2;
        sub_ln703_765_reg_4852 <= sub_ln703_765_fu_1832_p2;
        sub_ln703_reg_4017 <= sub_ln703_fu_248_p2;
        sub_ln703_reg_4017_pp0_iter2_reg <= sub_ln703_reg_4017;
        tmp_2_reg_3437 <= {{data_V_read_int_reg[31:16]}};
        tmp_3_reg_3443 <= {{data_V_read_int_reg[47:32]}};
        tmp_3_reg_3443_pp0_iter1_reg <= tmp_3_reg_3443;
        tmp_3_reg_3443_pp0_iter2_reg <= tmp_3_reg_3443_pp0_iter1_reg;
        tmp_4_reg_3454 <= {{data_V_read_int_reg[63:48]}};
        tmp_4_reg_3454_pp0_iter1_reg <= tmp_4_reg_3454;
        tmp_4_reg_3454_pp0_iter2_reg <= tmp_4_reg_3454_pp0_iter1_reg;
        tmp_4_reg_3454_pp0_iter3_reg <= tmp_4_reg_3454_pp0_iter2_reg;
        tmp_4_reg_3454_pp0_iter4_reg <= tmp_4_reg_3454_pp0_iter3_reg;
        trunc_ln203_reg_3431 <= trunc_ln203_fu_88_p1;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_ce_reg)) begin
        ap_return_0_int_reg <= add_ln703_752_fu_2673_p2;
        ap_return_10_int_reg <= acc_10_V_fu_2733_p2;
        ap_return_11_int_reg <= acc_11_V_fu_2738_p2;
        ap_return_12_int_reg <= acc_12_V_fu_2743_p2;
        ap_return_13_int_reg <= acc_13_V_fu_2748_p2;
        ap_return_14_int_reg <= acc_14_V_fu_2753_p2;
        ap_return_15_int_reg <= acc_15_V_fu_2758_p2;
        ap_return_16_int_reg <= acc_16_V_fu_2771_p2;
        ap_return_17_int_reg <= acc_17_V_fu_2777_p2;
        ap_return_18_int_reg <= acc_18_V_fu_2782_p2;
        ap_return_19_int_reg <= acc_19_V_fu_2787_p2;
        ap_return_1_int_reg <= acc_1_V_fu_2678_p2;
        ap_return_20_int_reg <= acc_20_V_fu_2797_p2;
        ap_return_21_int_reg <= acc_21_V_fu_2802_p2;
        ap_return_22_int_reg <= acc_22_V_fu_2807_p2;
        ap_return_23_int_reg <= acc_23_V_fu_2812_p2;
        ap_return_24_int_reg <= acc_24_V_fu_2817_p2;
        ap_return_25_int_reg <= acc_25_V_fu_2822_p2;
        ap_return_26_int_reg <= acc_26_V_fu_2827_p2;
        ap_return_27_int_reg <= acc_27_V_fu_2832_p2;
        ap_return_28_int_reg <= acc_28_V_fu_2837_p2;
        ap_return_29_int_reg <= acc_29_V_fu_2842_p2;
        ap_return_2_int_reg <= acc_2_V_fu_2683_p2;
        ap_return_30_int_reg <= acc_30_V_fu_2847_p2;
        ap_return_31_int_reg <= acc_31_V_fu_2852_p2;
        ap_return_32_int_reg <= acc_32_V_fu_2857_p2;
        ap_return_33_int_reg <= acc_33_V_fu_2862_p2;
        ap_return_34_int_reg <= acc_34_V_fu_2872_p2;
        ap_return_35_int_reg <= acc_35_V_fu_2877_p2;
        ap_return_36_int_reg <= acc_36_V_fu_2882_p2;
        ap_return_37_int_reg <= acc_37_V_fu_2887_p2;
        ap_return_38_int_reg <= acc_38_V_fu_2892_p2;
        ap_return_39_int_reg <= acc_39_V_fu_2897_p2;
        ap_return_3_int_reg <= acc_3_V_fu_2688_p2;
        ap_return_40_int_reg <= acc_40_V_fu_2902_p2;
        ap_return_41_int_reg <= acc_41_V_fu_2907_p2;
        ap_return_42_int_reg <= acc_42_V_fu_2912_p2;
        ap_return_43_int_reg <= acc_43_V_fu_2917_p2;
        ap_return_44_int_reg <= acc_44_V_fu_2922_p2;
        ap_return_45_int_reg <= acc_45_V_fu_2927_p2;
        ap_return_46_int_reg <= acc_46_V_fu_2932_p2;
        ap_return_47_int_reg <= acc_47_V_fu_2942_p2;
        ap_return_48_int_reg <= acc_48_V_fu_2952_p2;
        ap_return_49_int_reg <= acc_49_V_fu_2962_p2;
        ap_return_4_int_reg <= acc_4_V_fu_2698_p2;
        ap_return_50_int_reg <= acc_50_V_fu_2967_p2;
        ap_return_51_int_reg <= acc_51_V_fu_2972_p2;
        ap_return_52_int_reg <= acc_52_V_fu_2977_p2;
        ap_return_53_int_reg <= acc_53_V_fu_2982_p2;
        ap_return_54_int_reg <= acc_54_V_fu_2987_p2;
        ap_return_55_int_reg <= acc_55_V_fu_2997_p2;
        ap_return_56_int_reg <= acc_56_V_fu_3002_p2;
        ap_return_57_int_reg <= acc_57_V_fu_3007_p2;
        ap_return_58_int_reg <= acc_58_V_fu_3012_p2;
        ap_return_59_int_reg <= acc_59_V_fu_3017_p2;
        ap_return_5_int_reg <= acc_5_V_fu_2703_p2;
        ap_return_60_int_reg <= acc_60_V_fu_3022_p2;
        ap_return_61_int_reg <= acc_61_V_fu_3031_p2;
        ap_return_62_int_reg <= acc_62_V_fu_3037_p2;
        ap_return_63_int_reg <= acc_63_V_fu_3042_p2;
        ap_return_6_int_reg <= acc_6_V_fu_2708_p2;
        ap_return_7_int_reg <= acc_7_V_fu_2713_p2;
        ap_return_8_int_reg <= acc_8_V_fu_2718_p2;
        ap_return_9_int_reg <= acc_9_V_fu_2723_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_ce)) begin
        data_V_read_int_reg <= data_V_read;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_0 = ap_return_0_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_0 = add_ln703_752_fu_2673_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_1 = ap_return_1_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_1 = acc_1_V_fu_2678_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_10 = ap_return_10_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_10 = acc_10_V_fu_2733_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_11 = ap_return_11_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_11 = acc_11_V_fu_2738_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_12 = ap_return_12_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_12 = acc_12_V_fu_2743_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_13 = ap_return_13_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_13 = acc_13_V_fu_2748_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_14 = ap_return_14_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_14 = acc_14_V_fu_2753_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_15 = ap_return_15_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_15 = acc_15_V_fu_2758_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_16 = ap_return_16_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_16 = acc_16_V_fu_2771_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_17 = ap_return_17_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_17 = acc_17_V_fu_2777_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_18 = ap_return_18_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_18 = acc_18_V_fu_2782_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_19 = ap_return_19_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_19 = acc_19_V_fu_2787_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_2 = ap_return_2_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_2 = acc_2_V_fu_2683_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_20 = ap_return_20_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_20 = acc_20_V_fu_2797_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_21 = ap_return_21_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_21 = acc_21_V_fu_2802_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_22 = ap_return_22_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_22 = acc_22_V_fu_2807_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_23 = ap_return_23_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_23 = acc_23_V_fu_2812_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_24 = ap_return_24_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_24 = acc_24_V_fu_2817_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_25 = ap_return_25_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_25 = acc_25_V_fu_2822_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_26 = ap_return_26_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_26 = acc_26_V_fu_2827_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_27 = ap_return_27_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_27 = acc_27_V_fu_2832_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_28 = ap_return_28_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_28 = acc_28_V_fu_2837_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_29 = ap_return_29_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_29 = acc_29_V_fu_2842_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_3 = ap_return_3_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_3 = acc_3_V_fu_2688_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_30 = ap_return_30_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_30 = acc_30_V_fu_2847_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_31 = ap_return_31_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_31 = acc_31_V_fu_2852_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_32 = ap_return_32_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_32 = acc_32_V_fu_2857_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_33 = ap_return_33_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_33 = acc_33_V_fu_2862_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_34 = ap_return_34_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_34 = acc_34_V_fu_2872_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_35 = ap_return_35_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_35 = acc_35_V_fu_2877_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_36 = ap_return_36_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_36 = acc_36_V_fu_2882_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_37 = ap_return_37_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_37 = acc_37_V_fu_2887_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_38 = ap_return_38_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_38 = acc_38_V_fu_2892_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_39 = ap_return_39_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_39 = acc_39_V_fu_2897_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_4 = ap_return_4_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_4 = acc_4_V_fu_2698_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_40 = ap_return_40_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_40 = acc_40_V_fu_2902_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_41 = ap_return_41_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_41 = acc_41_V_fu_2907_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_42 = ap_return_42_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_42 = acc_42_V_fu_2912_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_43 = ap_return_43_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_43 = acc_43_V_fu_2917_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_44 = ap_return_44_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_44 = acc_44_V_fu_2922_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_45 = ap_return_45_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_45 = acc_45_V_fu_2927_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_46 = ap_return_46_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_46 = acc_46_V_fu_2932_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_47 = ap_return_47_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_47 = acc_47_V_fu_2942_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_48 = ap_return_48_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_48 = acc_48_V_fu_2952_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_49 = ap_return_49_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_49 = acc_49_V_fu_2962_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_5 = ap_return_5_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_5 = acc_5_V_fu_2703_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_50 = ap_return_50_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_50 = acc_50_V_fu_2967_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_51 = ap_return_51_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_51 = acc_51_V_fu_2972_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_52 = ap_return_52_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_52 = acc_52_V_fu_2977_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_53 = ap_return_53_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_53 = acc_53_V_fu_2982_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_54 = ap_return_54_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_54 = acc_54_V_fu_2987_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_55 = ap_return_55_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_55 = acc_55_V_fu_2997_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_56 = ap_return_56_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_56 = acc_56_V_fu_3002_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_57 = ap_return_57_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_57 = acc_57_V_fu_3007_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_58 = ap_return_58_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_58 = acc_58_V_fu_3012_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_59 = ap_return_59_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_59 = acc_59_V_fu_3017_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_6 = ap_return_6_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_6 = acc_6_V_fu_2708_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_60 = ap_return_60_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_60 = acc_60_V_fu_3022_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_61 = ap_return_61_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_61 = acc_61_V_fu_3031_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_62 = ap_return_62_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_62 = acc_62_V_fu_3037_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_63 = ap_return_63_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_63 = acc_63_V_fu_3042_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_7 = ap_return_7_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_7 = acc_7_V_fu_2713_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_8 = ap_return_8_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_8 = acc_8_V_fu_2718_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_9 = ap_return_9_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_9 = acc_9_V_fu_2723_p2;
    end
end

assign acc_10_V_fu_2733_p2 = (add_ln703_758_fu_2728_p2 + add_ln703_751_reg_4920);

assign acc_11_V_fu_2738_p2 = (sub_ln703_811_fu_2474_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_12_V_fu_2743_p2 = (mult_960_V_reg_3958_pp0_iter7_reg + sub_ln703_812_fu_2479_p2);

assign acc_13_V_fu_2748_p2 = (add_ln703_735_fu_2484_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_14_V_fu_2753_p2 = (sub_ln703_813_fu_2489_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_15_V_fu_2758_p2 = (sub_ln703_814_fu_2494_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_16_V_fu_2771_p2 = (add_ln703_761_fu_2763_p2 + add_ln703_762_fu_2767_p2);

assign acc_17_V_fu_2777_p2 = (sub_ln703_815_fu_2499_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_18_V_fu_2782_p2 = (add_ln703_736_fu_2504_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_19_V_fu_2787_p2 = (sub_ln703_790_fu_2299_p2 + add_ln703_751_reg_4920);

assign acc_1_V_fu_2678_p2 = (mult_960_V_reg_3958_pp0_iter7_reg + sub_ln703_805_fu_2439_p2);

assign acc_20_V_fu_2797_p2 = (add_ln703_765_fu_2792_p2 + add_ln703_751_reg_4920);

assign acc_21_V_fu_2802_p2 = (sub_ln703_816_fu_2509_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_22_V_fu_2807_p2 = (mult_960_V_reg_3958_pp0_iter7_reg + sub_ln703_817_fu_2514_p2);

assign acc_23_V_fu_2812_p2 = (sub_ln703_818_fu_2519_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_24_V_fu_2817_p2 = (sub_ln703_819_fu_2524_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_25_V_fu_2822_p2 = (sub_ln703_791_fu_2318_p2 + add_ln703_751_reg_4920);

assign acc_26_V_fu_2827_p2 = (add_ln703_738_fu_2528_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_27_V_fu_2832_p2 = (add_ln703_741_fu_2536_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_28_V_fu_2837_p2 = (sub_ln703_820_fu_2541_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_29_V_fu_2842_p2 = (sub_ln703_821_fu_2546_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_2_V_fu_2683_p2 = (sub_ln703_806_fu_2444_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_30_V_fu_2847_p2 = (mult_960_V_reg_3958_pp0_iter7_reg + sub_ln703_822_fu_2550_p2);

assign acc_31_V_fu_2852_p2 = (sub_ln703_823_fu_2555_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_32_V_fu_2857_p2 = (sub_ln703_824_fu_2560_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_33_V_fu_2862_p2 = (sub_ln703_825_fu_2564_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_34_V_fu_2872_p2 = (add_ln703_770_fu_2867_p2 + add_ln703_751_reg_4920);

assign acc_35_V_fu_2877_p2 = (add_ln703_742_fu_2569_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_36_V_fu_2882_p2 = (sub_ln703_793_fu_2356_p2 + add_ln703_751_reg_4920);

assign acc_37_V_fu_2887_p2 = (sub_ln703_826_fu_2574_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_38_V_fu_2892_p2 = (mult_960_V_reg_3958_pp0_iter7_reg + sub_ln703_827_fu_2579_p2);

assign acc_39_V_fu_2897_p2 = (add_ln703_743_fu_2583_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_3_V_fu_2688_p2 = (sub_ln703_807_fu_2449_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_40_V_fu_2902_p2 = (sub_ln703_828_fu_2588_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_41_V_fu_2907_p2 = (sub_ln703_829_fu_2593_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_42_V_fu_2912_p2 = (sub_ln703_830_fu_2598_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_43_V_fu_2917_p2 = (mult_960_V_reg_3958_pp0_iter7_reg + sub_ln703_831_fu_2602_p2);

assign acc_44_V_fu_2922_p2 = (sub_ln703_797_fu_2385_p2 + add_ln703_751_reg_4920);

assign acc_45_V_fu_2927_p2 = (sub_ln703_832_fu_2607_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_46_V_fu_2932_p2 = (add_ln703_744_fu_2612_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_47_V_fu_2942_p2 = (add_ln703_776_fu_2937_p2 + add_ln703_751_reg_4920);

assign acc_48_V_fu_2952_p2 = (add_ln703_778_fu_2947_p2 + add_ln703_751_reg_4920);

assign acc_49_V_fu_2962_p2 = (add_ln703_780_fu_2957_p2 + add_ln703_751_reg_4920);

assign acc_4_V_fu_2698_p2 = (add_ln703_754_fu_2693_p2 + add_ln703_751_reg_4920);

assign acc_50_V_fu_2967_p2 = (add_ln703_745_fu_2617_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_51_V_fu_2972_p2 = (add_ln703_746_fu_2622_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_52_V_fu_2977_p2 = (add_ln703_747_fu_2627_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_53_V_fu_2982_p2 = (add_ln703_748_fu_2632_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_54_V_fu_2987_p2 = (add_ln703_749_fu_2637_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_55_V_fu_2997_p2 = (add_ln703_782_fu_2992_p2 + add_ln703_751_reg_4920);

assign acc_56_V_fu_3002_p2 = (sub_ln703_833_fu_2642_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_57_V_fu_3007_p2 = (mult_960_V_reg_3958_pp0_iter7_reg + sub_ln703_834_fu_2646_p2);

assign acc_58_V_fu_3012_p2 = (sub_ln703_835_fu_2651_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_59_V_fu_3017_p2 = (sub_ln703_836_fu_2655_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_5_V_fu_2703_p2 = (sub_ln703_808_fu_2454_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_60_V_fu_3022_p2 = (sub_ln703_804_fu_2429_p2 + add_ln703_751_reg_4920);

assign acc_61_V_fu_3031_p2 = (add_ln703_786_fu_3027_p2 + add_ln703_762_fu_2767_p2);

assign acc_62_V_fu_3037_p2 = (sub_ln703_837_fu_2660_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_63_V_fu_3042_p2 = (sub_ln703_838_fu_2664_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_6_V_fu_2708_p2 = (sub_ln703_809_fu_2459_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign acc_7_V_fu_2713_p2 = (mult_960_V_reg_3958_pp0_iter7_reg + sub_ln703_810_fu_2464_p2);

assign acc_8_V_fu_2718_p2 = (sub_ln703_785_fu_2254_p2 + add_ln703_751_reg_4920);

assign acc_9_V_fu_2723_p2 = (add_ln703_734_fu_2469_p2 - mult_960_V_reg_3958_pp0_iter7_reg);

assign add_ln703_538_fu_280_p2 = (tmp_3_reg_3443_pp0_iter2_reg + sub_ln703_reg_4017_pp0_iter2_reg);

assign add_ln703_539_fu_260_p2 = (tmp_3_reg_3443 + add_ln703_reg_4010);

assign add_ln703_540_fu_288_p2 = (tmp_3_reg_3443_pp0_iter2_reg + sub_ln703_531_reg_4023_pp0_iter2_reg);

assign add_ln703_541_fu_348_p2 = (tmp_4_reg_3454_pp0_iter4_reg + sub_ln703_535_reg_4073_pp0_iter4_reg);

assign add_ln703_542_fu_352_p2 = (tmp_4_reg_3454_pp0_iter4_reg + sub_ln703_534_reg_4029_pp0_iter4_reg);

assign add_ln703_543_fu_272_p2 = (tmp_4_reg_3454_pp0_iter1_reg + add_ln703_539_reg_4035);

assign add_ln703_544_fu_312_p2 = (tmp_4_reg_3454_pp0_iter3_reg + sub_ln703_532_reg_4061);

assign add_ln703_545_fu_364_p2 = (tmp_4_reg_3454_pp0_iter4_reg + sub_ln703_533_reg_4042_pp0_iter4_reg);

assign add_ln703_546_fu_438_p2 = (mult_307_V_reg_3472_pp0_iter5_reg + sub_ln703_536_reg_4159);

assign add_ln703_547_fu_320_p2 = (mult_307_V_reg_3472_pp0_iter3_reg + tmp_4_reg_3454_pp0_iter3_reg);

assign add_ln703_548_fu_368_p2 = (add_ln703_538_reg_4067_pp0_iter4_reg + add_ln703_547_reg_4128);

assign add_ln703_549_fu_304_p2 = (mult_307_V_reg_3472_pp0_iter2_reg + add_ln703_543_reg_4054);

assign add_ln703_550_fu_384_p2 = (add_ln703_540_reg_4079_pp0_iter4_reg + add_ln703_547_reg_4128);

assign add_ln703_551_fu_393_p2 = (mult_307_V_reg_3472_pp0_iter4_reg + sub_ln703_542_fu_360_p2);

assign add_ln703_552_fu_454_p2 = (mult_307_V_reg_3472_pp0_iter5_reg + add_ln703_542_reg_4177);

assign add_ln703_553_fu_458_p2 = (mult_307_V_reg_3472_pp0_iter5_reg + sub_ln703_539_reg_4165);

assign add_ln703_554_fu_324_p2 = (mult_307_V_reg_3472_pp0_iter3_reg + sub_ln703_543_reg_4091);

assign add_ln703_555_fu_466_p2 = (mult_307_V_reg_3472_pp0_iter5_reg + sub_ln703_538_reg_4048_pp0_iter5_reg);

assign add_ln703_556_fu_478_p2 = (mult_320_V_reg_3500_pp0_iter5_reg + add_ln703_546_fu_438_p2);

assign add_ln703_557_fu_488_p2 = (mult_320_V_reg_3500_pp0_iter5_reg + sub_ln703_547_fu_446_p2);

assign add_ln703_558_fu_498_p2 = (mult_320_V_reg_3500_pp0_iter5_reg + add_ln703_548_reg_4188);

assign add_ln703_559_fu_332_p2 = (mult_320_V_reg_3500_pp0_iter3_reg + add_ln703_549_reg_4103);

assign add_ln703_560_fu_336_p2 = (mult_320_V_reg_3500_pp0_iter3_reg + mult_307_V_reg_3472_pp0_iter3_reg);

assign add_ln703_561_fu_510_p2 = (add_ln703_541_reg_4171 + add_ln703_560_reg_4153_pp0_iter5_reg);

assign add_ln703_562_fu_522_p2 = (mult_320_V_reg_3500_pp0_iter5_reg + sub_ln703_552_reg_4217);

assign add_ln703_563_fu_526_p2 = (mult_320_V_reg_3500_pp0_iter5_reg + add_ln703_551_reg_4222);

assign add_ln703_564_fu_406_p2 = (add_ln703_544_reg_4116 + add_ln703_560_reg_4153);

assign add_ln703_565_fu_554_p2 = (mult_320_V_reg_3500_pp0_iter5_reg + sub_ln703_544_reg_4122_pp0_iter5_reg);

assign add_ln703_566_fu_418_p2 = (mult_386_V_reg_3539_pp0_iter4_reg + sub_ln703_558_reg_4140);

assign add_ln703_567_fu_629_p2 = (mult_307_V_reg_3472_pp0_iter5_reg + sub_ln703_537_reg_4085_pp0_iter5_reg);

assign add_ln703_568_fu_426_p2 = (mult_386_V_reg_3539_pp0_iter4_reg + mult_320_V_reg_3500_pp0_iter4_reg);

assign add_ln703_569_fu_633_p2 = (add_ln703_567_fu_629_p2 + add_ln703_568_reg_4270);

assign add_ln703_570_fu_648_p2 = (mult_386_V_reg_3539_pp0_iter5_reg + sub_ln703_566_fu_535_p2);

assign add_ln703_571_fu_657_p2 = (sub_ln703_554_reg_4228 + add_ln703_568_reg_4270);

assign add_ln703_572_fu_670_p2 = (mult_386_V_reg_3539_pp0_iter5_reg + sub_ln703_569_fu_549_p2);

assign add_ln703_573_fu_675_p2 = (mult_386_V_reg_3539_pp0_iter5_reg + add_ln703_559_reg_4146_pp0_iter5_reg);

assign add_ln703_574_fu_679_p2 = (mult_386_V_reg_3539_pp0_iter5_reg + sub_ln703_570_reg_4246);

assign add_ln703_575_fu_698_p2 = (mult_386_V_reg_3539_pp0_iter5_reg + add_ln703_564_reg_4240);

assign add_ln703_576_fu_702_p2 = (mult_386_V_reg_3539_pp0_iter5_reg + sub_ln703_575_fu_577_p2);

assign add_ln703_577_fu_707_p2 = (mult_386_V_reg_3539_pp0_iter5_reg + sub_ln703_577_fu_581_p2);

assign add_ln703_578_fu_944_p2 = (mult_386_V_reg_3539_pp0_iter6_reg + add_ln703_558_reg_4298);

assign add_ln703_579_fu_716_p2 = (mult_386_V_reg_3539_pp0_iter5_reg + sub_ln703_576_reg_4252);

assign add_ln703_580_fu_730_p2 = (mult_449_V_reg_3582_pp0_iter5_reg + sub_ln703_584_reg_4264);

assign add_ln703_581_fu_744_p2 = (mult_449_V_reg_3582_pp0_iter5_reg + mult_386_V_reg_3539_pp0_iter5_reg);

assign add_ln703_582_fu_748_p2 = (sub_ln703_564_fu_518_p2 + add_ln703_581_fu_744_p2);

assign add_ln703_583_fu_754_p2 = (mult_449_V_reg_3582_pp0_iter5_reg + add_ln703_566_reg_4258);

assign add_ln703_584_fu_985_p2 = (mult_449_V_reg_3582_pp0_iter6_reg + sub_ln703_592_reg_4366);

assign add_ln703_585_fu_777_p2 = (mult_307_V_reg_3472_pp0_iter5_reg + sub_ln703_540_reg_4110_pp0_iter5_reg);

assign add_ln703_586_fu_781_p2 = (mult_320_V_reg_3500_pp0_iter5_reg + add_ln703_581_fu_744_p2);

assign add_ln703_587_fu_786_p2 = (add_ln703_585_fu_777_p2 + add_ln703_586_fu_781_p2);

assign add_ln703_588_fu_792_p2 = (mult_449_V_reg_3582_pp0_iter5_reg + sub_ln703_597_fu_688_p2);

assign add_ln703_589_fu_797_p2 = (mult_320_V_reg_3500_pp0_iter5_reg + sub_ln703_545_reg_4097_pp0_iter5_reg);

assign add_ln703_590_fu_801_p2 = (add_ln703_589_fu_797_p2 + add_ln703_581_fu_744_p2);

assign add_ln703_591_fu_1027_p2 = (mult_449_V_reg_3582_pp0_iter6_reg + add_ln703_573_reg_4387);

assign add_ln703_592_fu_1031_p2 = (mult_449_V_reg_3582_pp0_iter6_reg + sub_ln703_589_reg_4355);

assign add_ln703_593_fu_812_p2 = (sub_ln703_568_fu_545_p2 + add_ln703_581_fu_744_p2);

assign add_ln703_594_fu_823_p2 = (sub_ln703_557_reg_4234 + add_ln703_581_fu_744_p2);

assign add_ln703_595_fu_828_p2 = (mult_320_V_reg_3500_pp0_iter5_reg + add_ln703_550_reg_4211);

assign add_ln703_596_fu_832_p2 = (add_ln703_595_fu_828_p2 + add_ln703_581_fu_744_p2);

assign add_ln703_597_fu_434_p2 = (mult_512_V_reg_3629_pp0_iter4_reg + mult_449_V_reg_3582_pp0_iter4_reg);

assign add_ln703_598_fu_1052_p2 = (sub_ln703_579_reg_4324 + add_ln703_597_reg_4282_pp0_iter6_reg);

assign add_ln703_599_fu_1073_p2 = (mult_512_V_reg_3629_pp0_iter6_reg + sub_ln703_609_fu_965_p2);

assign add_ln703_600_fu_848_p2 = (mult_320_V_reg_3500_pp0_iter5_reg + add_ln703_554_reg_4134_pp0_iter5_reg);

assign add_ln703_601_fu_852_p2 = (mult_386_V_reg_3539_pp0_iter5_reg + add_ln703_597_reg_4282);

assign add_ln703_602_fu_856_p2 = (add_ln703_600_fu_848_p2 + add_ln703_601_fu_852_p2);

assign add_ln703_603_fu_1132_p2 = (sub_ln703_596_reg_4398 + add_ln703_597_reg_4282_pp0_iter6_reg);

assign add_ln703_604_fu_1140_p2 = (sub_ln703_598_fu_932_p2 + add_ln703_597_reg_4282_pp0_iter6_reg);

assign add_ln703_605_fu_862_p2 = (mult_320_V_reg_3500_pp0_iter5_reg + sub_ln703_549_reg_4194);

assign add_ln703_606_fu_866_p2 = (add_ln703_605_fu_862_p2 + add_ln703_601_fu_852_p2);

assign add_ln703_607_fu_1163_p2 = (mult_512_V_reg_3629_pp0_iter6_reg + sub_ln703_611_reg_4444);

assign add_ln703_608_fu_1176_p2 = (mult_512_V_reg_3629_pp0_iter6_reg + sub_ln703_631_fu_1039_p2);

assign add_ln703_609_fu_1181_p2 = (mult_512_V_reg_3629_pp0_iter6_reg + sub_ln703_632_reg_4491);

assign add_ln703_610_fu_1185_p2 = (sub_ln703_586_reg_4340 + add_ln703_597_reg_4282_pp0_iter6_reg);

assign add_ln703_611_fu_887_p2 = (mult_576_V_reg_3674_pp0_iter5_reg + mult_512_V_reg_3629_pp0_iter5_reg);

assign add_ln703_612_fu_1194_p2 = (sub_ln703_604_fu_952_p2 + add_ln703_611_reg_4521);

assign add_ln703_613_fu_1209_p2 = (mult_576_V_reg_3674_pp0_iter6_reg + sub_ln703_638_fu_1069_p2);

assign add_ln703_614_fu_1219_p2 = (mult_576_V_reg_3674_pp0_iter6_reg + sub_ln703_639_fu_1078_p2);

assign add_ln703_615_fu_1228_p2 = (mult_576_V_reg_3674_pp0_iter6_reg + sub_ln703_643_fu_1091_p2);

assign add_ln703_616_fu_1238_p2 = (sub_ln703_615_fu_977_p2 + add_ln703_611_reg_4521);

assign add_ln703_617_fu_1243_p2 = (sub_ln703_616_fu_981_p2 + add_ln703_611_reg_4521);

assign add_ln703_618_fu_1248_p2 = (add_ln703_580_reg_4433 + add_ln703_611_reg_4521);

assign add_ln703_619_fu_1252_p2 = (sub_ln703_617_reg_4460 + add_ln703_611_reg_4521);

assign add_ln703_620_fu_891_p2 = (mult_576_V_reg_3674_pp0_iter5_reg + sub_ln703_645_fu_843_p2);

assign add_ln703_621_fu_1256_p2 = (mult_576_V_reg_3674_pp0_iter6_reg + sub_ln703_646_fu_1099_p2);

assign add_ln703_622_fu_1271_p2 = (mult_576_V_reg_3674_pp0_iter6_reg + sub_ln703_648_fu_1108_p2);

assign add_ln703_623_fu_1276_p2 = (mult_576_V_reg_3674_pp0_iter6_reg + sub_ln703_649_fu_1113_p2);

assign add_ln703_624_fu_1286_p2 = (mult_576_V_reg_3674_pp0_iter6_reg + sub_ln703_652_fu_1127_p2);

assign add_ln703_625_fu_1311_p2 = (sub_ln703_629_fu_1022_p2 + add_ln703_611_reg_4521);

assign add_ln703_626_fu_1321_p2 = (mult_449_V_reg_3582_pp0_iter6_reg + sub_ln703_587_reg_4345);

assign add_ln703_627_fu_1325_p2 = (add_ln703_626_fu_1321_p2 + add_ln703_611_reg_4521);

assign add_ln703_628_fu_1350_p2 = (mult_449_V_reg_3582_pp0_iter6_reg + sub_ln703_601_fu_940_p2);

assign add_ln703_629_fu_1355_p2 = (add_ln703_628_fu_1350_p2 + add_ln703_611_reg_4521);

assign add_ln703_630_fu_1387_p2 = (sub_ln703_634_fu_1048_p2 + add_ln703_611_reg_4521);

assign add_ln703_631_fu_1397_p2 = (mult_640_V_reg_3716_pp0_iter6_reg + add_ln703_612_fu_1194_p2);

assign add_ln703_632_fu_1407_p2 = (mult_512_V_reg_3629_pp0_iter6_reg + sub_ln703_606_fu_956_p2);

assign add_ln703_633_fu_1412_p2 = (mult_640_V_reg_3716_pp0_iter6_reg + mult_576_V_reg_3674_pp0_iter6_reg);

assign add_ln703_634_fu_1416_p2 = (add_ln703_632_fu_1407_p2 + add_ln703_633_fu_1412_p2);

assign add_ln703_635_fu_1422_p2 = (sub_ln703_636_fu_1060_p2 + add_ln703_633_fu_1412_p2);

assign add_ln703_636_fu_1448_p2 = (sub_ln703_640_fu_1082_p2 + add_ln703_633_fu_1412_p2);

assign add_ln703_637_fu_906_p2 = (sub_ln703_551_reg_4205 + add_ln703_568_reg_4270);

assign add_ln703_638_fu_1454_p2 = (add_ln703_597_reg_4282_pp0_iter6_reg + add_ln703_633_fu_1412_p2);

assign add_ln703_639_fu_1459_p2 = (add_ln703_637_reg_4553 + add_ln703_638_fu_1454_p2);

assign add_ln703_640_fu_1469_p2 = (sub_ln703_642_fu_1086_p2 + add_ln703_633_fu_1412_p2);

assign add_ln703_641_fu_1480_p2 = (mult_640_V_reg_3716_pp0_iter6_reg + sub_ln703_668_fu_1233_p2);

assign add_ln703_642_fu_1505_p2 = (mult_640_V_reg_3716_pp0_iter6_reg + add_ln703_620_reg_4537);

assign add_ln703_643_fu_1529_p2 = (mult_449_V_reg_3582_pp0_iter6_reg + sub_ln703_585_reg_4334);

assign add_ln703_644_fu_1533_p2 = (mult_512_V_reg_3629_pp0_iter6_reg + add_ln703_633_fu_1412_p2);

assign add_ln703_645_fu_1538_p2 = (add_ln703_643_fu_1529_p2 + add_ln703_644_fu_1533_p2);

assign add_ln703_646_fu_1553_p2 = (sub_ln703_650_fu_1118_p2 + add_ln703_633_fu_1412_p2);

assign add_ln703_647_fu_1574_p2 = (mult_640_V_reg_3716_pp0_iter6_reg + sub_ln703_674_fu_1296_p2);

assign add_ln703_648_fu_1579_p2 = (mult_512_V_reg_3629_pp0_iter6_reg + sub_ln703_626_fu_1014_p2);

assign add_ln703_649_fu_1584_p2 = (add_ln703_648_fu_1579_p2 + add_ln703_633_fu_1412_p2);

assign add_ln703_650_fu_1590_p2 = (mult_640_V_reg_3716_pp0_iter6_reg + sub_ln703_677_fu_1306_p2);

assign add_ln703_651_fu_1595_p2 = (mult_512_V_reg_3629_pp0_iter6_reg + sub_ln703_628_fu_1018_p2);

assign add_ln703_652_fu_1600_p2 = (add_ln703_651_fu_1595_p2 + add_ln703_633_fu_1412_p2);

assign add_ln703_653_fu_1651_p2 = (mult_640_V_reg_3716_pp0_iter6_reg + sub_ln703_687_fu_1378_p2);

assign add_ln703_654_fu_1661_p2 = (mult_512_V_reg_3629_pp0_iter6_reg + sub_ln703_603_fu_948_p2);

assign add_ln703_655_fu_910_p2 = (mult_704_V_reg_3765_pp0_iter5_reg + mult_640_V_reg_3716_pp0_iter5_reg);

assign add_ln703_656_fu_1666_p2 = (mult_576_V_reg_3674_pp0_iter6_reg + add_ln703_655_reg_4558);

assign add_ln703_657_fu_1670_p2 = (add_ln703_654_fu_1661_p2 + add_ln703_656_fu_1666_p2);

assign add_ln703_658_fu_1696_p2 = (mult_704_V_reg_3765_pp0_iter6_reg + sub_ln703_694_fu_1443_p2);

assign add_ln703_659_fu_914_p2 = (sub_ln703_563_fu_514_p2 + add_ln703_581_fu_744_p2);

assign add_ln703_660_fu_1706_p2 = (add_ln703_611_reg_4521 + add_ln703_655_reg_4558);

assign add_ln703_661_fu_1710_p2 = (add_ln703_659_reg_4568 + add_ln703_660_fu_1706_p2);

assign add_ln703_662_fu_1730_p2 = (mult_512_V_reg_3629_pp0_iter6_reg + sub_ln703_614_fu_973_p2);

assign add_ln703_663_fu_1735_p2 = (add_ln703_662_fu_1730_p2 + add_ln703_656_fu_1666_p2);

assign add_ln703_664_fu_1991_p2 = (mult_704_V_reg_3765_pp0_iter7_reg + sub_ln703_699_reg_4618);

assign add_ln703_665_fu_1746_p2 = (mult_512_V_reg_3629_pp0_iter6_reg + sub_ln703_619_fu_989_p2);

assign add_ln703_666_fu_1751_p2 = (add_ln703_665_fu_1746_p2 + add_ln703_656_fu_1666_p2);

assign add_ln703_667_fu_1767_p2 = (sub_ln703_675_fu_1301_p2 + add_ln703_655_reg_4558);

assign add_ln703_668_fu_2035_p2 = (mult_704_V_reg_3765_pp0_iter7_reg + sub_ln703_712_reg_4688);

assign add_ln703_669_fu_1787_p2 = (sub_ln703_680_fu_1335_p2 + add_ln703_655_reg_4558);

assign add_ln703_670_fu_1802_p2 = (sub_ln703_685_fu_1370_p2 + add_ln703_655_reg_4558);

assign add_ln703_671_fu_2047_p2 = (mult_704_V_reg_3765_pp0_iter7_reg + sub_ln703_718_reg_4708);

assign add_ln703_672_fu_1812_p2 = (mult_704_V_reg_3765_pp0_iter6_reg + sub_ln703_719_fu_1656_p2);

assign add_ln703_673_fu_2068_p2 = (mult_770_V_reg_3814_pp0_iter7_reg + sub_ln703_725_reg_4728);

assign add_ln703_674_fu_1822_p2 = (mult_770_V_reg_3814_pp0_iter6_reg + mult_704_V_reg_3765_pp0_iter6_reg);

assign add_ln703_675_fu_2072_p2 = (sub_ln703_692_reg_4598 + add_ln703_674_reg_4839);

assign add_ln703_676_fu_2093_p2 = (sub_ln703_695_reg_4613 + add_ln703_674_reg_4839);

assign add_ln703_677_fu_2101_p2 = (mult_770_V_reg_3814_pp0_iter7_reg + sub_ln703_730_reg_4754);

assign add_ln703_678_fu_2109_p2 = (mult_770_V_reg_3814_pp0_iter7_reg + sub_ln703_732_reg_4769);

assign add_ln703_679_fu_1826_p2 = (sub_ln703_698_fu_1490_p2 + add_ln703_674_fu_1822_p2);

assign add_ln703_680_fu_2118_p2 = (mult_770_V_reg_3814_pp0_iter7_reg + sub_ln703_736_fu_2007_p2);

assign add_ln703_681_fu_2132_p2 = (mult_770_V_reg_3814_pp0_iter7_reg + sub_ln703_727_reg_4738);

assign add_ln703_682_fu_2136_p2 = (mult_770_V_reg_3814_pp0_iter7_reg + sub_ln703_740_fu_2019_p2);

assign add_ln703_683_fu_2146_p2 = (mult_770_V_reg_3814_pp0_iter7_reg + sub_ln703_742_reg_4779);

assign add_ln703_684_fu_2154_p2 = (mult_770_V_reg_3814_pp0_iter7_reg + sub_ln703_743_reg_4789);

assign add_ln703_685_fu_1837_p2 = (mult_576_V_reg_3674_pp0_iter6_reg + sub_ln703_654_fu_1145_p2);

assign add_ln703_686_fu_1842_p2 = (mult_640_V_reg_3716_pp0_iter6_reg + add_ln703_674_fu_1822_p2);

assign add_ln703_687_fu_1847_p2 = (add_ln703_685_fu_1837_p2 + add_ln703_686_fu_1842_p2);

assign add_ln703_688_fu_1853_p2 = (mult_640_V_reg_3716_pp0_iter6_reg + sub_ln703_679_fu_1330_p2);

assign add_ln703_689_fu_2181_p2 = (add_ln703_688_reg_4862 + add_ln703_674_reg_4839);

assign add_ln703_690_fu_2189_p2 = (mult_770_V_reg_3814_pp0_iter7_reg + sub_ln703_748_reg_4809);

assign add_ln703_691_fu_2193_p2 = (sub_ln703_714_reg_4693 + add_ln703_674_reg_4839);

assign add_ln703_692_fu_920_p2 = (mult_832_V_reg_3861_pp0_iter5_reg + mult_770_V_reg_3814_pp0_iter5_reg);

assign add_ln703_693_fu_2229_p2 = (sub_ln703_721_fu_1975_p2 + add_ln703_692_reg_4573_pp0_iter7_reg);

assign add_ln703_694_fu_2234_p2 = (mult_832_V_reg_3861_pp0_iter7_reg + sub_ln703_755_fu_2055_p2);

assign add_ln703_695_fu_2239_p2 = (mult_832_V_reg_3861_pp0_iter7_reg + sub_ln703_757_fu_2064_p2);

assign add_ln703_696_fu_2264_p2 = (sub_ln703_728_fu_1987_p2 + add_ln703_692_reg_4573_pp0_iter7_reg);

assign add_ln703_697_fu_2269_p2 = (mult_832_V_reg_3861_pp0_iter7_reg + sub_ln703_761_fu_2089_p2);

assign add_ln703_698_fu_2279_p2 = (mult_832_V_reg_3861_pp0_iter7_reg + sub_ln703_762_fu_2097_p2);

assign add_ln703_699_fu_2289_p2 = (mult_832_V_reg_3861_pp0_iter7_reg + sub_ln703_763_fu_2105_p2);

assign add_ln703_700_fu_2303_p2 = (sub_ln703_733_fu_1995_p2 + add_ln703_692_reg_4573_pp0_iter7_reg);

assign add_ln703_701_fu_2308_p2 = (sub_ln703_734_fu_1999_p2 + add_ln703_692_reg_4573_pp0_iter7_reg);

assign add_ln703_702_fu_2313_p2 = (sub_ln703_735_fu_2003_p2 + add_ln703_692_reg_4573_pp0_iter7_reg);

assign add_ln703_703_fu_1858_p2 = (mult_386_V_reg_3539_pp0_iter6_reg + sub_ln703_567_reg_4303);

assign add_ln703_704_fu_1862_p2 = (add_ln703_703_fu_1858_p2 + add_ln703_597_reg_4282_pp0_iter6_reg);

assign add_ln703_705_fu_1867_p2 = (mult_704_V_reg_3765_pp0_iter6_reg + add_ln703_692_reg_4573);

assign add_ln703_706_fu_1871_p2 = (add_ln703_633_fu_1412_p2 + add_ln703_705_fu_1867_p2);

assign add_ln703_707_fu_1877_p2 = (add_ln703_704_fu_1862_p2 + add_ln703_706_fu_1871_p2);

assign add_ln703_708_fu_2323_p2 = (mult_704_V_reg_3765_pp0_iter7_reg + sub_ln703_704_reg_4643);

assign add_ln703_709_fu_2327_p2 = (add_ln703_708_fu_2323_p2 + add_ln703_692_reg_4573_pp0_iter7_reg);

assign add_ln703_710_fu_1883_p2 = (mult_640_V_reg_3716_pp0_iter6_reg + sub_ln703_671_reg_4543);

assign add_ln703_711_fu_1887_p2 = (add_ln703_710_fu_1883_p2 + add_ln703_705_fu_1867_p2);

assign add_ln703_712_fu_2332_p2 = (sub_ln703_737_fu_2011_p2 + add_ln703_692_reg_4573_pp0_iter7_reg);

assign add_ln703_713_fu_2337_p2 = (mult_832_V_reg_3861_pp0_iter7_reg + sub_ln703_766_fu_2123_p2);

assign add_ln703_714_fu_1893_p2 = (sub_ln703_622_fu_997_p2 + add_ln703_611_reg_4521);

assign add_ln703_715_fu_1898_p2 = (add_ln703_655_reg_4558 + add_ln703_692_reg_4573);

assign add_ln703_716_fu_1902_p2 = (add_ln703_714_fu_1893_p2 + add_ln703_715_fu_1898_p2);

assign add_ln703_717_fu_2342_p2 = (mult_704_V_reg_3765_pp0_iter7_reg + sub_ln703_706_reg_4653);

assign add_ln703_718_fu_2346_p2 = (add_ln703_717_fu_2342_p2 + add_ln703_692_reg_4573_pp0_iter7_reg);

assign add_ln703_719_fu_2361_p2 = (mult_704_V_reg_3765_pp0_iter7_reg + sub_ln703_708_reg_4668);

assign add_ln703_720_fu_2365_p2 = (add_ln703_719_fu_2361_p2 + add_ln703_692_reg_4573_pp0_iter7_reg);

assign add_ln703_721_fu_1908_p2 = (mult_640_V_reg_3716_pp0_iter6_reg + sub_ln703_673_fu_1291_p2);

assign add_ln703_722_fu_1913_p2 = (add_ln703_721_fu_1908_p2 + add_ln703_705_fu_1867_p2);

assign add_ln703_723_fu_1919_p2 = (mult_640_V_reg_3716_pp0_iter6_reg + sub_ln703_676_reg_4548);

assign add_ln703_724_fu_1923_p2 = (add_ln703_723_fu_1919_p2 + add_ln703_705_fu_1867_p2);

assign add_ln703_725_fu_2389_p2 = (mult_832_V_reg_3861_pp0_iter7_reg + sub_ln703_770_fu_2158_p2);

assign add_ln703_726_fu_1929_p2 = (sub_ln703_660_reg_4506 + add_ln703_633_fu_1412_p2);

assign add_ln703_727_fu_1934_p2 = (add_ln703_726_fu_1929_p2 + add_ln703_705_fu_1867_p2);

assign add_ln703_728_fu_1940_p2 = (sub_ln703_633_fu_1043_p2 + add_ln703_611_reg_4521);

assign add_ln703_729_fu_1945_p2 = (add_ln703_728_fu_1940_p2 + add_ln703_715_fu_1898_p2);

assign add_ln703_730_fu_2424_p2 = (mult_832_V_reg_3861_pp0_iter7_reg + sub_ln703_779_fu_2211_p2);

assign add_ln703_731_fu_1951_p2 = (mult_640_V_reg_3716_pp0_iter6_reg + sub_ln703_688_fu_1382_p2);

assign add_ln703_732_fu_1956_p2 = (add_ln703_731_fu_1951_p2 + add_ln703_705_fu_1867_p2);

assign add_ln703_733_fu_2434_p2 = (mult_832_V_reg_3861_pp0_iter7_reg + sub_ln703_781_fu_2220_p2);

assign add_ln703_734_fu_2469_p2 = (mult_896_V_reg_3909_pp0_iter7_reg + sub_ln703_786_fu_2259_p2);

assign add_ln703_735_fu_2484_p2 = (mult_896_V_reg_3909_pp0_iter7_reg + sub_ln703_787_fu_2274_p2);

assign add_ln703_736_fu_2504_p2 = (mult_896_V_reg_3909_pp0_iter7_reg + sub_ln703_789_fu_2294_p2);

assign add_ln703_737_fu_1962_p2 = (mult_896_V_reg_3909_pp0_iter6_reg + mult_832_V_reg_3861_pp0_iter6_reg);

assign add_ln703_738_fu_2528_p2 = (sub_ln703_765_reg_4852 + add_ln703_737_reg_4907);

assign add_ln703_739_fu_1966_p2 = (mult_704_V_reg_3765_pp0_iter6_reg + sub_ln703_703_fu_1519_p2);

assign add_ln703_740_fu_2532_p2 = (mult_770_V_reg_3814_pp0_iter7_reg + add_ln703_737_reg_4907);

assign add_ln703_741_fu_2536_p2 = (add_ln703_739_reg_4915 + add_ln703_740_fu_2532_p2);

assign add_ln703_742_fu_2569_p2 = (mult_896_V_reg_3909_pp0_iter7_reg + sub_ln703_792_fu_2351_p2);

assign add_ln703_743_fu_2583_p2 = (sub_ln703_768_fu_2141_p2 + add_ln703_737_reg_4907);

assign add_ln703_744_fu_2612_p2 = (mult_896_V_reg_3909_pp0_iter7_reg + sub_ln703_798_fu_2394_p2);

assign add_ln703_745_fu_2617_p2 = (mult_896_V_reg_3909_pp0_iter7_reg + sub_ln703_799_fu_2399_p2);

assign add_ln703_746_fu_2622_p2 = (mult_896_V_reg_3909_pp0_iter7_reg + sub_ln703_800_fu_2404_p2);

assign add_ln703_747_fu_2627_p2 = (mult_896_V_reg_3909_pp0_iter7_reg + sub_ln703_801_fu_2409_p2);

assign add_ln703_748_fu_2632_p2 = (mult_896_V_reg_3909_pp0_iter7_reg + sub_ln703_802_fu_2414_p2);

assign add_ln703_749_fu_2637_p2 = (sub_ln703_776_fu_2197_p2 + add_ln703_737_reg_4907);

assign add_ln703_750_fu_2669_p2 = (mult_832_V_reg_3861_pp0_iter7_reg + sub_ln703_753_reg_4834);

assign add_ln703_751_fu_1971_p2 = (mult_960_V_reg_3958_pp0_iter6_reg + mult_896_V_reg_3909_pp0_iter6_reg);

assign add_ln703_752_fu_2673_p2 = (add_ln703_750_fu_2669_p2 + add_ln703_751_reg_4920);

assign add_ln703_754_fu_2693_p2 = (mult_832_V_reg_3861_pp0_iter7_reg + sub_ln703_756_fu_2059_p2);

assign add_ln703_758_fu_2728_p2 = (mult_832_V_reg_3861_pp0_iter7_reg + sub_ln703_760_fu_2085_p2);

assign add_ln703_761_fu_2763_p2 = (mult_770_V_reg_3814_pp0_iter7_reg + sub_ln703_731_reg_4759);

assign add_ln703_762_fu_2767_p2 = (mult_832_V_reg_3861_pp0_iter7_reg + add_ln703_751_reg_4920);

assign add_ln703_765_fu_2792_p2 = (mult_832_V_reg_3861_pp0_iter7_reg + sub_ln703_764_fu_2113_p2);

assign add_ln703_770_fu_2867_p2 = (mult_832_V_reg_3861_pp0_iter7_reg + sub_ln703_767_fu_2127_p2);

assign add_ln703_776_fu_2937_p2 = (mult_832_V_reg_3861_pp0_iter7_reg + sub_ln703_772_fu_2166_p2);

assign add_ln703_778_fu_2947_p2 = (mult_832_V_reg_3861_pp0_iter7_reg + sub_ln703_773_fu_2171_p2);

assign add_ln703_780_fu_2957_p2 = (mult_832_V_reg_3861_pp0_iter7_reg + sub_ln703_774_fu_2176_p2);

assign add_ln703_782_fu_2992_p2 = (mult_832_V_reg_3861_pp0_iter7_reg + sub_ln703_777_fu_2202_p2);

assign add_ln703_786_fu_3027_p2 = (mult_770_V_reg_3814_pp0_iter7_reg + sub_ln703_752_reg_4824);

assign add_ln703_fu_242_p2 = (tmp_2_fu_92_p4 + trunc_ln203_fu_88_p1);

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_state1_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter4 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter5 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage0_iter6 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage0_iter7 = ~(1'b1 == 1'b1);

assign ap_block_state9_pp0_stage0_iter8 = ~(1'b1 == 1'b1);

assign sub_ln703_531_fu_252_p2 = (tmp_2_reg_3437 - trunc_ln203_reg_3431);

assign sub_ln703_532_fu_276_p2 = (sub_ln703_reg_4017_pp0_iter2_reg - tmp_3_reg_3443_pp0_iter2_reg);

assign sub_ln703_533_fu_264_p2 = (sub_ln703_531_reg_4023 - tmp_3_reg_3443_pp0_iter1_reg);

assign sub_ln703_534_fu_256_p2 = (add_ln703_reg_4010 - tmp_3_reg_3443);

assign sub_ln703_535_fu_284_p2 = (tmp_3_reg_3443_pp0_iter2_reg - add_ln703_reg_4010_pp0_iter2_reg);

assign sub_ln703_536_fu_340_p2 = (sub_ln703_532_reg_4061_pp0_iter4_reg - tmp_4_reg_3454_pp0_iter4_reg);

assign sub_ln703_537_fu_292_p2 = (sub_ln703_533_reg_4042 - tmp_4_reg_3454_pp0_iter2_reg);

assign sub_ln703_538_fu_268_p2 = (sub_ln703_534_reg_4029 - tmp_4_reg_3454_pp0_iter1_reg);

assign sub_ln703_539_fu_344_p2 = (add_ln703_538_reg_4067_pp0_iter4_reg - tmp_4_reg_3454_pp0_iter4_reg);

assign sub_ln703_540_fu_308_p2 = (tmp_4_reg_3454_pp0_iter3_reg - add_ln703_539_reg_4035_pp0_iter3_reg);

assign sub_ln703_541_fu_356_p2 = (add_ln703_540_reg_4079_pp0_iter4_reg - tmp_4_reg_3454_pp0_iter4_reg);

assign sub_ln703_542_fu_360_p2 = (sub_ln703_535_reg_4073_pp0_iter4_reg - tmp_4_reg_3454_pp0_iter4_reg);

assign sub_ln703_543_fu_296_p2 = (add_ln703_539_reg_4035_pp0_iter2_reg - tmp_4_reg_3454_pp0_iter2_reg);

assign sub_ln703_544_fu_316_p2 = (sub_ln703_537_reg_4085 - mult_307_V_reg_3472_pp0_iter3_reg);

assign sub_ln703_545_fu_300_p2 = (sub_ln703_538_reg_4048 - mult_307_V_reg_3472_pp0_iter2_reg);

assign sub_ln703_546_fu_442_p2 = (sub_ln703_539_reg_4165 - mult_307_V_reg_3472_pp0_iter5_reg);

assign sub_ln703_547_fu_446_p2 = (add_ln703_541_reg_4171 - mult_307_V_reg_3472_pp0_iter5_reg);

assign sub_ln703_548_fu_450_p2 = (add_ln703_542_reg_4177 - mult_307_V_reg_3472_pp0_iter5_reg);

assign sub_ln703_549_fu_372_p2 = (add_ln703_543_reg_4054_pp0_iter4_reg - mult_307_V_reg_3472_pp0_iter4_reg);

assign sub_ln703_550_fu_376_p2 = (mult_307_V_reg_3472_pp0_iter4_reg - add_ln703_543_reg_4054_pp0_iter4_reg);

assign sub_ln703_551_fu_380_p2 = (sub_ln703_540_reg_4110 - mult_307_V_reg_3472_pp0_iter4_reg);

assign sub_ln703_552_fu_388_p2 = (sub_ln703_541_fu_356_p2 - mult_307_V_reg_3472_pp0_iter4_reg);

assign sub_ln703_553_fu_462_p2 = (add_ln703_544_reg_4116_pp0_iter5_reg - mult_307_V_reg_3472_pp0_iter5_reg);

assign sub_ln703_554_fu_398_p2 = (sub_ln703_543_reg_4091_pp0_iter4_reg - mult_307_V_reg_3472_pp0_iter4_reg);

assign sub_ln703_555_fu_470_p2 = (sub_ln703_536_reg_4159 - mult_307_V_reg_3472_pp0_iter5_reg);

assign sub_ln703_556_fu_474_p2 = (add_ln703_545_reg_4183 - mult_307_V_reg_3472_pp0_iter5_reg);

assign sub_ln703_557_fu_402_p2 = (sub_ln703_544_reg_4122 - mult_320_V_reg_3500_pp0_iter4_reg);

assign sub_ln703_558_fu_328_p2 = (sub_ln703_545_reg_4097 - mult_320_V_reg_3500_pp0_iter3_reg);

assign sub_ln703_559_fu_483_p2 = (sub_ln703_546_fu_442_p2 - mult_320_V_reg_3500_pp0_iter5_reg);

assign sub_ln703_560_fu_493_p2 = (sub_ln703_548_fu_450_p2 - mult_320_V_reg_3500_pp0_iter5_reg);

assign sub_ln703_561_fu_502_p2 = (sub_ln703_549_reg_4194 - mult_320_V_reg_3500_pp0_iter5_reg);

assign sub_ln703_562_fu_506_p2 = (sub_ln703_550_reg_4200 - mult_320_V_reg_3500_pp0_iter5_reg);

assign sub_ln703_563_fu_514_p2 = (add_ln703_550_reg_4211 - mult_320_V_reg_3500_pp0_iter5_reg);

assign sub_ln703_564_fu_518_p2 = (mult_320_V_reg_3500_pp0_iter5_reg - add_ln703_549_reg_4103_pp0_iter5_reg);

assign sub_ln703_565_fu_530_p2 = (add_ln703_552_fu_454_p2 - mult_320_V_reg_3500_pp0_iter5_reg);

assign sub_ln703_566_fu_535_p2 = (add_ln703_553_fu_458_p2 - mult_320_V_reg_3500_pp0_iter5_reg);

assign sub_ln703_567_fu_540_p2 = (sub_ln703_553_fu_462_p2 - mult_320_V_reg_3500_pp0_iter5_reg);

assign sub_ln703_568_fu_545_p2 = (sub_ln703_551_reg_4205 - mult_320_V_reg_3500_pp0_iter5_reg);

assign sub_ln703_569_fu_549_p2 = (add_ln703_546_fu_438_p2 - mult_320_V_reg_3500_pp0_iter5_reg);

assign sub_ln703_570_fu_410_p2 = (add_ln703_554_reg_4134 - mult_320_V_reg_3500_pp0_iter4_reg);

assign sub_ln703_571_fu_558_p2 = (add_ln703_555_fu_466_p2 - mult_320_V_reg_3500_pp0_iter5_reg);

assign sub_ln703_572_fu_563_p2 = (sub_ln703_554_reg_4228 - mult_320_V_reg_3500_pp0_iter5_reg);

assign sub_ln703_573_fu_567_p2 = (sub_ln703_555_fu_470_p2 - mult_320_V_reg_3500_pp0_iter5_reg);

assign sub_ln703_574_fu_572_p2 = (sub_ln703_556_fu_474_p2 - mult_320_V_reg_3500_pp0_iter5_reg);

assign sub_ln703_575_fu_577_p2 = (add_ln703_548_reg_4188 - mult_320_V_reg_3500_pp0_iter5_reg);

assign sub_ln703_576_fu_414_p2 = (add_ln703_549_reg_4103_pp0_iter4_reg - mult_320_V_reg_3500_pp0_iter4_reg);

assign sub_ln703_577_fu_581_p2 = (add_ln703_551_reg_4222 - mult_320_V_reg_3500_pp0_iter5_reg);

assign sub_ln703_578_fu_585_p2 = (add_ln703_556_fu_478_p2 - mult_386_V_reg_3539_pp0_iter5_reg);

assign sub_ln703_579_fu_590_p2 = (sub_ln703_557_reg_4234 - mult_386_V_reg_3539_pp0_iter5_reg);

assign sub_ln703_580_fu_594_p2 = (sub_ln703_559_fu_483_p2 - mult_386_V_reg_3539_pp0_iter5_reg);

assign sub_ln703_581_fu_924_p2 = (add_ln703_557_reg_4293 - mult_386_V_reg_3539_pp0_iter6_reg);

assign sub_ln703_582_fu_599_p2 = (sub_ln703_560_fu_493_p2 - mult_386_V_reg_3539_pp0_iter5_reg);

assign sub_ln703_583_fu_604_p2 = (add_ln703_558_fu_498_p2 - mult_386_V_reg_3539_pp0_iter5_reg);

assign sub_ln703_584_fu_422_p2 = (add_ln703_559_reg_4146 - mult_386_V_reg_3539_pp0_iter4_reg);

assign sub_ln703_585_fu_609_p2 = (sub_ln703_561_fu_502_p2 - mult_386_V_reg_3539_pp0_iter5_reg);

assign sub_ln703_586_fu_614_p2 = (sub_ln703_562_fu_506_p2 - mult_386_V_reg_3539_pp0_iter5_reg);

assign sub_ln703_587_fu_619_p2 = (add_ln703_561_fu_510_p2 - mult_386_V_reg_3539_pp0_iter5_reg);

assign sub_ln703_588_fu_624_p2 = (add_ln703_562_fu_522_p2 - mult_386_V_reg_3539_pp0_iter5_reg);

assign sub_ln703_589_fu_638_p2 = (add_ln703_563_fu_526_p2 - mult_386_V_reg_3539_pp0_iter5_reg);

assign sub_ln703_590_fu_643_p2 = (sub_ln703_565_fu_530_p2 - mult_386_V_reg_3539_pp0_iter5_reg);

assign sub_ln703_591_fu_430_p2 = (mult_386_V_reg_3539_pp0_iter4_reg - add_ln703_559_reg_4146);

assign sub_ln703_592_fu_653_p2 = (sub_ln703_558_reg_4140_pp0_iter5_reg - mult_386_V_reg_3539_pp0_iter5_reg);

assign sub_ln703_593_fu_661_p2 = (sub_ln703_568_fu_545_p2 - mult_386_V_reg_3539_pp0_iter5_reg);

assign sub_ln703_594_fu_666_p2 = (add_ln703_564_reg_4240 - mult_386_V_reg_3539_pp0_iter5_reg);

assign sub_ln703_595_fu_928_p2 = (sub_ln703_567_reg_4303 - mult_386_V_reg_3539_pp0_iter6_reg);

assign sub_ln703_596_fu_683_p2 = (add_ln703_565_fu_554_p2 - mult_386_V_reg_3539_pp0_iter5_reg);

assign sub_ln703_597_fu_688_p2 = (sub_ln703_571_fu_558_p2 - mult_386_V_reg_3539_pp0_iter5_reg);

assign sub_ln703_598_fu_932_p2 = (sub_ln703_572_reg_4309 - mult_386_V_reg_3539_pp0_iter6_reg);

assign sub_ln703_599_fu_693_p2 = (sub_ln703_573_fu_567_p2 - mult_386_V_reg_3539_pp0_iter5_reg);

assign sub_ln703_600_fu_936_p2 = (sub_ln703_574_reg_4314 - mult_386_V_reg_3539_pp0_iter6_reg);

assign sub_ln703_601_fu_940_p2 = (sub_ln703_576_reg_4252_pp0_iter6_reg - mult_386_V_reg_3539_pp0_iter6_reg);

assign sub_ln703_602_fu_712_p2 = (sub_ln703_570_reg_4246 - mult_386_V_reg_3539_pp0_iter5_reg);

assign sub_ln703_603_fu_948_p2 = (sub_ln703_578_reg_4319 - mult_449_V_reg_3582_pp0_iter6_reg);

assign sub_ln703_604_fu_952_p2 = (add_ln703_566_reg_4258_pp0_iter6_reg - mult_449_V_reg_3582_pp0_iter6_reg);

assign sub_ln703_605_fu_720_p2 = (sub_ln703_580_fu_594_p2 - mult_449_V_reg_3582_pp0_iter5_reg);

assign sub_ln703_606_fu_956_p2 = (sub_ln703_581_fu_924_p2 - mult_449_V_reg_3582_pp0_iter6_reg);

assign sub_ln703_607_fu_961_p2 = (sub_ln703_582_reg_4329 - mult_449_V_reg_3582_pp0_iter6_reg);

assign sub_ln703_608_fu_725_p2 = (sub_ln703_583_fu_604_p2 - mult_449_V_reg_3582_pp0_iter5_reg);

assign sub_ln703_609_fu_965_p2 = (sub_ln703_585_reg_4334 - mult_449_V_reg_3582_pp0_iter6_reg);

assign sub_ln703_610_fu_734_p2 = (sub_ln703_586_fu_614_p2 - mult_449_V_reg_3582_pp0_iter5_reg);

assign sub_ln703_611_fu_739_p2 = (sub_ln703_587_fu_619_p2 - mult_449_V_reg_3582_pp0_iter5_reg);

assign sub_ln703_612_fu_969_p2 = (sub_ln703_588_reg_4350 - mult_449_V_reg_3582_pp0_iter6_reg);

assign sub_ln703_613_fu_758_p2 = (add_ln703_569_fu_633_p2 - mult_449_V_reg_3582_pp0_iter5_reg);

assign sub_ln703_614_fu_973_p2 = (sub_ln703_589_reg_4355 - mult_449_V_reg_3582_pp0_iter6_reg);

assign sub_ln703_615_fu_977_p2 = (sub_ln703_590_reg_4361 - mult_449_V_reg_3582_pp0_iter6_reg);

assign sub_ln703_616_fu_981_p2 = (sub_ln703_584_reg_4264_pp0_iter6_reg - mult_449_V_reg_3582_pp0_iter6_reg);

assign sub_ln703_617_fu_763_p2 = (add_ln703_570_fu_648_p2 - mult_449_V_reg_3582_pp0_iter5_reg);

assign sub_ln703_618_fu_768_p2 = (sub_ln703_591_reg_4277 - mult_449_V_reg_3582_pp0_iter5_reg);

assign sub_ln703_619_fu_989_p2 = (add_ln703_571_reg_4372 - mult_449_V_reg_3582_pp0_iter6_reg);

assign sub_ln703_620_fu_772_p2 = (sub_ln703_593_fu_661_p2 - mult_449_V_reg_3582_pp0_iter5_reg);

assign sub_ln703_621_fu_993_p2 = (sub_ln703_594_reg_4377 - mult_449_V_reg_3582_pp0_iter6_reg);

assign sub_ln703_622_fu_997_p2 = (sub_ln703_595_fu_928_p2 - mult_449_V_reg_3582_pp0_iter6_reg);

assign sub_ln703_623_fu_1002_p2 = (add_ln703_572_reg_4382 - mult_449_V_reg_3582_pp0_iter6_reg);

assign sub_ln703_624_fu_1006_p2 = (add_ln703_573_reg_4387 - mult_449_V_reg_3582_pp0_iter6_reg);

assign sub_ln703_625_fu_1010_p2 = (add_ln703_574_reg_4393 - mult_449_V_reg_3582_pp0_iter6_reg);

assign sub_ln703_626_fu_1014_p2 = (sub_ln703_599_reg_4403 - mult_449_V_reg_3582_pp0_iter6_reg);

assign sub_ln703_627_fu_807_p2 = (add_ln703_575_fu_698_p2 - mult_449_V_reg_3582_pp0_iter5_reg);

assign sub_ln703_628_fu_1018_p2 = (sub_ln703_592_reg_4366 - mult_449_V_reg_3582_pp0_iter6_reg);

assign sub_ln703_629_fu_1022_p2 = (sub_ln703_600_fu_936_p2 - mult_449_V_reg_3582_pp0_iter6_reg);

assign sub_ln703_630_fu_1035_p2 = (add_ln703_576_reg_4408 - mult_449_V_reg_3582_pp0_iter6_reg);

assign sub_ln703_631_fu_1039_p2 = (add_ln703_577_reg_4413 - mult_449_V_reg_3582_pp0_iter6_reg);

assign sub_ln703_632_fu_818_p2 = (sub_ln703_602_fu_712_p2 - mult_449_V_reg_3582_pp0_iter5_reg);

assign sub_ln703_633_fu_1043_p2 = (add_ln703_578_fu_944_p2 - mult_449_V_reg_3582_pp0_iter6_reg);

assign sub_ln703_634_fu_1048_p2 = (add_ln703_579_reg_4418 - mult_449_V_reg_3582_pp0_iter6_reg);

assign sub_ln703_635_fu_1056_p2 = (sub_ln703_605_reg_4423 - mult_512_V_reg_3629_pp0_iter6_reg);

assign sub_ln703_636_fu_1060_p2 = (sub_ln703_607_fu_961_p2 - mult_512_V_reg_3629_pp0_iter6_reg);

assign sub_ln703_637_fu_1065_p2 = (sub_ln703_608_reg_4428 - mult_512_V_reg_3629_pp0_iter6_reg);

assign sub_ln703_638_fu_1069_p2 = (add_ln703_580_reg_4433 - mult_512_V_reg_3629_pp0_iter6_reg);

assign sub_ln703_639_fu_1078_p2 = (sub_ln703_610_reg_4439 - mult_512_V_reg_3629_pp0_iter6_reg);

assign sub_ln703_640_fu_1082_p2 = (sub_ln703_611_reg_4444 - mult_512_V_reg_3629_pp0_iter6_reg);

assign sub_ln703_641_fu_838_p2 = (add_ln703_582_fu_748_p2 - mult_512_V_reg_3629_pp0_iter5_reg);

assign sub_ln703_642_fu_1086_p2 = (sub_ln703_612_fu_969_p2 - mult_512_V_reg_3629_pp0_iter6_reg);

assign sub_ln703_643_fu_1091_p2 = (add_ln703_583_reg_4450 - mult_512_V_reg_3629_pp0_iter6_reg);

assign sub_ln703_644_fu_1095_p2 = (sub_ln703_613_reg_4455 - mult_512_V_reg_3629_pp0_iter6_reg);

assign sub_ln703_645_fu_843_p2 = (sub_ln703_618_fu_768_p2 - mult_512_V_reg_3629_pp0_iter5_reg);

assign sub_ln703_646_fu_1099_p2 = (add_ln703_584_fu_985_p2 - mult_512_V_reg_3629_pp0_iter6_reg);

assign sub_ln703_647_fu_1104_p2 = (sub_ln703_620_reg_4466 - mult_512_V_reg_3629_pp0_iter6_reg);

assign sub_ln703_648_fu_1108_p2 = (sub_ln703_621_fu_993_p2 - mult_512_V_reg_3629_pp0_iter6_reg);

assign sub_ln703_649_fu_1113_p2 = (sub_ln703_623_fu_1002_p2 - mult_512_V_reg_3629_pp0_iter6_reg);

assign sub_ln703_650_fu_1118_p2 = (add_ln703_587_reg_4471 - mult_512_V_reg_3629_pp0_iter6_reg);

assign sub_ln703_651_fu_1122_p2 = (sub_ln703_624_fu_1006_p2 - mult_512_V_reg_3629_pp0_iter6_reg);

assign sub_ln703_652_fu_1127_p2 = (sub_ln703_625_fu_1010_p2 - mult_512_V_reg_3629_pp0_iter6_reg);

assign sub_ln703_653_fu_1136_p2 = (add_ln703_588_reg_4476 - mult_512_V_reg_3629_pp0_iter6_reg);

assign sub_ln703_654_fu_1145_p2 = (add_ln703_590_reg_4481 - mult_512_V_reg_3629_pp0_iter6_reg);

assign sub_ln703_655_fu_1149_p2 = (sub_ln703_627_reg_4486 - mult_512_V_reg_3629_pp0_iter6_reg);

assign sub_ln703_656_fu_1153_p2 = (add_ln703_591_fu_1027_p2 - mult_512_V_reg_3629_pp0_iter6_reg);

assign sub_ln703_657_fu_1158_p2 = (add_ln703_592_fu_1031_p2 - mult_512_V_reg_3629_pp0_iter6_reg);

assign sub_ln703_658_fu_1167_p2 = (sub_ln703_617_reg_4460 - mult_512_V_reg_3629_pp0_iter6_reg);

assign sub_ln703_659_fu_1171_p2 = (sub_ln703_630_fu_1035_p2 - mult_512_V_reg_3629_pp0_iter6_reg);

assign sub_ln703_660_fu_872_p2 = (add_ln703_593_fu_812_p2 - mult_512_V_reg_3629_pp0_iter5_reg);

assign sub_ln703_661_fu_877_p2 = (add_ln703_594_fu_823_p2 - mult_512_V_reg_3629_pp0_iter5_reg);

assign sub_ln703_662_fu_882_p2 = (add_ln703_596_fu_832_p2 - mult_512_V_reg_3629_pp0_iter5_reg);

assign sub_ln703_663_fu_1189_p2 = (add_ln703_598_fu_1052_p2 - mult_576_V_reg_3674_pp0_iter6_reg);

assign sub_ln703_664_fu_1199_p2 = (sub_ln703_635_fu_1056_p2 - mult_576_V_reg_3674_pp0_iter6_reg);

assign sub_ln703_665_fu_1204_p2 = (sub_ln703_637_fu_1065_p2 - mult_576_V_reg_3674_pp0_iter6_reg);

assign sub_ln703_666_fu_1214_p2 = (add_ln703_599_fu_1073_p2 - mult_576_V_reg_3674_pp0_iter6_reg);

assign sub_ln703_667_fu_1224_p2 = (sub_ln703_641_reg_4496 - mult_576_V_reg_3674_pp0_iter6_reg);

assign sub_ln703_668_fu_1233_p2 = (sub_ln703_644_fu_1095_p2 - mult_576_V_reg_3674_pp0_iter6_reg);

assign sub_ln703_669_fu_1261_p2 = (sub_ln703_636_fu_1060_p2 - mult_576_V_reg_3674_pp0_iter6_reg);

assign sub_ln703_670_fu_1266_p2 = (sub_ln703_647_fu_1104_p2 - mult_576_V_reg_3674_pp0_iter6_reg);

assign sub_ln703_671_fu_896_p2 = (add_ln703_602_fu_856_p2 - mult_576_V_reg_3674_pp0_iter5_reg);

assign sub_ln703_672_fu_1281_p2 = (sub_ln703_651_fu_1122_p2 - mult_576_V_reg_3674_pp0_iter6_reg);

assign sub_ln703_673_fu_1291_p2 = (add_ln703_603_fu_1132_p2 - mult_576_V_reg_3674_pp0_iter6_reg);

assign sub_ln703_674_fu_1296_p2 = (sub_ln703_653_fu_1136_p2 - mult_576_V_reg_3674_pp0_iter6_reg);

assign sub_ln703_675_fu_1301_p2 = (add_ln703_604_fu_1140_p2 - mult_576_V_reg_3674_pp0_iter6_reg);

assign sub_ln703_676_fu_901_p2 = (add_ln703_606_fu_866_p2 - mult_576_V_reg_3674_pp0_iter5_reg);

assign sub_ln703_677_fu_1306_p2 = (sub_ln703_655_fu_1149_p2 - mult_576_V_reg_3674_pp0_iter6_reg);

assign sub_ln703_678_fu_1316_p2 = (sub_ln703_656_fu_1153_p2 - mult_576_V_reg_3674_pp0_iter6_reg);

assign sub_ln703_679_fu_1330_p2 = (sub_ln703_657_fu_1158_p2 - mult_576_V_reg_3674_pp0_iter6_reg);

assign sub_ln703_680_fu_1335_p2 = (add_ln703_607_fu_1163_p2 - mult_576_V_reg_3674_pp0_iter6_reg);

assign sub_ln703_681_fu_1340_p2 = (sub_ln703_658_fu_1167_p2 - mult_576_V_reg_3674_pp0_iter6_reg);

assign sub_ln703_682_fu_1345_p2 = (sub_ln703_659_fu_1171_p2 - mult_576_V_reg_3674_pp0_iter6_reg);

assign sub_ln703_683_fu_1360_p2 = (add_ln703_608_fu_1176_p2 - mult_576_V_reg_3674_pp0_iter6_reg);

assign sub_ln703_684_fu_1365_p2 = (add_ln703_609_fu_1181_p2 - mult_576_V_reg_3674_pp0_iter6_reg);

assign sub_ln703_685_fu_1370_p2 = (sub_ln703_661_reg_4511 - mult_576_V_reg_3674_pp0_iter6_reg);

assign sub_ln703_686_fu_1374_p2 = (sub_ln703_662_reg_4516 - mult_576_V_reg_3674_pp0_iter6_reg);

assign sub_ln703_687_fu_1378_p2 = (sub_ln703_645_reg_4501 - mult_576_V_reg_3674_pp0_iter6_reg);

assign sub_ln703_688_fu_1382_p2 = (add_ln703_610_fu_1185_p2 - mult_576_V_reg_3674_pp0_iter6_reg);

assign sub_ln703_689_fu_1392_p2 = (sub_ln703_663_fu_1189_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_690_fu_1402_p2 = (sub_ln703_664_fu_1199_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_691_fu_1428_p2 = (sub_ln703_665_fu_1204_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_692_fu_1433_p2 = (add_ln703_613_fu_1209_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_693_fu_1438_p2 = (sub_ln703_666_fu_1214_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_694_fu_1443_p2 = (add_ln703_614_fu_1219_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_695_fu_1464_p2 = (sub_ln703_667_fu_1224_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_696_fu_1475_p2 = (add_ln703_615_fu_1228_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_697_fu_1485_p2 = (add_ln703_616_fu_1238_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_698_fu_1490_p2 = (add_ln703_617_fu_1243_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_699_fu_1495_p2 = (add_ln703_618_fu_1248_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_700_fu_1500_p2 = (add_ln703_619_fu_1252_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_701_fu_1509_p2 = (add_ln703_621_fu_1256_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_702_fu_1514_p2 = (sub_ln703_669_fu_1261_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_703_fu_1519_p2 = (sub_ln703_670_fu_1266_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_704_fu_1524_p2 = (add_ln703_622_fu_1271_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_705_fu_1544_p2 = (add_ln703_620_reg_4537 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_706_fu_1548_p2 = (add_ln703_623_fu_1276_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_707_fu_1559_p2 = (sub_ln703_672_fu_1281_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_708_fu_1564_p2 = (add_ln703_624_fu_1286_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_709_fu_1569_p2 = (add_ln703_612_fu_1194_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_710_fu_1606_p2 = (add_ln703_625_fu_1311_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_711_fu_1611_p2 = (sub_ln703_678_fu_1316_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_712_fu_1616_p2 = (add_ln703_627_fu_1325_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_713_fu_1621_p2 = (sub_ln703_681_fu_1340_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_714_fu_1626_p2 = (sub_ln703_682_fu_1345_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_715_fu_1631_p2 = (add_ln703_629_fu_1355_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_716_fu_1636_p2 = (sub_ln703_683_fu_1360_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_717_fu_1641_p2 = (sub_ln703_684_fu_1365_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_718_fu_1646_p2 = (sub_ln703_686_fu_1374_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_719_fu_1656_p2 = (add_ln703_630_fu_1387_p2 - mult_640_V_reg_3716_pp0_iter6_reg);

assign sub_ln703_720_fu_1676_p2 = (sub_ln703_689_fu_1392_p2 - mult_704_V_reg_3765_pp0_iter6_reg);

assign sub_ln703_721_fu_1975_p2 = (add_ln703_631_reg_4588 - mult_704_V_reg_3765_pp0_iter7_reg);

assign sub_ln703_722_fu_1681_p2 = (sub_ln703_690_fu_1402_p2 - mult_704_V_reg_3765_pp0_iter6_reg);

assign sub_ln703_723_fu_1979_p2 = (add_ln703_634_reg_4593 - mult_704_V_reg_3765_pp0_iter7_reg);

assign sub_ln703_724_fu_1686_p2 = (add_ln703_635_fu_1422_p2 - mult_704_V_reg_3765_pp0_iter6_reg);

assign sub_ln703_725_fu_1691_p2 = (sub_ln703_691_fu_1428_p2 - mult_704_V_reg_3765_pp0_iter6_reg);

assign sub_ln703_726_fu_1983_p2 = (sub_ln703_693_reg_4603 - mult_704_V_reg_3765_pp0_iter7_reg);

assign sub_ln703_727_fu_1701_p2 = (add_ln703_636_fu_1448_p2 - mult_704_V_reg_3765_pp0_iter6_reg);

assign sub_ln703_728_fu_1987_p2 = (add_ln703_639_reg_4608 - mult_704_V_reg_3765_pp0_iter7_reg);

assign sub_ln703_729_fu_1715_p2 = (add_ln703_640_fu_1469_p2 - mult_704_V_reg_3765_pp0_iter6_reg);

assign sub_ln703_730_fu_1720_p2 = (sub_ln703_696_fu_1475_p2 - mult_704_V_reg_3765_pp0_iter6_reg);

assign sub_ln703_731_fu_1725_p2 = (add_ln703_641_fu_1480_p2 - mult_704_V_reg_3765_pp0_iter6_reg);

assign sub_ln703_732_fu_1741_p2 = (sub_ln703_697_fu_1485_p2 - mult_704_V_reg_3765_pp0_iter6_reg);

assign sub_ln703_733_fu_1995_p2 = (sub_ln703_700_reg_4623 - mult_704_V_reg_3765_pp0_iter7_reg);

assign sub_ln703_734_fu_1999_p2 = (add_ln703_642_reg_4628 - mult_704_V_reg_3765_pp0_iter7_reg);

assign sub_ln703_735_fu_2003_p2 = (sub_ln703_701_reg_4633 - mult_704_V_reg_3765_pp0_iter7_reg);

assign sub_ln703_736_fu_2007_p2 = (sub_ln703_702_reg_4638 - mult_704_V_reg_3765_pp0_iter7_reg);

assign sub_ln703_737_fu_2011_p2 = (add_ln703_645_reg_4648 - mult_704_V_reg_3765_pp0_iter7_reg);

assign sub_ln703_738_fu_1757_p2 = (sub_ln703_705_fu_1544_p2 - mult_704_V_reg_3765_pp0_iter6_reg);

assign sub_ln703_739_fu_2015_p2 = (add_ln703_646_reg_4658 - mult_704_V_reg_3765_pp0_iter7_reg);

assign sub_ln703_740_fu_2019_p2 = (sub_ln703_707_reg_4663 - mult_704_V_reg_3765_pp0_iter7_reg);

assign sub_ln703_741_fu_2023_p2 = (sub_ln703_709_reg_4673 - mult_704_V_reg_3765_pp0_iter7_reg);

assign sub_ln703_742_fu_1762_p2 = (add_ln703_647_fu_1574_p2 - mult_704_V_reg_3765_pp0_iter6_reg);

assign sub_ln703_743_fu_1772_p2 = (add_ln703_649_fu_1584_p2 - mult_704_V_reg_3765_pp0_iter6_reg);

assign sub_ln703_744_fu_1777_p2 = (add_ln703_650_fu_1590_p2 - mult_704_V_reg_3765_pp0_iter6_reg);

assign sub_ln703_745_fu_1782_p2 = (add_ln703_652_fu_1600_p2 - mult_704_V_reg_3765_pp0_iter6_reg);

assign sub_ln703_746_fu_2027_p2 = (sub_ln703_710_reg_4678 - mult_704_V_reg_3765_pp0_iter7_reg);

assign sub_ln703_747_fu_2031_p2 = (sub_ln703_711_reg_4683 - mult_704_V_reg_3765_pp0_iter7_reg);

assign sub_ln703_748_fu_1792_p2 = (sub_ln703_713_fu_1621_p2 - mult_704_V_reg_3765_pp0_iter6_reg);

assign sub_ln703_749_fu_2039_p2 = (sub_ln703_715_reg_4698 - mult_704_V_reg_3765_pp0_iter7_reg);

assign sub_ln703_750_fu_2043_p2 = (sub_ln703_716_reg_4703 - mult_704_V_reg_3765_pp0_iter7_reg);

assign sub_ln703_751_fu_1797_p2 = (sub_ln703_717_fu_1641_p2 - mult_704_V_reg_3765_pp0_iter6_reg);

assign sub_ln703_752_fu_1807_p2 = (add_ln703_653_fu_1651_p2 - mult_704_V_reg_3765_pp0_iter6_reg);

assign sub_ln703_753_fu_1817_p2 = (add_ln703_657_fu_1670_p2 - mult_770_V_reg_3814_pp0_iter6_reg);

assign sub_ln703_754_fu_2051_p2 = (sub_ln703_720_reg_4713 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_755_fu_2055_p2 = (sub_ln703_722_reg_4718 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_756_fu_2059_p2 = (sub_ln703_723_fu_1979_p2 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_757_fu_2064_p2 = (sub_ln703_724_reg_4723 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_758_fu_2076_p2 = (sub_ln703_726_fu_1983_p2 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_759_fu_2081_p2 = (add_ln703_658_reg_4733 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_760_fu_2085_p2 = (sub_ln703_727_reg_4738 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_761_fu_2089_p2 = (add_ln703_661_reg_4744 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_762_fu_2097_p2 = (sub_ln703_729_reg_4749 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_763_fu_2105_p2 = (add_ln703_663_reg_4764 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_764_fu_2113_p2 = (add_ln703_664_fu_1991_p2 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_765_fu_1832_p2 = (add_ln703_666_fu_1751_p2 - mult_770_V_reg_3814_pp0_iter6_reg);

assign sub_ln703_766_fu_2123_p2 = (sub_ln703_738_reg_4774 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_767_fu_2127_p2 = (sub_ln703_739_fu_2015_p2 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_768_fu_2141_p2 = (sub_ln703_741_fu_2023_p2 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_769_fu_2150_p2 = (add_ln703_667_reg_4784 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_770_fu_2158_p2 = (sub_ln703_744_reg_4794 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_771_fu_2162_p2 = (sub_ln703_745_reg_4799 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_772_fu_2166_p2 = (sub_ln703_746_fu_2027_p2 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_773_fu_2171_p2 = (sub_ln703_747_fu_2031_p2 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_774_fu_2176_p2 = (add_ln703_668_fu_2035_p2 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_775_fu_2185_p2 = (add_ln703_669_reg_4804 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_776_fu_2197_p2 = (sub_ln703_749_fu_2039_p2 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_777_fu_2202_p2 = (sub_ln703_750_fu_2043_p2 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_778_fu_2207_p2 = (sub_ln703_751_reg_4814 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_779_fu_2211_p2 = (add_ln703_670_reg_4819 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_780_fu_2215_p2 = (add_ln703_671_fu_2047_p2 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_781_fu_2220_p2 = (add_ln703_672_reg_4829 - mult_770_V_reg_3814_pp0_iter7_reg);

assign sub_ln703_782_fu_2224_p2 = (sub_ln703_754_fu_2051_p2 - mult_832_V_reg_3861_pp0_iter7_reg);

assign sub_ln703_783_fu_2244_p2 = (add_ln703_673_fu_2068_p2 - mult_832_V_reg_3861_pp0_iter7_reg);

assign sub_ln703_784_fu_2249_p2 = (add_ln703_675_fu_2072_p2 - mult_832_V_reg_3861_pp0_iter7_reg);

assign sub_ln703_785_fu_2254_p2 = (sub_ln703_758_fu_2076_p2 - mult_832_V_reg_3861_pp0_iter7_reg);

assign sub_ln703_786_fu_2259_p2 = (sub_ln703_759_fu_2081_p2 - mult_832_V_reg_3861_pp0_iter7_reg);

assign sub_ln703_787_fu_2274_p2 = (add_ln703_676_fu_2093_p2 - mult_832_V_reg_3861_pp0_iter7_reg);

assign sub_ln703_788_fu_2284_p2 = (add_ln703_677_fu_2101_p2 - mult_832_V_reg_3861_pp0_iter7_reg);

assign sub_ln703_789_fu_2294_p2 = (add_ln703_678_fu_2109_p2 - mult_832_V_reg_3861_pp0_iter7_reg);

assign sub_ln703_790_fu_2299_p2 = (add_ln703_679_reg_4847 - mult_832_V_reg_3861_pp0_iter7_reg);

assign sub_ln703_791_fu_2318_p2 = (add_ln703_680_fu_2118_p2 - mult_832_V_reg_3861_pp0_iter7_reg);

assign sub_ln703_792_fu_2351_p2 = (add_ln703_681_fu_2132_p2 - mult_832_V_reg_3861_pp0_iter7_reg);

assign sub_ln703_793_fu_2356_p2 = (add_ln703_682_fu_2136_p2 - mult_832_V_reg_3861_pp0_iter7_reg);

assign sub_ln703_794_fu_2370_p2 = (add_ln703_683_fu_2146_p2 - mult_832_V_reg_3861_pp0_iter7_reg);

assign sub_ln703_795_fu_2375_p2 = (sub_ln703_769_fu_2150_p2 - mult_832_V_reg_3861_pp0_iter7_reg);

assign sub_ln703_796_fu_2380_p2 = (add_ln703_684_fu_2154_p2 - mult_832_V_reg_3861_pp0_iter7_reg);

assign sub_ln703_797_fu_2385_p2 = (add_ln703_687_reg_4857 - mult_832_V_reg_3861_pp0_iter7_reg);

assign sub_ln703_798_fu_2394_p2 = (sub_ln703_771_fu_2162_p2 - mult_832_V_reg_3861_pp0_iter7_reg);

assign sub_ln703_799_fu_2399_p2 = (add_ln703_689_fu_2181_p2 - mult_832_V_reg_3861_pp0_iter7_reg);

assign sub_ln703_800_fu_2404_p2 = (sub_ln703_775_fu_2185_p2 - mult_832_V_reg_3861_pp0_iter7_reg);

assign sub_ln703_801_fu_2409_p2 = (add_ln703_690_fu_2189_p2 - mult_832_V_reg_3861_pp0_iter7_reg);

assign sub_ln703_802_fu_2414_p2 = (add_ln703_691_fu_2193_p2 - mult_832_V_reg_3861_pp0_iter7_reg);

assign sub_ln703_803_fu_2419_p2 = (sub_ln703_778_fu_2207_p2 - mult_832_V_reg_3861_pp0_iter7_reg);

assign sub_ln703_804_fu_2429_p2 = (sub_ln703_780_fu_2215_p2 - mult_832_V_reg_3861_pp0_iter7_reg);

assign sub_ln703_805_fu_2439_p2 = (sub_ln703_782_fu_2224_p2 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_806_fu_2444_p2 = (add_ln703_693_fu_2229_p2 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_807_fu_2449_p2 = (add_ln703_694_fu_2234_p2 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_808_fu_2454_p2 = (add_ln703_695_fu_2239_p2 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_809_fu_2459_p2 = (sub_ln703_783_fu_2244_p2 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_810_fu_2464_p2 = (sub_ln703_784_fu_2249_p2 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_811_fu_2474_p2 = (add_ln703_696_fu_2264_p2 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_812_fu_2479_p2 = (add_ln703_697_fu_2269_p2 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_813_fu_2489_p2 = (add_ln703_698_fu_2279_p2 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_814_fu_2494_p2 = (sub_ln703_788_fu_2284_p2 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_815_fu_2499_p2 = (add_ln703_699_fu_2289_p2 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_816_fu_2509_p2 = (add_ln703_700_fu_2303_p2 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_817_fu_2514_p2 = (add_ln703_701_fu_2308_p2 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_818_fu_2519_p2 = (add_ln703_702_fu_2313_p2 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_819_fu_2524_p2 = (add_ln703_707_reg_4867 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_820_fu_2541_p2 = (add_ln703_709_fu_2327_p2 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_821_fu_2546_p2 = (add_ln703_711_reg_4872 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_822_fu_2550_p2 = (add_ln703_712_fu_2332_p2 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_823_fu_2555_p2 = (add_ln703_713_fu_2337_p2 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_824_fu_2560_p2 = (add_ln703_716_reg_4877 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_825_fu_2564_p2 = (add_ln703_718_fu_2346_p2 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_826_fu_2574_p2 = (add_ln703_720_fu_2365_p2 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_827_fu_2579_p2 = (add_ln703_722_reg_4882 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_828_fu_2588_p2 = (sub_ln703_794_fu_2370_p2 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_829_fu_2593_p2 = (sub_ln703_795_fu_2375_p2 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_830_fu_2598_p2 = (add_ln703_724_reg_4887 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_831_fu_2602_p2 = (sub_ln703_796_fu_2380_p2 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_832_fu_2607_p2 = (add_ln703_725_fu_2389_p2 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_833_fu_2642_p2 = (add_ln703_727_reg_4892 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_834_fu_2646_p2 = (sub_ln703_803_fu_2419_p2 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_835_fu_2651_p2 = (add_ln703_729_reg_4897 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_836_fu_2655_p2 = (add_ln703_730_fu_2424_p2 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_837_fu_2660_p2 = (add_ln703_732_reg_4902 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_838_fu_2664_p2 = (add_ln703_733_fu_2434_p2 - mult_896_V_reg_3909_pp0_iter7_reg);

assign sub_ln703_fu_248_p2 = (trunc_ln203_reg_3431 - tmp_2_reg_3437);

assign tmp_2_fu_92_p4 = {{data_V_read_int_reg[31:16]}};

assign trunc_ln203_fu_88_p1 = data_V_read_int_reg[15:0];

endmodule //dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_1
