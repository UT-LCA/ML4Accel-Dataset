`define M     593         // M is the degree of the irreducible polynomial
`define WIDTH (2*`M-1)    // width for a GF(3^M) element
`define WIDTH_D0 1187
`define M     593         // M is the degree of the irreducible polynomial
`define WIDTH (2*`M-1)    // width for a GF(3^M) element
`define WIDTH_D0 1187
`define M     593         // M is the degree of the irreducible polynomial
`define WIDTH (2*`M-1)    // width for a GF(3^M) element
`define WIDTH_D0 1187
`define M     593         // M is the degree of the irreducible polynomial
`define WIDTH (2*`M-1)    // width for a GF(3^M) element
`define WIDTH_D0 1187
`define M     593         // M is the degree of the irreducible polynomial
`define WIDTH (2*`M-1)    // width for a GF(3^M) element
`define WIDTH_D0 1187

module v0(a, c);
    input [1185:0] a;
    output [1185:0] c;
    assign c[1:0] = a[1:0];
    assign c[3:2] = a[1113:1112];
    assign c[5:4] = a[793:792];
    assign c[7:6] = a[3:2];
    assign c[9:8] = a[1115:1114];
    assign c[11:10] = a[1041:1040];
    assign c[13:12] = {a[720], a[721]};
    assign c[15:14] = a[401:400];
    assign c[17:16] = a[1043:1042];
    assign c[19:18] = {a[722], a[723]};
    assign c[21:20] = a[403:402];
    assign c[23:22] = a[1045:1044];
    assign c[25:24] = {a[724], a[725]};
    assign c[27:26] = a[1121:1120];
    assign c[29:28] = a[801:800];
    assign c[31:30] = {a[726], a[727]};
    assign c[33:32] = a[1123:1122];
    assign c[35:34] = a[803:802];
    assign c[37:36] = {a[728], a[729]};
    assign c[39:38] = a[1125:1124];
    assign c[41:40] = a[805:804];
    assign c[43:42] = {a[730], a[731]};
    assign c[45:44] = a[1127:1126];
    assign c[47:46] = a[807:806];
    assign c[49:48] = a[17:16];
    assign c[51:50] = a[1129:1128];
    assign c[53:52] = a[809:808];
    assign c[55:54] = a[19:18];
    assign c[57:56] = a[1131:1130];
    assign c[59:58] = a[1057:1056];
    assign c[61:60] = {a[736], a[737]};
    assign c[63:62] = a[417:416];
    assign c[65:64] = a[1059:1058];
    assign c[67:66] = {a[738], a[739]};
    assign c[69:68] = a[419:418];
    assign c[71:70] = a[1061:1060];
    assign c[73:72] = {a[740], a[741]};
    assign c[75:74] = a[1137:1136];
    assign c[77:76] = a[817:816];
    assign c[79:78] = {a[742], a[743]};
    assign c[81:80] = a[1139:1138];
    assign c[83:82] = a[819:818];
    assign c[85:84] = {a[744], a[745]};
    assign c[87:86] = a[1141:1140];
    assign c[89:88] = a[821:820];
    assign c[91:90] = {a[746], a[747]};
    assign c[93:92] = a[1143:1142];
    assign c[95:94] = a[823:822];
    assign c[97:96] = a[33:32];
    assign c[99:98] = a[1145:1144];
    assign c[101:100] = a[825:824];
    assign c[103:102] = a[35:34];
    assign c[105:104] = a[1147:1146];
    assign c[107:106] = a[1073:1072];
    assign c[109:108] = {a[752], a[753]};
    assign c[111:110] = a[433:432];
    assign c[113:112] = a[1075:1074];
    assign c[115:114] = {a[754], a[755]};
    assign c[117:116] = a[435:434];
    assign c[119:118] = a[1077:1076];
    assign c[121:120] = {a[756], a[757]};
    assign c[123:122] = a[1153:1152];
    assign c[125:124] = a[833:832];
    assign c[127:126] = {a[758], a[759]};
    assign c[129:128] = a[1155:1154];
    assign c[131:130] = a[835:834];
    assign c[133:132] = {a[760], a[761]};
    assign c[135:134] = a[1157:1156];
    assign c[137:136] = a[837:836];
    assign c[139:138] = {a[762], a[763]};
    assign c[141:140] = a[1159:1158];
    assign c[143:142] = a[839:838];
    assign c[145:144] = a[49:48];
    assign c[147:146] = a[1161:1160];
    assign c[149:148] = a[841:840];
    assign c[151:150] = a[51:50];
    assign c[153:152] = a[1163:1162];
    assign c[155:154] = a[1089:1088];
    assign c[157:156] = {a[768], a[769]};
    assign c[159:158] = a[449:448];
    assign c[161:160] = a[1091:1090];
    assign c[163:162] = {a[770], a[771]};
    assign c[165:164] = a[451:450];
    assign c[167:166] = a[1093:1092];
    assign c[169:168] = {a[772], a[773]};
    assign c[171:170] = a[1169:1168];
    assign c[173:172] = a[849:848];
    assign c[175:174] = {a[774], a[775]};
    assign c[177:176] = a[1171:1170];
    assign c[179:178] = a[851:850];
    assign c[181:180] = {a[776], a[777]};
    assign c[183:182] = a[1173:1172];
    assign c[185:184] = a[853:852];
    assign c[187:186] = {a[778], a[779]};
    assign c[189:188] = a[1175:1174];
    assign c[191:190] = a[855:854];
    assign c[193:192] = a[65:64];
    assign c[195:194] = a[1177:1176];
    assign c[197:196] = a[857:856];
    assign c[199:198] = a[67:66];
    assign c[201:200] = a[1179:1178];
    assign c[203:202] = a[1105:1104];
    assign c[205:204] = {a[784], a[785]};
    assign c[207:206] = a[465:464];
    assign c[209:208] = a[1107:1106];
    assign c[211:210] = {a[786], a[787]};
    assign c[213:212] = a[467:466];
    assign c[215:214] = a[1109:1108];
    assign c[217:216] = {a[788], a[789]};
    assign c[219:218] = a[1185:1184];
    assign c[221:220] = a[865:864];
    assign c[223:222] = {a[790], a[791]};
    assign c[225:224] = a[471:470];
    assign c[227:226] = a[867:866];
    assign c[229:228] = a[793:792];
    assign c[231:230] = a[473:472];
    assign c[233:232] = a[869:868];
    assign c[235:234] = {a[1040], a[1041]};
    assign c[237:236] = a[721:720];
    assign c[239:238] = {a[400], a[401]};
    assign c[241:240] = a[81:80];
    assign c[243:242] = a[723:722];
    assign c[245:244] = {a[402], a[403]};
    assign c[247:246] = a[83:82];
    assign c[249:248] = a[725:724];
    assign c[251:250] = {a[404], a[405]};
    assign c[253:252] = a[801:800];
    assign c[255:254] = a[481:480];
    assign c[257:256] = {a[406], a[407]};
    assign c[259:258] = a[803:802];
    assign c[261:260] = a[483:482];
    assign c[263:262] = {a[408], a[409]};
    assign c[265:264] = a[805:804];
    assign c[267:266] = a[485:484];
    assign c[269:268] = a[881:880];
    assign c[271:270] = a[807:806];
    assign c[273:272] = a[487:486];
    assign c[275:274] = a[883:882];
    assign c[277:276] = a[809:808];
    assign c[279:278] = a[489:488];
    assign c[281:280] = a[885:884];
    assign c[283:282] = {a[1056], a[1057]};
    assign c[285:284] = a[737:736];
    assign c[287:286] = {a[416], a[417]};
    assign c[289:288] = a[97:96];
    assign c[291:290] = a[739:738];
    assign c[293:292] = {a[418], a[419]};
    assign c[295:294] = a[99:98];
    assign c[297:296] = a[741:740];
    assign c[299:298] = {a[420], a[421]};
    assign c[301:300] = a[817:816];
    assign c[303:302] = a[497:496];
    assign c[305:304] = {a[422], a[423]};
    assign c[307:306] = a[819:818];
    assign c[309:308] = a[499:498];
    assign c[311:310] = {a[424], a[425]};
    assign c[313:312] = a[821:820];
    assign c[315:314] = a[501:500];
    assign c[317:316] = a[897:896];
    assign c[319:318] = a[823:822];
    assign c[321:320] = a[503:502];
    assign c[323:322] = a[899:898];
    assign c[325:324] = a[825:824];
    assign c[327:326] = a[505:504];
    assign c[329:328] = a[901:900];
    assign c[331:330] = {a[1072], a[1073]};
    assign c[333:332] = a[753:752];
    assign c[335:334] = {a[432], a[433]};
    assign c[337:336] = a[113:112];
    assign c[339:338] = a[755:754];
    assign c[341:340] = {a[434], a[435]};
    assign c[343:342] = a[115:114];
    assign c[345:344] = a[757:756];
    assign c[347:346] = {a[436], a[437]};
    assign c[349:348] = a[833:832];
    assign c[351:350] = a[513:512];
    assign c[353:352] = {a[438], a[439]};
    assign c[355:354] = a[835:834];
    assign c[357:356] = a[515:514];
    assign c[359:358] = {a[440], a[441]};
    assign c[361:360] = a[837:836];
    assign c[363:362] = a[517:516];
    assign c[365:364] = a[913:912];
    assign c[367:366] = a[839:838];
    assign c[369:368] = a[519:518];
    assign c[371:370] = a[915:914];
    assign c[373:372] = a[841:840];
    assign c[375:374] = a[521:520];
    assign c[377:376] = a[917:916];
    assign c[379:378] = {a[1088], a[1089]};
    assign c[381:380] = a[769:768];
    assign c[383:382] = {a[448], a[449]};
    assign c[385:384] = a[129:128];
    assign c[387:386] = a[771:770];
    assign c[389:388] = {a[450], a[451]};
    assign c[391:390] = a[131:130];
    assign c[393:392] = a[773:772];
    assign c[395:394] = {a[452], a[453]};
    assign c[397:396] = a[849:848];
    assign c[399:398] = a[529:528];
    assign c[401:400] = {a[454], a[455]};
    assign c[403:402] = a[851:850];
    assign c[405:404] = a[531:530];
    assign c[407:406] = {a[456], a[457]};
    assign c[409:408] = a[853:852];
    assign c[411:410] = a[533:532];
    assign c[413:412] = a[929:928];
    assign c[415:414] = a[855:854];
    assign c[417:416] = a[535:534];
    assign c[419:418] = a[931:930];
    assign c[421:420] = a[857:856];
    assign c[423:422] = a[537:536];
    assign c[425:424] = a[933:932];
    assign c[427:426] = {a[1104], a[1105]};
    assign c[429:428] = a[785:784];
    assign c[431:430] = {a[464], a[465]};
    assign c[433:432] = a[145:144];
    assign c[435:434] = a[787:786];
    assign c[437:436] = {a[466], a[467]};
    assign c[439:438] = a[147:146];
    assign c[441:440] = a[789:788];
    assign c[443:442] = {a[468], a[469]};
    assign c[445:444] = a[865:864];
    assign c[447:446] = a[545:544];
    assign c[449:448] = {a[470], a[471]};
    assign c[451:450] = a[867:866];
    assign c[453:452] = a[547:546];
    assign c[455:454] = {a[472], a[473]};
    assign c[457:456] = a[869:868];
    assign c[459:458] = a[549:548];
    assign c[461:460] = a[945:944];
    assign c[463:462] = a[871:870];
    assign c[465:464] = a[551:550];
    assign c[467:466] = a[947:946];
    assign c[469:468] = a[873:872];
    assign c[471:470] = a[553:552];
    assign c[473:472] = a[949:948];
    assign c[475:474] = {a[1120], a[1121]};
    assign c[477:476] = a[801:800];
    assign c[479:478] = {a[480], a[481]};
    assign c[481:480] = a[161:160];
    assign c[483:482] = a[803:802];
    assign c[485:484] = {a[482], a[483]};
    assign c[487:486] = a[163:162];
    assign c[489:488] = a[805:804];
    assign c[491:490] = {a[484], a[485]};
    assign c[493:492] = a[881:880];
    assign c[495:494] = a[561:560];
    assign c[497:496] = {a[486], a[487]};
    assign c[499:498] = a[883:882];
    assign c[501:500] = a[563:562];
    assign c[503:502] = {a[488], a[489]};
    assign c[505:504] = a[885:884];
    assign c[507:506] = a[565:564];
    assign c[509:508] = a[961:960];
    assign c[511:510] = a[887:886];
    assign c[513:512] = a[567:566];
    assign c[515:514] = a[963:962];
    assign c[517:516] = a[889:888];
    assign c[519:518] = a[569:568];
    assign c[521:520] = a[965:964];
    assign c[523:522] = {a[1136], a[1137]};
    assign c[525:524] = a[817:816];
    assign c[527:526] = {a[496], a[497]};
    assign c[529:528] = a[177:176];
    assign c[531:530] = a[819:818];
    assign c[533:532] = {a[498], a[499]};
    assign c[535:534] = a[179:178];
    assign c[537:536] = a[821:820];
    assign c[539:538] = {a[500], a[501]};
    assign c[541:540] = a[897:896];
    assign c[543:542] = a[577:576];
    assign c[545:544] = {a[502], a[503]};
    assign c[547:546] = a[899:898];
    assign c[549:548] = a[579:578];
    assign c[551:550] = {a[504], a[505]};
    assign c[553:552] = a[901:900];
    assign c[555:554] = a[581:580];
    assign c[557:556] = a[977:976];
    assign c[559:558] = a[903:902];
    assign c[561:560] = a[583:582];
    assign c[563:562] = a[979:978];
    assign c[565:564] = a[905:904];
    assign c[567:566] = a[585:584];
    assign c[569:568] = a[981:980];
    assign c[571:570] = {a[1152], a[1153]};
    assign c[573:572] = a[833:832];
    assign c[575:574] = {a[512], a[513]};
    assign c[577:576] = a[193:192];
    assign c[579:578] = a[835:834];
    assign c[581:580] = {a[514], a[515]};
    assign c[583:582] = a[195:194];
    assign c[585:584] = a[837:836];
    assign c[587:586] = {a[516], a[517]};
    assign c[589:588] = a[913:912];
    assign c[591:590] = a[593:592];
    assign c[593:592] = {a[518], a[519]};
    assign c[595:594] = a[915:914];
    assign c[597:596] = a[595:594];
    assign c[599:598] = {a[520], a[521]};
    assign c[601:600] = a[917:916];
    assign c[603:602] = a[597:596];
    assign c[605:604] = a[993:992];
    assign c[607:606] = a[919:918];
    assign c[609:608] = a[599:598];
    assign c[611:610] = a[995:994];
    assign c[613:612] = a[921:920];
    assign c[615:614] = a[601:600];
    assign c[617:616] = a[997:996];
    assign c[619:618] = {a[1168], a[1169]};
    assign c[621:620] = a[849:848];
    assign c[623:622] = {a[528], a[529]};
    assign c[625:624] = a[209:208];
    assign c[627:626] = a[851:850];
    assign c[629:628] = {a[530], a[531]};
    assign c[631:630] = a[211:210];
    assign c[633:632] = a[853:852];
    assign c[635:634] = {a[532], a[533]};
    assign c[637:636] = a[929:928];
    assign c[639:638] = a[609:608];
    assign c[641:640] = {a[534], a[535]};
    assign c[643:642] = a[931:930];
    assign c[645:644] = a[611:610];
    assign c[647:646] = {a[536], a[537]};
    assign c[649:648] = a[933:932];
    assign c[651:650] = a[613:612];
    assign c[653:652] = a[1009:1008];
    assign c[655:654] = a[935:934];
    assign c[657:656] = a[615:614];
    assign c[659:658] = a[1011:1010];
    assign c[661:660] = a[937:936];
    assign c[663:662] = a[617:616];
    assign c[665:664] = a[1013:1012];
    assign c[667:666] = {a[1184], a[1185]};
    assign c[669:668] = a[865:864];
    assign c[671:670] = {a[544], a[545]};
    assign c[673:672] = a[225:224];
    assign c[675:674] = a[867:866];
    assign c[677:676] = {a[546], a[547]};
    assign c[679:678] = a[227:226];
    assign c[681:680] = a[869:868];
    assign c[683:682] = {a[548], a[549]};
    assign c[685:684] = a[945:944];
    assign c[687:686] = a[625:624];
    assign c[689:688] = {a[550], a[551]};
    assign c[691:690] = a[947:946];
    assign c[693:692] = a[627:626];
    assign c[695:694] = {a[552], a[553]};
    assign c[697:696] = a[949:948];
    assign c[699:698] = a[629:628];
    assign c[701:700] = a[1025:1024];
    assign c[703:702] = a[951:950];
    assign c[705:704] = a[631:630];
    assign c[707:706] = a[1027:1026];
    assign c[709:708] = a[953:952];
    assign c[711:710] = a[633:632];
    assign c[713:712] = a[1029:1028];
    assign c[715:714] = a[955:954];
    assign c[717:716] = a[881:880];
    assign c[719:718] = {a[560], a[561]};
    assign c[721:720] = a[241:240];
    assign c[723:722] = a[883:882];
    assign c[725:724] = {a[562], a[563]};
    assign c[727:726] = a[243:242];
    assign c[729:728] = a[885:884];
    assign c[731:730] = {a[564], a[565]};
    assign c[733:732] = a[961:960];
    assign c[735:734] = a[641:640];
    assign c[737:736] = {a[566], a[567]};
    assign c[739:738] = a[963:962];
    assign c[741:740] = a[643:642];
    assign c[743:742] = {a[568], a[569]};
    assign c[745:744] = a[965:964];
    assign c[747:746] = a[645:644];
    assign c[749:748] = a[1041:1040];
    assign c[751:750] = a[967:966];
    assign c[753:752] = a[647:646];
    assign c[755:754] = a[1043:1042];
    assign c[757:756] = a[969:968];
    assign c[759:758] = a[649:648];
    assign c[761:760] = a[1045:1044];
    assign c[763:762] = a[971:970];
    assign c[765:764] = a[897:896];
    assign c[767:766] = {a[576], a[577]};
    assign c[769:768] = a[257:256];
    assign c[771:770] = a[899:898];
    assign c[773:772] = {a[578], a[579]};
    assign c[775:774] = a[259:258];
    assign c[777:776] = a[901:900];
    assign c[779:778] = {a[580], a[581]};
    assign c[781:780] = a[977:976];
    assign c[783:782] = a[657:656];
    assign c[785:784] = {a[582], a[583]};
    assign c[787:786] = a[979:978];
    assign c[789:788] = a[659:658];
    assign c[791:790] = {a[584], a[585]};
    assign c[793:792] = a[981:980];
    assign c[795:794] = a[661:660];
    assign c[797:796] = a[1057:1056];
    assign c[799:798] = a[983:982];
    assign c[801:800] = a[663:662];
    assign c[803:802] = a[1059:1058];
    assign c[805:804] = a[985:984];
    assign c[807:806] = a[665:664];
    assign c[809:808] = a[1061:1060];
    assign c[811:810] = a[987:986];
    assign c[813:812] = a[913:912];
    assign c[815:814] = {a[592], a[593]};
    assign c[817:816] = a[273:272];
    assign c[819:818] = a[915:914];
    assign c[821:820] = {a[594], a[595]};
    assign c[823:822] = a[275:274];
    assign c[825:824] = a[917:916];
    assign c[827:826] = {a[596], a[597]};
    assign c[829:828] = a[993:992];
    assign c[831:830] = a[673:672];
    assign c[833:832] = {a[598], a[599]};
    assign c[835:834] = a[995:994];
    assign c[837:836] = a[675:674];
    assign c[839:838] = {a[600], a[601]};
    assign c[841:840] = a[997:996];
    assign c[843:842] = a[677:676];
    assign c[845:844] = a[1073:1072];
    assign c[847:846] = a[999:998];
    assign c[849:848] = a[679:678];
    assign c[851:850] = a[1075:1074];
    assign c[853:852] = a[1001:1000];
    assign c[855:854] = a[681:680];
    assign c[857:856] = a[1077:1076];
    assign c[859:858] = a[1003:1002];
    assign c[861:860] = a[929:928];
    assign c[863:862] = {a[608], a[609]};
    assign c[865:864] = a[289:288];
    assign c[867:866] = a[931:930];
    assign c[869:868] = {a[610], a[611]};
    assign c[871:870] = a[291:290];
    assign c[873:872] = a[933:932];
    assign c[875:874] = {a[612], a[613]};
    assign c[877:876] = a[1009:1008];
    assign c[879:878] = a[689:688];
    assign c[881:880] = {a[614], a[615]};
    assign c[883:882] = a[1011:1010];
    assign c[885:884] = a[691:690];
    assign c[887:886] = {a[616], a[617]};
    assign c[889:888] = a[1013:1012];
    assign c[891:890] = a[693:692];
    assign c[893:892] = a[1089:1088];
    assign c[895:894] = a[1015:1014];
    assign c[897:896] = a[695:694];
    assign c[899:898] = a[1091:1090];
    assign c[901:900] = a[1017:1016];
    assign c[903:902] = a[697:696];
    assign c[905:904] = a[1093:1092];
    assign c[907:906] = a[1019:1018];
    assign c[909:908] = a[945:944];
    assign c[911:910] = {a[624], a[625]};
    assign c[913:912] = a[305:304];
    assign c[915:914] = a[947:946];
    assign c[917:916] = {a[626], a[627]};
    assign c[919:918] = a[307:306];
    assign c[921:920] = a[949:948];
    assign c[923:922] = {a[628], a[629]};
    assign c[925:924] = a[1025:1024];
    assign c[927:926] = a[705:704];
    assign c[929:928] = {a[630], a[631]};
    assign c[931:930] = a[1027:1026];
    assign c[933:932] = a[707:706];
    assign c[935:934] = {a[632], a[633]};
    assign c[937:936] = a[1029:1028];
    assign c[939:938] = a[709:708];
    assign c[941:940] = a[1105:1104];
    assign c[943:942] = a[1031:1030];
    assign c[945:944] = a[711:710];
    assign c[947:946] = a[1107:1106];
    assign c[949:948] = a[1033:1032];
    assign c[951:950] = a[713:712];
    assign c[953:952] = a[1109:1108];
    assign c[955:954] = a[1035:1034];
    assign c[957:956] = a[961:960];
    assign c[959:958] = {a[640], a[641]};
    assign c[961:960] = a[321:320];
    assign c[963:962] = a[963:962];
    assign c[965:964] = {a[642], a[643]};
    assign c[967:966] = a[323:322];
    assign c[969:968] = a[965:964];
    assign c[971:970] = {a[644], a[645]};
    assign c[973:972] = a[1041:1040];
    assign c[975:974] = a[721:720];
    assign c[977:976] = {a[646], a[647]};
    assign c[979:978] = a[1043:1042];
    assign c[981:980] = a[723:722];
    assign c[983:982] = {a[648], a[649]};
    assign c[985:984] = a[1045:1044];
    assign c[987:986] = a[725:724];
    assign c[989:988] = a[1121:1120];
    assign c[991:990] = a[1047:1046];
    assign c[993:992] = a[727:726];
    assign c[995:994] = a[1123:1122];
    assign c[997:996] = a[1049:1048];
    assign c[999:998] = a[729:728];
    assign c[1001:1000] = a[1125:1124];
    assign c[1003:1002] = a[1051:1050];
    assign c[1005:1004] = a[977:976];
    assign c[1007:1006] = {a[656], a[657]};
    assign c[1009:1008] = a[337:336];
    assign c[1011:1010] = a[979:978];
    assign c[1013:1012] = {a[658], a[659]};
    assign c[1015:1014] = a[339:338];
    assign c[1017:1016] = a[981:980];
    assign c[1019:1018] = {a[660], a[661]};
    assign c[1021:1020] = a[1057:1056];
    assign c[1023:1022] = a[737:736];
    assign c[1025:1024] = {a[662], a[663]};
    assign c[1027:1026] = a[1059:1058];
    assign c[1029:1028] = a[739:738];
    assign c[1031:1030] = {a[664], a[665]};
    assign c[1033:1032] = a[1061:1060];
    assign c[1035:1034] = a[741:740];
    assign c[1037:1036] = a[1137:1136];
    assign c[1039:1038] = a[1063:1062];
    assign c[1041:1040] = a[743:742];
    assign c[1043:1042] = a[1139:1138];
    assign c[1045:1044] = a[1065:1064];
    assign c[1047:1046] = a[745:744];
    assign c[1049:1048] = a[1141:1140];
    assign c[1051:1050] = a[1067:1066];
    assign c[1053:1052] = a[993:992];
    assign c[1055:1054] = {a[672], a[673]};
    assign c[1057:1056] = a[353:352];
    assign c[1059:1058] = a[995:994];
    assign c[1061:1060] = {a[674], a[675]};
    assign c[1063:1062] = a[355:354];
    assign c[1065:1064] = a[997:996];
    assign c[1067:1066] = {a[676], a[677]};
    assign c[1069:1068] = a[1073:1072];
    assign c[1071:1070] = a[753:752];
    assign c[1073:1072] = {a[678], a[679]};
    assign c[1075:1074] = a[1075:1074];
    assign c[1077:1076] = a[755:754];
    assign c[1079:1078] = {a[680], a[681]};
    assign c[1081:1080] = a[1077:1076];
    assign c[1083:1082] = a[757:756];
    assign c[1085:1084] = a[1153:1152];
    assign c[1087:1086] = a[1079:1078];
    assign c[1089:1088] = a[759:758];
    assign c[1091:1090] = a[1155:1154];
    assign c[1093:1092] = a[1081:1080];
    assign c[1095:1094] = a[761:760];
    assign c[1097:1096] = a[1157:1156];
    assign c[1099:1098] = a[1083:1082];
    assign c[1101:1100] = a[1009:1008];
    assign c[1103:1102] = {a[688], a[689]};
    assign c[1105:1104] = a[369:368];
    assign c[1107:1106] = a[1011:1010];
    assign c[1109:1108] = {a[690], a[691]};
    assign c[1111:1110] = a[371:370];
    assign c[1113:1112] = a[1013:1012];
    assign c[1115:1114] = {a[692], a[693]};
    assign c[1117:1116] = a[1089:1088];
    assign c[1119:1118] = a[769:768];
    assign c[1121:1120] = {a[694], a[695]};
    assign c[1123:1122] = a[1091:1090];
    assign c[1125:1124] = a[771:770];
    assign c[1127:1126] = {a[696], a[697]};
    assign c[1129:1128] = a[1093:1092];
    assign c[1131:1130] = a[773:772];
    assign c[1133:1132] = a[1169:1168];
    assign c[1135:1134] = a[1095:1094];
    assign c[1137:1136] = a[775:774];
    assign c[1139:1138] = a[1171:1170];
    assign c[1141:1140] = a[1097:1096];
    assign c[1143:1142] = a[777:776];
    assign c[1145:1144] = a[1173:1172];
    assign c[1147:1146] = a[1099:1098];
    assign c[1149:1148] = a[1025:1024];
    assign c[1151:1150] = {a[704], a[705]};
    assign c[1153:1152] = a[385:384];
    assign c[1155:1154] = a[1027:1026];
    assign c[1157:1156] = {a[706], a[707]};
    assign c[1159:1158] = a[387:386];
    assign c[1161:1160] = a[1029:1028];
    assign c[1163:1162] = {a[708], a[709]};
    assign c[1165:1164] = a[1105:1104];
    assign c[1167:1166] = a[785:784];
    assign c[1169:1168] = {a[710], a[711]};
    assign c[1171:1170] = a[1107:1106];
    assign c[1173:1172] = a[787:786];
    assign c[1175:1174] = {a[712], a[713]};
    assign c[1177:1176] = a[1109:1108];
    assign c[1179:1178] = a[789:788];
    assign c[1181:1180] = a[1185:1184];
    assign c[1183:1182] = a[1111:1110];
    assign c[1185:1184] = a[791:790];
endmodule
