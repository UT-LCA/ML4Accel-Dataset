
module dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2 (
        ap_clk,
        ap_rst,
        data_0_V_read,
        data_1_V_read,
        data_2_V_read,
        data_3_V_read,
        data_4_V_read,
        data_5_V_read,
        data_6_V_read,
        data_7_V_read,
        data_8_V_read,
        data_9_V_read,
        data_10_V_read,
        data_11_V_read,
        data_12_V_read,
        data_13_V_read,
        data_14_V_read,
        data_15_V_read,
        data_16_V_read,
        data_17_V_read,
        data_18_V_read,
        data_19_V_read,
        data_20_V_read,
        data_21_V_read,
        data_22_V_read,
        data_23_V_read,
        data_24_V_read,
        data_25_V_read,
        data_26_V_read,
        data_27_V_read,
        data_28_V_read,
        data_29_V_read,
        data_30_V_read,
        data_31_V_read,
        ap_return_0,
        ap_return_1,
        ap_return_2,
        ap_return_3,
        ap_return_4,
        ap_return_5,
        ap_return_6,
        ap_return_7,
        ap_return_8,
        ap_return_9,
        ap_return_10,
        ap_return_11,
        ap_return_12,
        ap_return_13,
        ap_return_14,
        ap_return_15,
        ap_return_16,
        ap_return_17,
        ap_return_18,
        ap_return_19,
        ap_return_20,
        ap_return_21,
        ap_return_22,
        ap_return_23,
        ap_return_24,
        ap_return_25,
        ap_return_26,
        ap_return_27,
        ap_return_28,
        ap_return_29,
        ap_return_30,
        ap_return_31,
        ap_ce
);


input   ap_clk;
input   ap_rst;
input  [15:0] data_0_V_read;
input  [15:0] data_1_V_read;
input  [15:0] data_2_V_read;
input  [15:0] data_3_V_read;
input  [15:0] data_4_V_read;
input  [15:0] data_5_V_read;
input  [15:0] data_6_V_read;
input  [15:0] data_7_V_read;
input  [15:0] data_8_V_read;
input  [15:0] data_9_V_read;
input  [15:0] data_10_V_read;
input  [15:0] data_11_V_read;
input  [15:0] data_12_V_read;
input  [15:0] data_13_V_read;
input  [15:0] data_14_V_read;
input  [15:0] data_15_V_read;
input  [15:0] data_16_V_read;
input  [15:0] data_17_V_read;
input  [15:0] data_18_V_read;
input  [15:0] data_19_V_read;
input  [15:0] data_20_V_read;
input  [15:0] data_21_V_read;
input  [15:0] data_22_V_read;
input  [15:0] data_23_V_read;
input  [15:0] data_24_V_read;
input  [15:0] data_25_V_read;
input  [15:0] data_26_V_read;
input  [15:0] data_27_V_read;
input  [15:0] data_28_V_read;
input  [15:0] data_29_V_read;
input  [15:0] data_30_V_read;
input  [15:0] data_31_V_read;
output  [15:0] ap_return_0;
output  [15:0] ap_return_1;
output  [15:0] ap_return_2;
output  [15:0] ap_return_3;
output  [15:0] ap_return_4;
output  [15:0] ap_return_5;
output  [15:0] ap_return_6;
output  [15:0] ap_return_7;
output  [15:0] ap_return_8;
output  [15:0] ap_return_9;
output  [15:0] ap_return_10;
output  [15:0] ap_return_11;
output  [15:0] ap_return_12;
output  [15:0] ap_return_13;
output  [15:0] ap_return_14;
output  [15:0] ap_return_15;
output  [15:0] ap_return_16;
output  [15:0] ap_return_17;
output  [15:0] ap_return_18;
output  [15:0] ap_return_19;
output  [15:0] ap_return_20;
output  [15:0] ap_return_21;
output  [15:0] ap_return_22;
output  [15:0] ap_return_23;
output  [15:0] ap_return_24;
output  [15:0] ap_return_25;
output  [15:0] ap_return_26;
output  [15:0] ap_return_27;
output  [15:0] ap_return_28;
output  [15:0] ap_return_29;
output  [15:0] ap_return_30;
output  [15:0] ap_return_31;
input   ap_ce;

reg[15:0] ap_return_0;
reg[15:0] ap_return_1;
reg[15:0] ap_return_2;
reg[15:0] ap_return_3;
reg[15:0] ap_return_4;
reg[15:0] ap_return_5;
reg[15:0] ap_return_6;
reg[15:0] ap_return_7;
reg[15:0] ap_return_8;
reg[15:0] ap_return_9;
reg[15:0] ap_return_10;
reg[15:0] ap_return_11;
reg[15:0] ap_return_12;
reg[15:0] ap_return_13;
reg[15:0] ap_return_14;
reg[15:0] ap_return_15;
reg[15:0] ap_return_16;
reg[15:0] ap_return_17;
reg[15:0] ap_return_18;
reg[15:0] ap_return_19;
reg[15:0] ap_return_20;
reg[15:0] ap_return_21;
reg[15:0] ap_return_22;
reg[15:0] ap_return_23;
reg[15:0] ap_return_24;
reg[15:0] ap_return_25;
reg[15:0] ap_return_26;
reg[15:0] ap_return_27;
reg[15:0] ap_return_28;
reg[15:0] ap_return_29;
reg[15:0] ap_return_30;
reg[15:0] ap_return_31;

reg   [15:0] data_31_V_read32_reg_4221;
wire    ap_block_state1_pp0_stage0_iter0;
wire    ap_block_state2_pp0_stage0_iter1;
wire    ap_block_state3_pp0_stage0_iter2;
wire    ap_block_state4_pp0_stage0_iter3;
wire    ap_block_state5_pp0_stage0_iter4;
wire    ap_block_state6_pp0_stage0_iter5;
wire    ap_block_state7_pp0_stage0_iter6;
wire    ap_block_state8_pp0_stage0_iter7;
wire    ap_block_state9_pp0_stage0_iter8;
wire    ap_block_state10_pp0_stage0_iter9;
wire    ap_block_pp0_stage0_11001;
reg   [15:0] data_31_V_read32_reg_4221_pp0_iter1_reg;
reg   [15:0] data_31_V_read32_reg_4221_pp0_iter2_reg;
reg   [15:0] data_31_V_read32_reg_4221_pp0_iter3_reg;
reg   [15:0] data_31_V_read32_reg_4221_pp0_iter4_reg;
reg   [15:0] data_31_V_read32_reg_4221_pp0_iter5_reg;
reg   [15:0] data_31_V_read32_reg_4221_pp0_iter6_reg;
reg   [15:0] data_31_V_read32_reg_4221_pp0_iter7_reg;
reg   [15:0] data_31_V_read32_reg_4221_pp0_iter8_reg;
reg   [15:0] data_30_V_read31_reg_4250;
reg   [15:0] data_30_V_read31_reg_4250_pp0_iter1_reg;
reg   [15:0] data_30_V_read31_reg_4250_pp0_iter2_reg;
reg   [15:0] data_30_V_read31_reg_4250_pp0_iter3_reg;
reg   [15:0] data_30_V_read31_reg_4250_pp0_iter4_reg;
reg   [15:0] data_30_V_read31_reg_4250_pp0_iter5_reg;
reg   [15:0] data_30_V_read31_reg_4250_pp0_iter6_reg;
reg   [15:0] data_30_V_read31_reg_4250_pp0_iter7_reg;
reg   [15:0] data_30_V_read31_reg_4250_pp0_iter8_reg;
reg   [15:0] data_29_V_read_7_reg_4279;
reg   [15:0] data_29_V_read_7_reg_4279_pp0_iter1_reg;
reg   [15:0] data_29_V_read_7_reg_4279_pp0_iter2_reg;
reg   [15:0] data_29_V_read_7_reg_4279_pp0_iter3_reg;
reg   [15:0] data_29_V_read_7_reg_4279_pp0_iter4_reg;
reg   [15:0] data_29_V_read_7_reg_4279_pp0_iter5_reg;
reg   [15:0] data_29_V_read_7_reg_4279_pp0_iter6_reg;
reg   [15:0] data_29_V_read_7_reg_4279_pp0_iter7_reg;
reg   [15:0] data_29_V_read_7_reg_4279_pp0_iter8_reg;
reg   [15:0] data_28_V_read_7_reg_4313;
reg   [15:0] data_28_V_read_7_reg_4313_pp0_iter1_reg;
reg   [15:0] data_28_V_read_7_reg_4313_pp0_iter2_reg;
reg   [15:0] data_28_V_read_7_reg_4313_pp0_iter3_reg;
reg   [15:0] data_28_V_read_7_reg_4313_pp0_iter4_reg;
reg   [15:0] data_28_V_read_7_reg_4313_pp0_iter5_reg;
reg   [15:0] data_28_V_read_7_reg_4313_pp0_iter6_reg;
reg   [15:0] data_28_V_read_7_reg_4313_pp0_iter7_reg;
reg   [15:0] data_28_V_read_7_reg_4313_pp0_iter8_reg;
reg   [15:0] data_27_V_read_8_reg_4342;
reg   [15:0] data_27_V_read_8_reg_4342_pp0_iter1_reg;
reg   [15:0] data_27_V_read_8_reg_4342_pp0_iter2_reg;
reg   [15:0] data_27_V_read_8_reg_4342_pp0_iter3_reg;
reg   [15:0] data_27_V_read_8_reg_4342_pp0_iter4_reg;
reg   [15:0] data_27_V_read_8_reg_4342_pp0_iter5_reg;
reg   [15:0] data_27_V_read_8_reg_4342_pp0_iter6_reg;
reg   [15:0] data_27_V_read_8_reg_4342_pp0_iter7_reg;
reg   [15:0] data_26_V_read27_reg_4365;
reg   [15:0] data_26_V_read27_reg_4365_pp0_iter1_reg;
reg   [15:0] data_26_V_read27_reg_4365_pp0_iter2_reg;
reg   [15:0] data_26_V_read27_reg_4365_pp0_iter3_reg;
reg   [15:0] data_26_V_read27_reg_4365_pp0_iter4_reg;
reg   [15:0] data_26_V_read27_reg_4365_pp0_iter5_reg;
reg   [15:0] data_26_V_read27_reg_4365_pp0_iter6_reg;
reg   [15:0] data_26_V_read27_reg_4365_pp0_iter7_reg;
reg   [15:0] data_25_V_read26_reg_4391;
reg   [15:0] data_25_V_read26_reg_4391_pp0_iter1_reg;
reg   [15:0] data_25_V_read26_reg_4391_pp0_iter2_reg;
reg   [15:0] data_25_V_read26_reg_4391_pp0_iter3_reg;
reg   [15:0] data_25_V_read26_reg_4391_pp0_iter4_reg;
reg   [15:0] data_25_V_read26_reg_4391_pp0_iter5_reg;
reg   [15:0] data_25_V_read26_reg_4391_pp0_iter6_reg;
reg   [15:0] data_25_V_read26_reg_4391_pp0_iter7_reg;
reg   [15:0] data_24_V_read25_reg_4421;
reg   [15:0] data_24_V_read25_reg_4421_pp0_iter1_reg;
reg   [15:0] data_24_V_read25_reg_4421_pp0_iter2_reg;
reg   [15:0] data_24_V_read25_reg_4421_pp0_iter3_reg;
reg   [15:0] data_24_V_read25_reg_4421_pp0_iter4_reg;
reg   [15:0] data_24_V_read25_reg_4421_pp0_iter5_reg;
reg   [15:0] data_24_V_read25_reg_4421_pp0_iter6_reg;
reg   [15:0] data_24_V_read25_reg_4421_pp0_iter7_reg;
reg   [15:0] data_23_V_read24_reg_4451;
reg   [15:0] data_23_V_read24_reg_4451_pp0_iter1_reg;
reg   [15:0] data_23_V_read24_reg_4451_pp0_iter2_reg;
reg   [15:0] data_23_V_read24_reg_4451_pp0_iter3_reg;
reg   [15:0] data_23_V_read24_reg_4451_pp0_iter4_reg;
reg   [15:0] data_23_V_read24_reg_4451_pp0_iter5_reg;
reg   [15:0] data_23_V_read24_reg_4451_pp0_iter6_reg;
reg   [15:0] data_23_V_read24_reg_4451_pp0_iter7_reg;
reg   [15:0] data_22_V_read23_reg_4483;
reg   [15:0] data_22_V_read23_reg_4483_pp0_iter1_reg;
reg   [15:0] data_22_V_read23_reg_4483_pp0_iter2_reg;
reg   [15:0] data_22_V_read23_reg_4483_pp0_iter3_reg;
reg   [15:0] data_22_V_read23_reg_4483_pp0_iter4_reg;
reg   [15:0] data_22_V_read23_reg_4483_pp0_iter5_reg;
reg   [15:0] data_22_V_read23_reg_4483_pp0_iter6_reg;
reg   [15:0] data_22_V_read23_reg_4483_pp0_iter7_reg;
reg   [15:0] data_21_V_read22_reg_4512;
reg   [15:0] data_21_V_read22_reg_4512_pp0_iter1_reg;
reg   [15:0] data_21_V_read22_reg_4512_pp0_iter2_reg;
reg   [15:0] data_21_V_read22_reg_4512_pp0_iter3_reg;
reg   [15:0] data_21_V_read22_reg_4512_pp0_iter4_reg;
reg   [15:0] data_21_V_read22_reg_4512_pp0_iter5_reg;
reg   [15:0] data_21_V_read22_reg_4512_pp0_iter6_reg;
reg   [15:0] data_20_V_read21_reg_4539;
reg   [15:0] data_20_V_read21_reg_4539_pp0_iter1_reg;
reg   [15:0] data_20_V_read21_reg_4539_pp0_iter2_reg;
reg   [15:0] data_20_V_read21_reg_4539_pp0_iter3_reg;
reg   [15:0] data_20_V_read21_reg_4539_pp0_iter4_reg;
reg   [15:0] data_20_V_read21_reg_4539_pp0_iter5_reg;
reg   [15:0] data_20_V_read21_reg_4539_pp0_iter6_reg;
reg   [15:0] data_19_V_read_7_reg_4567;
reg   [15:0] data_19_V_read_7_reg_4567_pp0_iter1_reg;
reg   [15:0] data_19_V_read_7_reg_4567_pp0_iter2_reg;
reg   [15:0] data_19_V_read_7_reg_4567_pp0_iter3_reg;
reg   [15:0] data_19_V_read_7_reg_4567_pp0_iter4_reg;
reg   [15:0] data_19_V_read_7_reg_4567_pp0_iter5_reg;
reg   [15:0] data_19_V_read_7_reg_4567_pp0_iter6_reg;
reg   [15:0] data_18_V_read_7_reg_4594;
reg   [15:0] data_18_V_read_7_reg_4594_pp0_iter1_reg;
reg   [15:0] data_18_V_read_7_reg_4594_pp0_iter2_reg;
reg   [15:0] data_18_V_read_7_reg_4594_pp0_iter3_reg;
reg   [15:0] data_18_V_read_7_reg_4594_pp0_iter4_reg;
reg   [15:0] data_18_V_read_7_reg_4594_pp0_iter5_reg;
reg   [15:0] data_18_V_read_7_reg_4594_pp0_iter6_reg;
reg   [15:0] data_17_V_read_8_reg_4621;
reg   [15:0] data_17_V_read_8_reg_4621_pp0_iter1_reg;
reg   [15:0] data_17_V_read_8_reg_4621_pp0_iter2_reg;
reg   [15:0] data_17_V_read_8_reg_4621_pp0_iter3_reg;
reg   [15:0] data_17_V_read_8_reg_4621_pp0_iter4_reg;
reg   [15:0] data_17_V_read_8_reg_4621_pp0_iter5_reg;
reg   [15:0] data_17_V_read_8_reg_4621_pp0_iter6_reg;
reg   [15:0] data_16_V_read17_reg_4650;
reg   [15:0] data_16_V_read17_reg_4650_pp0_iter1_reg;
reg   [15:0] data_16_V_read17_reg_4650_pp0_iter2_reg;
reg   [15:0] data_16_V_read17_reg_4650_pp0_iter3_reg;
reg   [15:0] data_16_V_read17_reg_4650_pp0_iter4_reg;
reg   [15:0] data_16_V_read17_reg_4650_pp0_iter5_reg;
reg   [15:0] data_15_V_read16_reg_4682;
reg   [15:0] data_15_V_read16_reg_4682_pp0_iter1_reg;
reg   [15:0] data_15_V_read16_reg_4682_pp0_iter2_reg;
reg   [15:0] data_15_V_read16_reg_4682_pp0_iter3_reg;
reg   [15:0] data_15_V_read16_reg_4682_pp0_iter4_reg;
reg   [15:0] data_15_V_read16_reg_4682_pp0_iter5_reg;
reg   [15:0] data_14_V_read15_reg_4714;
reg   [15:0] data_14_V_read15_reg_4714_pp0_iter1_reg;
reg   [15:0] data_14_V_read15_reg_4714_pp0_iter2_reg;
reg   [15:0] data_14_V_read15_reg_4714_pp0_iter3_reg;
reg   [15:0] data_14_V_read15_reg_4714_pp0_iter4_reg;
reg   [15:0] data_14_V_read15_reg_4714_pp0_iter5_reg;
reg   [15:0] data_13_V_read14_reg_4745;
reg   [15:0] data_13_V_read14_reg_4745_pp0_iter1_reg;
reg   [15:0] data_13_V_read14_reg_4745_pp0_iter2_reg;
reg   [15:0] data_13_V_read14_reg_4745_pp0_iter3_reg;
reg   [15:0] data_13_V_read14_reg_4745_pp0_iter4_reg;
reg   [15:0] data_13_V_read14_reg_4745_pp0_iter5_reg;
reg   [15:0] data_12_V_read13_reg_4778;
reg   [15:0] data_12_V_read13_reg_4778_pp0_iter1_reg;
reg   [15:0] data_12_V_read13_reg_4778_pp0_iter2_reg;
reg   [15:0] data_12_V_read13_reg_4778_pp0_iter3_reg;
reg   [15:0] data_12_V_read13_reg_4778_pp0_iter4_reg;
reg   [15:0] data_11_V_read12_reg_4808;
reg   [15:0] data_11_V_read12_reg_4808_pp0_iter1_reg;
reg   [15:0] data_11_V_read12_reg_4808_pp0_iter2_reg;
reg   [15:0] data_11_V_read12_reg_4808_pp0_iter3_reg;
reg   [15:0] data_11_V_read12_reg_4808_pp0_iter4_reg;
reg   [15:0] data_10_V_read11_reg_4832;
reg   [15:0] data_10_V_read11_reg_4832_pp0_iter1_reg;
reg   [15:0] data_10_V_read11_reg_4832_pp0_iter2_reg;
reg   [15:0] data_10_V_read11_reg_4832_pp0_iter3_reg;
reg   [15:0] data_10_V_read11_reg_4832_pp0_iter4_reg;
reg   [15:0] data_9_V_read_7_reg_4859;
reg   [15:0] data_9_V_read_7_reg_4859_pp0_iter1_reg;
reg   [15:0] data_9_V_read_7_reg_4859_pp0_iter2_reg;
reg   [15:0] data_9_V_read_7_reg_4859_pp0_iter3_reg;
reg   [15:0] data_9_V_read_7_reg_4859_pp0_iter4_reg;
reg   [15:0] data_8_V_read_7_reg_4887;
reg   [15:0] data_8_V_read_7_reg_4887_pp0_iter1_reg;
reg   [15:0] data_8_V_read_7_reg_4887_pp0_iter2_reg;
reg   [15:0] data_8_V_read_7_reg_4887_pp0_iter3_reg;
reg   [15:0] data_7_V_read_8_reg_4916;
reg   [15:0] data_7_V_read_8_reg_4916_pp0_iter1_reg;
reg   [15:0] data_7_V_read_8_reg_4916_pp0_iter2_reg;
reg   [15:0] data_7_V_read_8_reg_4916_pp0_iter3_reg;
reg   [15:0] data_6_V_read_8_reg_4944;
reg   [15:0] data_6_V_read_8_reg_4944_pp0_iter1_reg;
reg   [15:0] data_6_V_read_8_reg_4944_pp0_iter2_reg;
reg   [15:0] data_6_V_read_8_reg_4944_pp0_iter3_reg;
reg   [15:0] data_5_V_read_8_reg_4969;
reg   [15:0] data_5_V_read_8_reg_4969_pp0_iter1_reg;
reg   [15:0] data_5_V_read_8_reg_4969_pp0_iter2_reg;
reg   [15:0] data_5_V_read_8_reg_4969_pp0_iter3_reg;
reg   [15:0] data_4_V_read_9_reg_4998;
reg   [15:0] data_4_V_read_9_reg_4998_pp0_iter1_reg;
reg   [15:0] data_4_V_read_9_reg_4998_pp0_iter2_reg;
reg   [15:0] data_3_V_read_9_reg_5019;
reg   [15:0] data_3_V_read_9_reg_5019_pp0_iter1_reg;
reg   [15:0] data_3_V_read_9_reg_5019_pp0_iter2_reg;
reg   [15:0] data_2_V_read_9_reg_5035;
wire   [15:0] sub_ln703_fu_274_p2;
reg   [15:0] sub_ln703_reg_5046;
wire   [15:0] add_ln703_fu_280_p2;
reg   [15:0] add_ln703_reg_5052;
wire   [15:0] sub_ln703_73_fu_286_p2;
reg   [15:0] sub_ln703_73_reg_5059;
wire   [15:0] sub_ln703_74_fu_292_p2;
reg   [15:0] sub_ln703_74_reg_5065;
reg   [15:0] sub_ln703_74_reg_5065_pp0_iter2_reg;
wire   [15:0] sub_ln703_76_fu_300_p2;
reg   [15:0] sub_ln703_76_reg_5071;
reg   [15:0] sub_ln703_76_reg_5071_pp0_iter2_reg;
wire   [15:0] add_ln703_200_fu_304_p2;
reg   [15:0] add_ln703_200_reg_5077;
reg   [15:0] add_ln703_200_reg_5077_pp0_iter2_reg;
wire   [15:0] sub_ln703_77_fu_308_p2;
reg   [15:0] sub_ln703_77_reg_5084;
wire   [15:0] add_ln703_201_fu_312_p2;
reg   [15:0] add_ln703_201_reg_5090;
reg   [15:0] add_ln703_201_reg_5090_pp0_iter2_reg;
wire   [15:0] add_ln703_202_fu_316_p2;
reg   [15:0] add_ln703_202_reg_5096;
reg   [15:0] add_ln703_202_reg_5096_pp0_iter2_reg;
wire   [15:0] add_ln703_204_fu_320_p2;
reg   [15:0] add_ln703_204_reg_5101;
reg   [15:0] add_ln703_204_reg_5101_pp0_iter2_reg;
wire   [15:0] add_ln703_207_fu_325_p2;
reg   [15:0] add_ln703_207_reg_5107;
reg   [15:0] add_ln703_207_reg_5107_pp0_iter2_reg;
wire   [15:0] add_ln703_203_fu_329_p2;
reg   [15:0] add_ln703_203_reg_5113;
wire   [15:0] add_ln703_205_fu_333_p2;
reg   [15:0] add_ln703_205_reg_5119;
wire   [15:0] sub_ln703_79_fu_337_p2;
reg   [15:0] sub_ln703_79_reg_5125;
wire   [15:0] add_ln703_206_fu_341_p2;
reg   [15:0] add_ln703_206_reg_5131;
wire   [15:0] add_ln703_208_fu_345_p2;
reg   [15:0] add_ln703_208_reg_5137;
wire   [15:0] add_ln703_210_fu_349_p2;
reg   [15:0] add_ln703_210_reg_5143;
reg   [15:0] add_ln703_210_reg_5143_pp0_iter3_reg;
wire   [15:0] add_ln703_233_fu_353_p2;
reg   [15:0] add_ln703_233_reg_5149;
reg   [15:0] add_ln703_233_reg_5149_pp0_iter3_reg;
wire   [15:0] add_ln703_247_fu_357_p2;
reg   [15:0] add_ln703_247_reg_5159;
reg   [15:0] add_ln703_247_reg_5159_pp0_iter3_reg;
wire   [15:0] sub_ln703_89_fu_402_p2;
reg   [15:0] sub_ln703_89_reg_5166;
wire   [15:0] sub_ln703_91_fu_411_p2;
reg   [15:0] sub_ln703_91_reg_5172;
wire   [15:0] add_ln703_209_fu_416_p2;
reg   [15:0] add_ln703_209_reg_5178;
wire   [15:0] add_ln703_211_fu_420_p2;
reg   [15:0] add_ln703_211_reg_5184;
wire   [15:0] add_ln703_213_fu_429_p2;
reg   [15:0] add_ln703_213_reg_5189;
wire   [15:0] add_ln703_214_fu_433_p2;
reg   [15:0] add_ln703_214_reg_5194;
wire   [15:0] sub_ln703_93_fu_442_p2;
reg   [15:0] sub_ln703_93_reg_5200;
wire   [15:0] sub_ln703_94_fu_446_p2;
reg   [15:0] sub_ln703_94_reg_5205;
wire   [15:0] sub_ln703_96_fu_456_p2;
reg   [15:0] sub_ln703_96_reg_5210;
wire   [15:0] add_ln703_216_fu_461_p2;
reg   [15:0] add_ln703_216_reg_5215;
wire   [15:0] add_ln703_220_fu_484_p2;
reg   [15:0] add_ln703_220_reg_5221;
wire   [15:0] sub_ln703_105_fu_489_p2;
reg   [15:0] sub_ln703_105_reg_5226;
wire   [15:0] add_ln703_223_fu_507_p2;
reg   [15:0] add_ln703_223_reg_5231;
wire   [15:0] add_ln703_225_fu_513_p2;
reg   [15:0] add_ln703_225_reg_5237;
wire   [15:0] add_ln703_227_fu_522_p2;
reg   [15:0] add_ln703_227_reg_5242;
wire   [15:0] sub_ln703_113_fu_533_p2;
reg   [15:0] sub_ln703_113_reg_5247;
wire   [15:0] sub_ln703_114_fu_549_p2;
reg   [15:0] sub_ln703_114_reg_5253;
wire   [15:0] sub_ln703_117_fu_554_p2;
reg   [15:0] sub_ln703_117_reg_5259;
wire   [15:0] add_ln703_234_fu_564_p2;
reg   [15:0] add_ln703_234_reg_5264;
wire   [15:0] add_ln703_238_fu_569_p2;
reg   [15:0] add_ln703_238_reg_5269;
wire   [15:0] sub_ln703_126_fu_574_p2;
reg   [15:0] sub_ln703_126_reg_5274;
wire   [15:0] sub_ln703_129_fu_579_p2;
reg   [15:0] sub_ln703_129_reg_5279;
wire   [15:0] sub_ln703_133_fu_584_p2;
reg   [15:0] sub_ln703_133_reg_5284;
wire   [15:0] add_ln703_251_fu_589_p2;
reg   [15:0] add_ln703_251_reg_5289;
wire   [15:0] add_ln703_258_fu_593_p2;
reg   [15:0] add_ln703_258_reg_5295;
wire   [15:0] add_ln703_272_fu_597_p2;
reg   [15:0] add_ln703_272_reg_5304;
reg   [15:0] add_ln703_272_reg_5304_pp0_iter4_reg;
wire   [15:0] add_ln703_304_fu_601_p2;
reg   [15:0] add_ln703_304_reg_5314;
wire   [15:0] add_ln703_246_fu_787_p2;
reg   [15:0] add_ln703_246_reg_5320;
wire   [15:0] sub_ln703_138_fu_816_p2;
reg   [15:0] sub_ln703_138_reg_5325;
wire   [15:0] sub_ln703_141_fu_835_p2;
reg   [15:0] sub_ln703_141_reg_5330;
wire   [15:0] sub_ln703_143_fu_844_p2;
reg   [15:0] sub_ln703_143_reg_5335;
wire   [15:0] sub_ln703_144_fu_858_p2;
reg   [15:0] sub_ln703_144_reg_5340;
wire   [15:0] sub_ln703_145_fu_863_p2;
reg   [15:0] sub_ln703_145_reg_5345;
wire   [15:0] sub_ln703_149_fu_901_p2;
reg   [15:0] sub_ln703_149_reg_5350;
wire   [15:0] sub_ln703_154_fu_920_p2;
reg   [15:0] sub_ln703_154_reg_5355;
wire   [15:0] add_ln703_261_fu_955_p2;
reg   [15:0] add_ln703_261_reg_5360;
wire   [15:0] sub_ln703_161_fu_960_p2;
reg   [15:0] sub_ln703_161_reg_5365;
wire   [15:0] sub_ln703_162_fu_980_p2;
reg   [15:0] sub_ln703_162_reg_5370;
wire   [15:0] sub_ln703_166_fu_1000_p2;
reg   [15:0] sub_ln703_166_reg_5375;
wire   [15:0] sub_ln703_171_fu_1015_p2;
reg   [15:0] sub_ln703_171_reg_5380;
wire   [15:0] sub_ln703_173_fu_1025_p2;
reg   [15:0] sub_ln703_173_reg_5385;
wire   [15:0] sub_ln703_176_fu_1040_p2;
reg   [15:0] sub_ln703_176_reg_5390;
wire   [15:0] sub_ln703_180_fu_1045_p2;
reg   [15:0] sub_ln703_180_reg_5395;
wire   [15:0] sub_ln703_181_fu_1050_p2;
reg   [15:0] sub_ln703_181_reg_5400;
wire   [15:0] add_ln703_267_fu_1055_p2;
reg   [15:0] add_ln703_267_reg_5405;
wire   [15:0] sub_ln703_182_fu_1060_p2;
reg   [15:0] sub_ln703_182_reg_5410;
wire   [15:0] add_ln703_268_fu_1065_p2;
reg   [15:0] add_ln703_268_reg_5415;
wire   [15:0] add_ln703_274_fu_1089_p2;
reg   [15:0] add_ln703_274_reg_5420;
wire   [15:0] sub_ln703_185_fu_1095_p2;
reg   [15:0] sub_ln703_185_reg_5425;
wire   [15:0] add_ln703_276_fu_1100_p2;
reg   [15:0] add_ln703_276_reg_5430;
wire   [15:0] add_ln703_278_fu_1105_p2;
reg   [15:0] add_ln703_278_reg_5435;
wire   [15:0] sub_ln703_187_fu_1110_p2;
reg   [15:0] sub_ln703_187_reg_5440;
wire   [15:0] sub_ln703_189_fu_1115_p2;
reg   [15:0] sub_ln703_189_reg_5445;
wire   [15:0] sub_ln703_191_fu_1120_p2;
reg   [15:0] sub_ln703_191_reg_5450;
wire   [15:0] add_ln703_281_fu_1129_p2;
reg   [15:0] add_ln703_281_reg_5455;
wire   [15:0] add_ln703_283_fu_1140_p2;
reg   [15:0] add_ln703_283_reg_5460;
wire   [15:0] sub_ln703_198_fu_1146_p2;
reg   [15:0] sub_ln703_198_reg_5465;
wire   [15:0] sub_ln703_199_fu_1151_p2;
reg   [15:0] sub_ln703_199_reg_5470;
wire   [15:0] add_ln703_288_fu_1156_p2;
reg   [15:0] add_ln703_288_reg_5475;
wire   [15:0] add_ln703_309_fu_1179_p2;
reg   [15:0] add_ln703_309_reg_5484;
wire   [15:0] add_ln703_314_fu_1183_p2;
reg   [15:0] add_ln703_314_reg_5490;
wire   [15:0] add_ln703_316_fu_1187_p2;
reg   [15:0] add_ln703_316_reg_5496;
wire   [15:0] sub_ln703_246_fu_1193_p2;
reg   [15:0] sub_ln703_246_reg_5501;
wire   [15:0] add_ln703_323_fu_1198_p2;
reg   [15:0] add_ln703_323_reg_5506;
wire   [15:0] sub_ln703_200_fu_1326_p2;
reg   [15:0] sub_ln703_200_reg_5515;
wire   [15:0] sub_ln703_203_fu_1339_p2;
reg   [15:0] sub_ln703_203_reg_5520;
wire   [15:0] add_ln703_287_fu_1354_p2;
reg   [15:0] add_ln703_287_reg_5525;
wire   [15:0] add_ln703_291_fu_1371_p2;
reg   [15:0] add_ln703_291_reg_5530;
wire   [15:0] sub_ln703_207_fu_1384_p2;
reg   [15:0] sub_ln703_207_reg_5535;
wire   [15:0] sub_ln703_212_fu_1412_p2;
reg   [15:0] sub_ln703_212_reg_5540;
wire   [15:0] sub_ln703_215_fu_1441_p2;
reg   [15:0] sub_ln703_215_reg_5545;
wire   [15:0] add_ln703_301_fu_1494_p2;
reg   [15:0] add_ln703_301_reg_5550;
wire   [15:0] add_ln703_307_fu_1504_p2;
reg   [15:0] add_ln703_307_reg_5555;
wire   [15:0] sub_ln703_229_fu_1518_p2;
reg   [15:0] sub_ln703_229_reg_5560;
wire   [15:0] sub_ln703_237_fu_1571_p2;
reg   [15:0] sub_ln703_237_reg_5565;
wire   [15:0] sub_ln703_238_fu_1576_p2;
reg   [15:0] sub_ln703_238_reg_5570;
wire   [15:0] sub_ln703_252_fu_1616_p2;
reg   [15:0] sub_ln703_252_reg_5575;
wire   [15:0] sub_ln703_253_fu_1621_p2;
reg   [15:0] sub_ln703_253_reg_5580;
wire   [15:0] sub_ln703_254_fu_1626_p2;
reg   [15:0] sub_ln703_254_reg_5585;
wire   [15:0] add_ln703_321_fu_1636_p2;
reg   [15:0] add_ln703_321_reg_5590;
wire   [15:0] sub_ln703_257_fu_1641_p2;
reg   [15:0] sub_ln703_257_reg_5595;
wire   [15:0] sub_ln703_261_fu_1646_p2;
reg   [15:0] sub_ln703_261_reg_5600;
wire   [15:0] sub_ln703_262_fu_1651_p2;
reg   [15:0] sub_ln703_262_reg_5605;
wire   [15:0] sub_ln703_263_fu_1671_p2;
reg   [15:0] sub_ln703_263_reg_5610;
wire   [15:0] sub_ln703_265_fu_1676_p2;
reg   [15:0] sub_ln703_265_reg_5615;
wire   [15:0] sub_ln703_266_fu_1681_p2;
reg   [15:0] sub_ln703_266_reg_5620;
wire   [15:0] add_ln703_326_fu_1686_p2;
reg   [15:0] add_ln703_326_reg_5625;
wire   [15:0] sub_ln703_270_fu_1695_p2;
reg   [15:0] sub_ln703_270_reg_5630;
wire   [15:0] sub_ln703_272_fu_1700_p2;
reg   [15:0] sub_ln703_272_reg_5635;
wire   [15:0] add_ln703_330_fu_1710_p2;
reg   [15:0] add_ln703_330_reg_5640;
wire   [15:0] add_ln703_335_fu_1730_p2;
reg   [15:0] add_ln703_335_reg_5645;
wire   [15:0] sub_ln703_278_fu_1735_p2;
reg   [15:0] sub_ln703_278_reg_5650;
wire   [15:0] add_ln703_339_fu_1740_p2;
reg   [15:0] add_ln703_339_reg_5655;
wire   [15:0] add_ln703_343_fu_1745_p2;
reg   [15:0] add_ln703_343_reg_5660;
wire   [15:0] sub_ln703_289_fu_1750_p2;
reg   [15:0] sub_ln703_289_reg_5665;
wire   [15:0] sub_ln703_290_fu_1755_p2;
reg   [15:0] sub_ln703_290_reg_5670;
wire   [15:0] add_ln703_347_fu_1760_p2;
reg   [15:0] add_ln703_347_reg_5675;
wire   [15:0] add_ln703_357_fu_1764_p2;
reg   [15:0] add_ln703_357_reg_5683;
reg   [15:0] add_ln703_357_reg_5683_pp0_iter6_reg;
wire   [15:0] add_ln703_371_fu_1768_p2;
reg   [15:0] add_ln703_371_reg_5691;
wire   [15:0] add_ln703_384_fu_1772_p2;
reg   [15:0] add_ln703_384_reg_5701;
reg   [15:0] add_ln703_384_reg_5701_pp0_iter6_reg;
wire   [15:0] add_ln703_394_fu_1776_p2;
reg   [15:0] add_ln703_394_reg_5710;
reg   [15:0] add_ln703_394_reg_5710_pp0_iter6_reg;
wire   [15:0] add_ln703_404_fu_1780_p2;
reg   [15:0] add_ln703_404_reg_5718;
reg   [15:0] add_ln703_404_reg_5718_pp0_iter6_reg;
wire   [15:0] sub_ln703_276_fu_1918_p2;
reg   [15:0] sub_ln703_276_reg_5728;
wire   [15:0] sub_ln703_283_fu_1975_p2;
reg   [15:0] sub_ln703_283_reg_5733;
wire   [15:0] sub_ln703_288_fu_2003_p2;
reg   [15:0] sub_ln703_288_reg_5738;
wire   [15:0] add_ln703_353_fu_2060_p2;
reg   [15:0] add_ln703_353_reg_5743;
wire   [15:0] sub_ln703_300_fu_2075_p2;
reg   [15:0] sub_ln703_300_reg_5748;
wire   [15:0] add_ln703_354_fu_2080_p2;
reg   [15:0] add_ln703_354_reg_5753;
wire   [15:0] sub_ln703_302_fu_2089_p2;
reg   [15:0] sub_ln703_302_reg_5758;
wire   [15:0] sub_ln703_304_fu_2099_p2;
reg   [15:0] sub_ln703_304_reg_5763;
wire   [15:0] add_ln703_359_fu_2127_p2;
reg   [15:0] add_ln703_359_reg_5768;
wire   [15:0] sub_ln703_309_fu_2148_p2;
reg   [15:0] sub_ln703_309_reg_5773;
wire   [15:0] sub_ln703_311_fu_2173_p2;
reg   [15:0] sub_ln703_311_reg_5778;
wire   [15:0] sub_ln703_318_fu_2203_p2;
reg   [15:0] sub_ln703_318_reg_5783;
wire   [15:0] sub_ln703_321_fu_2218_p2;
reg   [15:0] sub_ln703_321_reg_5788;
wire   [15:0] add_ln703_372_fu_2228_p2;
reg   [15:0] add_ln703_372_reg_5793;
wire   [15:0] sub_ln703_323_fu_2233_p2;
reg   [15:0] sub_ln703_323_reg_5798;
wire   [15:0] sub_ln703_324_fu_2238_p2;
reg   [15:0] sub_ln703_324_reg_5803;
wire   [15:0] sub_ln703_325_fu_2243_p2;
reg   [15:0] sub_ln703_325_reg_5808;
wire   [15:0] sub_ln703_327_fu_2248_p2;
reg   [15:0] sub_ln703_327_reg_5813;
wire   [15:0] sub_ln703_328_fu_2253_p2;
reg   [15:0] sub_ln703_328_reg_5818;
wire   [15:0] sub_ln703_331_fu_2258_p2;
reg   [15:0] sub_ln703_331_reg_5823;
wire   [15:0] sub_ln703_332_fu_2273_p2;
reg   [15:0] sub_ln703_332_reg_5828;
wire   [15:0] add_ln703_377_fu_2283_p2;
reg   [15:0] add_ln703_377_reg_5833;
wire   [15:0] add_ln703_379_fu_2292_p2;
reg   [15:0] add_ln703_379_reg_5838;
wire   [15:0] sub_ln703_335_fu_2302_p2;
reg   [15:0] sub_ln703_335_reg_5843;
wire   [15:0] add_ln703_381_fu_2307_p2;
reg   [15:0] add_ln703_381_reg_5848;
wire   [15:0] sub_ln703_343_fu_2312_p2;
reg   [15:0] sub_ln703_343_reg_5853;
wire   [15:0] add_ln703_390_fu_2326_p2;
reg   [15:0] add_ln703_390_reg_5858;
wire   [15:0] sub_ln703_346_fu_2332_p2;
reg   [15:0] sub_ln703_346_reg_5863;
wire   [15:0] add_ln703_400_fu_2346_p2;
reg   [15:0] add_ln703_400_reg_5868;
wire   [15:0] add_ln703_413_fu_2361_p2;
reg   [15:0] add_ln703_413_reg_5873;
wire   [15:0] add_ln703_415_fu_2372_p2;
reg   [15:0] add_ln703_415_reg_5878;
wire   [15:0] add_ln703_427_fu_2383_p2;
reg   [15:0] add_ln703_427_reg_5883;
wire   [15:0] add_ln703_428_fu_2389_p2;
reg   [15:0] add_ln703_428_reg_5888;
wire   [15:0] add_ln703_435_fu_2393_p2;
reg   [15:0] add_ln703_435_reg_5894;
wire   [15:0] add_ln703_446_fu_2397_p2;
reg   [15:0] add_ln703_446_reg_5901;
wire   [15:0] add_ln703_462_fu_2401_p2;
reg   [15:0] add_ln703_462_reg_5909;
reg   [15:0] add_ln703_462_reg_5909_pp0_iter7_reg;
reg   [15:0] add_ln703_462_reg_5909_pp0_iter8_reg;
wire   [15:0] sub_ln703_356_fu_2603_p2;
reg   [15:0] sub_ln703_356_reg_5921;
wire   [15:0] sub_ln703_357_fu_2608_p2;
reg   [15:0] sub_ln703_357_reg_5926;
wire   [15:0] add_ln703_402_fu_2631_p2;
reg   [15:0] add_ln703_402_reg_5931;
wire   [15:0] sub_ln703_361_fu_2636_p2;
reg   [15:0] sub_ln703_361_reg_5936;
wire   [15:0] sub_ln703_366_fu_2684_p2;
reg   [15:0] sub_ln703_366_reg_5941;
wire   [15:0] sub_ln703_369_fu_2699_p2;
reg   [15:0] sub_ln703_369_reg_5946;
wire   [15:0] add_ln703_410_fu_2709_p2;
reg   [15:0] add_ln703_410_reg_5951;
wire   [15:0] sub_ln703_374_fu_2728_p2;
reg   [15:0] sub_ln703_374_reg_5956;
wire   [15:0] add_ln703_418_fu_2741_p2;
reg   [15:0] add_ln703_418_reg_5961;
wire   [15:0] sub_ln703_375_fu_2747_p2;
reg   [15:0] sub_ln703_375_reg_5966;
wire   [15:0] sub_ln703_379_fu_2781_p2;
reg   [15:0] sub_ln703_379_reg_5971;
wire   [15:0] sub_ln703_381_fu_2791_p2;
reg   [15:0] sub_ln703_381_reg_5976;
wire   [15:0] add_ln703_424_fu_2806_p2;
reg   [15:0] add_ln703_424_reg_5981;
wire   [15:0] sub_ln703_385_fu_2811_p2;
reg   [15:0] sub_ln703_385_reg_5986;
wire   [15:0] sub_ln703_386_fu_2816_p2;
reg   [15:0] sub_ln703_386_reg_5991;
wire   [15:0] sub_ln703_389_fu_2839_p2;
reg   [15:0] sub_ln703_389_reg_5996;
wire   [15:0] sub_ln703_392_fu_2848_p2;
reg   [15:0] sub_ln703_392_reg_6001;
wire   [15:0] sub_ln703_397_fu_2863_p2;
reg   [15:0] sub_ln703_397_reg_6006;
wire   [15:0] add_ln703_434_fu_2873_p2;
reg   [15:0] add_ln703_434_reg_6011;
wire   [15:0] sub_ln703_402_fu_2878_p2;
reg   [15:0] sub_ln703_402_reg_6016;
wire   [15:0] add_ln703_436_fu_2883_p2;
reg   [15:0] add_ln703_436_reg_6021;
wire   [15:0] sub_ln703_408_fu_2893_p2;
reg   [15:0] sub_ln703_408_reg_6026;
wire   [15:0] sub_ln703_409_fu_2898_p2;
reg   [15:0] sub_ln703_409_reg_6031;
wire   [15:0] sub_ln703_411_fu_2903_p2;
reg   [15:0] sub_ln703_411_reg_6036;
wire   [15:0] add_ln703_442_fu_2917_p2;
reg   [15:0] add_ln703_442_reg_6041;
wire   [15:0] sub_ln703_416_fu_2923_p2;
reg   [15:0] sub_ln703_416_reg_6046;
wire   [15:0] add_ln703_444_fu_2928_p2;
reg   [15:0] add_ln703_444_reg_6051;
wire   [15:0] add_ln703_447_fu_2933_p2;
reg   [15:0] add_ln703_447_reg_6056;
wire   [15:0] sub_ln703_426_fu_2938_p2;
reg   [15:0] sub_ln703_426_reg_6061;
wire   [15:0] add_ln703_451_fu_2943_p2;
reg   [15:0] add_ln703_451_reg_6066;
reg   [15:0] add_ln703_451_reg_6066_pp0_iter8_reg;
wire   [15:0] add_ln703_480_fu_2961_p2;
reg   [15:0] add_ln703_480_reg_6072;
reg   [15:0] add_ln703_480_reg_6072_pp0_iter8_reg;
wire   [15:0] add_ln703_482_fu_2967_p2;
reg   [15:0] add_ln703_482_reg_6077;
wire   [15:0] add_ln703_491_fu_2971_p2;
reg   [15:0] add_ln703_491_reg_6087;
reg   [15:0] add_ln703_491_reg_6087_pp0_iter8_reg;
wire   [15:0] add_ln703_509_fu_2976_p2;
reg   [15:0] add_ln703_509_reg_6092;
reg   [15:0] add_ln703_509_reg_6092_pp0_iter8_reg;
wire   [15:0] add_ln703_516_fu_2980_p2;
reg   [15:0] add_ln703_516_reg_6103;
reg   [15:0] add_ln703_516_reg_6103_pp0_iter8_reg;
wire   [15:0] sub_ln703_428_fu_3163_p2;
reg   [15:0] sub_ln703_428_reg_6108;
wire   [15:0] sub_ln703_434_fu_3199_p2;
reg   [15:0] sub_ln703_434_reg_6113;
wire   [15:0] sub_ln703_448_fu_3308_p2;
reg   [15:0] sub_ln703_448_reg_6118;
wire   [15:0] sub_ln703_450_fu_3318_p2;
reg   [15:0] sub_ln703_450_reg_6123;
wire   [15:0] add_ln703_463_fu_3328_p2;
reg   [15:0] add_ln703_463_reg_6128;
wire   [15:0] add_ln703_464_fu_3333_p2;
reg   [15:0] add_ln703_464_reg_6133;
wire   [15:0] add_ln703_465_fu_3338_p2;
reg   [15:0] add_ln703_465_reg_6138;
wire   [15:0] sub_ln703_451_fu_3343_p2;
reg   [15:0] sub_ln703_451_reg_6143;
wire   [15:0] sub_ln703_452_fu_3348_p2;
reg   [15:0] sub_ln703_452_reg_6148;
wire   [15:0] sub_ln703_453_fu_3353_p2;
reg   [15:0] sub_ln703_453_reg_6153;
wire   [15:0] add_ln703_467_fu_3363_p2;
reg   [15:0] add_ln703_467_reg_6158;
wire   [15:0] sub_ln703_454_fu_3368_p2;
reg   [15:0] sub_ln703_454_reg_6163;
wire   [15:0] sub_ln703_455_fu_3373_p2;
reg   [15:0] sub_ln703_455_reg_6168;
wire   [15:0] add_ln703_468_fu_3378_p2;
reg   [15:0] add_ln703_468_reg_6173;
wire   [15:0] sub_ln703_456_fu_3388_p2;
reg   [15:0] sub_ln703_456_reg_6178;
wire   [15:0] sub_ln703_457_fu_3393_p2;
reg   [15:0] sub_ln703_457_reg_6183;
wire   [15:0] add_ln703_471_fu_3403_p2;
reg   [15:0] add_ln703_471_reg_6188;
wire   [15:0] sub_ln703_458_fu_3408_p2;
reg   [15:0] sub_ln703_458_reg_6193;
wire   [15:0] sub_ln703_459_fu_3418_p2;
reg   [15:0] sub_ln703_459_reg_6198;
wire   [15:0] add_ln703_475_fu_3432_p2;
reg   [15:0] add_ln703_475_reg_6203;
wire   [15:0] sub_ln703_461_fu_3438_p2;
reg   [15:0] sub_ln703_461_reg_6208;
wire   [15:0] add_ln703_483_fu_3448_p2;
reg   [15:0] add_ln703_483_reg_6213;
wire   [15:0] sub_ln703_469_fu_3463_p2;
reg   [15:0] sub_ln703_469_reg_6218;
wire   [15:0] add_ln703_492_fu_3478_p2;
reg   [15:0] add_ln703_492_reg_6223;
wire   [15:0] sub_ln703_474_fu_3482_p2;
reg   [15:0] sub_ln703_474_reg_6229;
wire   [15:0] add_ln703_496_fu_3497_p2;
reg   [15:0] add_ln703_496_reg_6234;
wire   [15:0] add_ln703_497_fu_3501_p2;
reg   [15:0] add_ln703_497_reg_6239;
wire   [15:0] sub_ln703_486_fu_3507_p2;
reg   [15:0] sub_ln703_486_reg_6244;
wire   [15:0] sub_ln703_487_fu_3512_p2;
reg   [15:0] sub_ln703_487_reg_6249;
wire   [15:0] sub_ln703_491_fu_3517_p2;
reg   [15:0] sub_ln703_491_reg_6254;
wire   [15:0] sub_ln703_500_fu_3522_p2;
reg   [15:0] sub_ln703_500_reg_6259;
wire   [15:0] add_ln703_510_fu_3527_p2;
reg   [15:0] add_ln703_510_reg_6264;
wire    ap_block_pp0_stage0;
wire   [15:0] sub_ln703_75_fu_296_p2;
wire   [15:0] sub_ln703_78_fu_361_p2;
wire   [15:0] sub_ln703_80_fu_365_p2;
wire   [15:0] sub_ln703_81_fu_369_p2;
wire   [15:0] sub_ln703_82_fu_373_p2;
wire   [15:0] sub_ln703_84_fu_381_p2;
wire   [15:0] sub_ln703_86_fu_389_p2;
wire   [15:0] sub_ln703_87_fu_393_p2;
wire   [15:0] sub_ln703_88_fu_398_p2;
wire   [15:0] sub_ln703_90_fu_406_p2;
wire   [15:0] add_ln703_212_fu_425_p2;
wire   [15:0] sub_ln703_92_fu_437_p2;
wire   [15:0] add_ln703_222_fu_503_p2;
wire   [15:0] sub_ln703_85_fu_385_p2;
wire   [15:0] sub_ln703_98_fu_466_p2;
wire   [15:0] add_ln703_226_fu_518_p2;
wire   [15:0] add_ln703_217_fu_470_p2;
wire   [15:0] add_ln703_218_fu_474_p2;
wire   [15:0] sub_ln703_83_fu_377_p2;
wire   [15:0] add_ln703_230_fu_538_p2;
wire   [15:0] add_ln703_219_fu_479_p2;
wire   [15:0] sub_ln703_106_fu_494_p2;
wire   [15:0] add_ln703_221_fu_499_p2;
wire   [15:0] sub_ln703_95_fu_451_p2;
wire   [15:0] sub_ln703_112_fu_528_p2;
wire   [15:0] add_ln703_231_fu_543_p2;
wire   [15:0] sub_ln703_118_fu_559_p2;
wire   [15:0] add_ln703_215_fu_605_p2;
wire   [15:0] sub_ln703_97_fu_609_p2;
wire   [15:0] sub_ln703_99_fu_613_p2;
wire   [15:0] sub_ln703_100_fu_617_p2;
wire   [15:0] sub_ln703_101_fu_621_p2;
wire   [15:0] sub_ln703_103_fu_629_p2;
wire   [15:0] sub_ln703_108_fu_641_p2;
wire   [15:0] add_ln703_224_fu_645_p2;
wire   [15:0] sub_ln703_110_fu_654_p2;
wire   [15:0] sub_ln703_111_fu_658_p2;
wire   [15:0] add_ln703_228_fu_663_p2;
wire   [15:0] add_ln703_229_fu_668_p2;
wire   [15:0] add_ln703_232_fu_673_p2;
wire   [15:0] sub_ln703_102_fu_625_p2;
wire   [15:0] sub_ln703_115_fu_678_p2;
wire   [15:0] sub_ln703_116_fu_683_p2;
wire   [15:0] sub_ln703_107_fu_637_p2;
wire   [15:0] add_ln703_243_fu_774_p2;
wire   [15:0] sub_ln703_119_fu_687_p2;
wire   [15:0] sub_ln703_121_fu_696_p2;
wire   [15:0] sub_ln703_109_fu_649_p2;
wire   [15:0] add_ln703_235_fu_701_p2;
wire   [15:0] sub_ln703_122_fu_705_p2;
wire   [15:0] add_ln703_236_fu_710_p2;
wire   [15:0] add_ln703_237_fu_715_p2;
wire   [15:0] sub_ln703_123_fu_719_p2;
wire   [15:0] sub_ln703_125_fu_727_p2;
wire   [15:0] sub_ln703_128_fu_736_p2;
wire   [15:0] add_ln703_250_fu_849_p2;
wire   [15:0] add_ln703_239_fu_750_p2;
wire   [15:0] add_ln703_240_fu_755_p2;
wire   [15:0] sub_ln703_132_fu_760_p2;
wire   [15:0] add_ln703_253_fu_873_p2;
wire   [15:0] add_ln703_241_fu_765_p2;
wire   [15:0] add_ln703_255_fu_887_p2;
wire   [15:0] add_ln703_242_fu_769_p2;
wire   [15:0] add_ln703_244_fu_778_p2;
wire   [15:0] add_ln703_245_fu_783_p2;
wire   [15:0] sub_ln703_134_fu_792_p2;
wire   [15:0] add_ln703_248_fu_801_p2;
wire   [15:0] sub_ln703_139_fu_821_p2;
wire   [15:0] sub_ln703_140_fu_826_p2;
wire   [15:0] add_ln703_249_fu_830_p2;
wire   [15:0] sub_ln703_124_fu_723_p2;
wire   [15:0] sub_ln703_142_fu_840_p2;
wire   [15:0] sub_ln703_127_fu_732_p2;
wire   [15:0] sub_ln703_131_fu_745_p2;
wire   [15:0] add_ln703_252_fu_853_p2;
wire   [15:0] sub_ln703_104_fu_633_p2;
wire   [15:0] add_ln703_263_fu_970_p2;
wire   [15:0] add_ln703_262_fu_965_p2;
wire   [15:0] sub_ln703_146_fu_868_p2;
wire   [15:0] add_ln703_254_fu_877_p2;
wire   [15:0] sub_ln703_147_fu_882_p2;
wire   [15:0] add_ln703_256_fu_891_p2;
wire   [15:0] sub_ln703_148_fu_896_p2;
wire   [15:0] sub_ln703_151_fu_911_p2;
wire   [15:0] sub_ln703_153_fu_915_p2;
wire   [15:0] add_ln703_257_fu_925_p2;
wire   [15:0] sub_ln703_156_fu_930_p2;
wire   [15:0] sub_ln703_157_fu_935_p2;
wire   [15:0] add_ln703_259_fu_940_p2;
wire   [15:0] sub_ln703_159_fu_945_p2;
wire   [15:0] add_ln703_260_fu_950_p2;
wire   [15:0] add_ln703_264_fu_974_p2;
wire   [15:0] sub_ln703_163_fu_985_p2;
wire   [15:0] sub_ln703_164_fu_990_p2;
wire   [15:0] sub_ln703_165_fu_995_p2;
wire   [15:0] sub_ln703_150_fu_906_p2;
wire   [15:0] sub_ln703_168_fu_1005_p2;
wire   [15:0] sub_ln703_120_fu_691_p2;
wire   [15:0] add_ln703_273_fu_1085_p2;
wire   [15:0] add_ln703_271_fu_1080_p2;
wire   [15:0] add_ln703_265_fu_1010_p2;
wire   [15:0] sub_ln703_136_fu_806_p2;
wire   [15:0] sub_ln703_137_fu_811_p2;
wire   [15:0] sub_ln703_172_fu_1020_p2;
wire   [15:0] sub_ln703_174_fu_1030_p2;
wire   [15:0] sub_ln703_175_fu_1035_p2;
wire   [15:0] add_ln703_280_fu_1125_p2;
wire   [15:0] sub_ln703_130_fu_741_p2;
wire   [15:0] add_ln703_282_fu_1135_p2;
wire   [15:0] add_ln703_269_fu_1069_p2;
wire   [15:0] sub_ln703_184_fu_1075_p2;
wire   [15:0] add_ln703_302_fu_1160_p2;
wire   [15:0] add_ln703_305_fu_1169_p2;
wire   [15:0] add_ln703_303_fu_1164_p2;
wire   [15:0] sub_ln703_135_fu_796_p2;
wire   [15:0] add_ln703_306_fu_1173_p2;
wire   [15:0] sub_ln703_152_fu_1202_p2;
wire   [15:0] sub_ln703_155_fu_1206_p2;
wire   [15:0] sub_ln703_158_fu_1210_p2;
wire   [15:0] sub_ln703_160_fu_1214_p2;
wire   [15:0] sub_ln703_167_fu_1218_p2;
wire   [15:0] sub_ln703_169_fu_1222_p2;
wire   [15:0] sub_ln703_170_fu_1227_p2;
wire   [15:0] add_ln703_266_fu_1232_p2;
wire   [15:0] sub_ln703_177_fu_1237_p2;
wire   [15:0] sub_ln703_179_fu_1246_p2;
wire   [15:0] add_ln703_284_fu_1296_p2;
wire   [15:0] sub_ln703_183_fu_1250_p2;
wire   [15:0] add_ln703_270_fu_1255_p2;
wire   [15:0] add_ln703_275_fu_1260_p2;
wire   [15:0] add_ln703_277_fu_1264_p2;
wire   [15:0] add_ln703_279_fu_1268_p2;
wire   [15:0] sub_ln703_186_fu_1272_p2;
wire   [15:0] sub_ln703_190_fu_1281_p2;
wire   [15:0] sub_ln703_192_fu_1286_p2;
wire   [15:0] sub_ln703_178_fu_1242_p2;
wire   [15:0] sub_ln703_193_fu_1291_p2;
wire   [15:0] add_ln703_285_fu_1300_p2;
wire   [15:0] add_ln703_286_fu_1305_p2;
wire   [15:0] sub_ln703_194_fu_1309_p2;
wire   [15:0] sub_ln703_195_fu_1313_p2;
wire   [15:0] sub_ln703_196_fu_1317_p2;
wire   [15:0] add_ln703_296_fu_1432_p2;
wire   [15:0] sub_ln703_197_fu_1321_p2;
wire   [15:0] sub_ln703_202_fu_1335_p2;
wire   [15:0] sub_ln703_204_fu_1344_p2;
wire   [15:0] sub_ln703_205_fu_1349_p2;
wire   [15:0] add_ln703_289_fu_1359_p2;
wire   [15:0] sub_ln703_206_fu_1363_p2;
wire   [15:0] add_ln703_290_fu_1367_p2;
wire   [15:0] add_ln703_292_fu_1376_p2;
wire   [15:0] add_ln703_293_fu_1380_p2;
wire   [15:0] sub_ln703_208_fu_1389_p2;
wire   [15:0] add_ln703_294_fu_1397_p2;
wire   [15:0] sub_ln703_210_fu_1402_p2;
wire   [15:0] add_ln703_308_fu_1509_p2;
wire   [15:0] sub_ln703_211_fu_1407_p2;
wire   [15:0] add_ln703_311_fu_1523_p2;
wire   [15:0] sub_ln703_213_fu_1417_p2;
wire   [15:0] add_ln703_295_fu_1427_p2;
wire   [15:0] add_ln703_297_fu_1436_p2;
wire   [15:0] sub_ln703_217_fu_1450_p2;
wire   [15:0] sub_ln703_201_fu_1331_p2;
wire   [15:0] add_ln703_298_fu_1454_p2;
wire   [15:0] add_ln703_317_fu_1562_p2;
wire   [15:0] sub_ln703_220_fu_1459_p2;
wire   [15:0] add_ln703_299_fu_1464_p2;
wire   [15:0] sub_ln703_222_fu_1469_p2;
wire   [15:0] add_ln703_300_fu_1474_p2;
wire   [15:0] sub_ln703_223_fu_1479_p2;
wire   [15:0] sub_ln703_225_fu_1484_p2;
wire   [15:0] sub_ln703_226_fu_1489_p2;
wire   [15:0] add_ln703_310_fu_1513_p2;
wire   [15:0] add_ln703_312_fu_1527_p2;
wire   [15:0] add_ln703_313_fu_1532_p2;
wire   [15:0] sub_ln703_231_fu_1537_p2;
wire   [15:0] sub_ln703_232_fu_1542_p2;
wire   [15:0] add_ln703_315_fu_1552_p2;
wire   [15:0] sub_ln703_236_fu_1557_p2;
wire   [15:0] add_ln703_318_fu_1566_p2;
wire   [15:0] sub_ln703_240_fu_1581_p2;
wire   [15:0] sub_ln703_241_fu_1586_p2;
wire   [15:0] sub_ln703_188_fu_1277_p2;
wire   [15:0] add_ln703_324_fu_1661_p2;
wire   [15:0] add_ln703_322_fu_1656_p2;
wire   [15:0] add_ln703_319_fu_1591_p2;
wire   [15:0] sub_ln703_242_fu_1596_p2;
wire   [15:0] sub_ln703_243_fu_1601_p2;
wire   [15:0] sub_ln703_228_fu_1499_p2;
wire   [15:0] sub_ln703_248_fu_1606_p2;
wire   [15:0] sub_ln703_251_fu_1611_p2;
wire   [15:0] sub_ln703_214_fu_1422_p2;
wire   [15:0] add_ln703_329_fu_1705_p2;
wire   [15:0] sub_ln703_216_fu_1446_p2;
wire   [15:0] add_ln703_332_fu_1715_p2;
wire   [15:0] sub_ln703_234_fu_1547_p2;
wire   [15:0] sub_ln703_256_fu_1631_p2;
wire   [15:0] add_ln703_325_fu_1665_p2;
wire   [15:0] sub_ln703_209_fu_1393_p2;
wire   [15:0] sub_ln703_268_fu_1691_p2;
wire   [15:0] add_ln703_333_fu_1720_p2;
wire   [15:0] add_ln703_334_fu_1725_p2;
wire   [15:0] sub_ln703_218_fu_1784_p2;
wire   [15:0] sub_ln703_221_fu_1792_p2;
wire   [15:0] sub_ln703_224_fu_1796_p2;
wire   [15:0] sub_ln703_227_fu_1800_p2;
wire   [15:0] sub_ln703_230_fu_1804_p2;
wire   [15:0] sub_ln703_233_fu_1808_p2;
wire   [15:0] sub_ln703_239_fu_1817_p2;
wire   [15:0] add_ln703_320_fu_1822_p2;
wire   [15:0] sub_ln703_245_fu_1832_p2;
wire   [15:0] sub_ln703_247_fu_1836_p2;
wire   [15:0] sub_ln703_249_fu_1840_p2;
wire   [15:0] sub_ln703_250_fu_1844_p2;
wire   [15:0] sub_ln703_255_fu_1849_p2;
wire   [15:0] sub_ln703_258_fu_1854_p2;
wire   [15:0] sub_ln703_260_fu_1862_p2;
wire   [15:0] add_ln703_340_fu_1943_p2;
wire   [15:0] add_ln703_341_fu_1947_p2;
wire   [15:0] sub_ln703_269_fu_1877_p2;
wire   [15:0] sub_ln703_271_fu_1882_p2;
wire   [15:0] add_ln703_327_fu_1887_p2;
wire   [15:0] add_ln703_328_fu_1892_p2;
wire   [15:0] sub_ln703_273_fu_1896_p2;
wire   [15:0] add_ln703_331_fu_1900_p2;
wire   [15:0] sub_ln703_274_fu_1904_p2;
wire   [15:0] sub_ln703_275_fu_1909_p2;
wire   [15:0] sub_ln703_219_fu_1788_p2;
wire   [15:0] add_ln703_350_fu_2026_p2;
wire   [15:0] add_ln703_349_fu_2021_p2;
wire   [15:0] add_ln703_336_fu_1913_p2;
wire   [15:0] add_ln703_337_fu_1923_p2;
wire   [15:0] sub_ln703_277_fu_1927_p2;
wire   [15:0] sub_ln703_279_fu_1931_p2;
wire   [15:0] sub_ln703_264_fu_1867_p2;
wire   [15:0] sub_ln703_280_fu_1935_p2;
wire   [15:0] add_ln703_338_fu_1939_p2;
wire   [15:0] add_ln703_342_fu_1952_p2;
wire   [15:0] sub_ln703_281_fu_1957_p2;
wire   [15:0] sub_ln703_282_fu_1961_p2;
wire   [15:0] add_ln703_344_fu_1966_p2;
wire   [15:0] add_ln703_345_fu_1970_p2;
wire   [15:0] sub_ln703_286_fu_1989_p2;
wire   [15:0] add_ln703_346_fu_1993_p2;
wire   [15:0] sub_ln703_235_fu_1812_p2;
wire   [15:0] add_ln703_358_fu_2123_p2;
wire   [15:0] add_ln703_356_fu_2118_p2;
wire   [15:0] sub_ln703_291_fu_2008_p2;
wire   [15:0] sub_ln703_292_fu_2012_p2;
wire   [15:0] add_ln703_348_fu_2017_p2;
wire   [15:0] add_ln703_351_fu_2030_p2;
wire   [15:0] sub_ln703_259_fu_1858_p2;
wire   [15:0] add_ln703_361_fu_2153_p2;
wire   [15:0] sub_ln703_295_fu_2041_p2;
wire   [15:0] sub_ln703_296_fu_2046_p2;
wire   [15:0] add_ln703_352_fu_2051_p2;
wire   [15:0] sub_ln703_297_fu_2055_p2;
wire   [15:0] sub_ln703_298_fu_2065_p2;
wire   [15:0] sub_ln703_301_fu_2085_p2;
wire   [15:0] sub_ln703_303_fu_2094_p2;
wire   [15:0] sub_ln703_305_fu_2104_p2;
wire   [15:0] sub_ln703_306_fu_2109_p2;
wire   [15:0] add_ln703_355_fu_2114_p2;
wire   [15:0] sub_ln703_307_fu_2133_p2;
wire   [15:0] add_ln703_360_fu_2138_p2;
wire   [15:0] sub_ln703_308_fu_2143_p2;
wire   [15:0] sub_ln703_293_fu_2036_p2;
wire   [15:0] add_ln703_362_fu_2158_p2;
wire   [15:0] add_ln703_363_fu_2163_p2;
wire   [15:0] sub_ln703_310_fu_2168_p2;
wire   [15:0] add_ln703_364_fu_2178_p2;
wire   [15:0] add_ln703_365_fu_2183_p2;
wire   [15:0] add_ln703_366_fu_2193_p2;
wire   [15:0] sub_ln703_284_fu_1980_p2;
wire   [15:0] add_ln703_374_fu_2263_p2;
wire   [15:0] add_ln703_367_fu_2198_p2;
wire   [15:0] sub_ln703_287_fu_1998_p2;
wire   [15:0] add_ln703_376_fu_2278_p2;
wire   [15:0] add_ln703_378_fu_2288_p2;
wire   [15:0] sub_ln703_319_fu_2208_p2;
wire   [15:0] add_ln703_369_fu_2213_p2;
wire   [15:0] sub_ln703_322_fu_2223_p2;
wire   [15:0] add_ln703_375_fu_2268_p2;
wire   [15:0] sub_ln703_285_fu_1984_p2;
wire   [15:0] add_ln703_389_fu_2322_p2;
wire   [15:0] add_ln703_388_fu_2317_p2;
wire   [15:0] add_ln703_380_fu_2297_p2;
wire   [15:0] sub_ln703_267_fu_1872_p2;
wire   [15:0] add_ln703_399_fu_2342_p2;
wire   [15:0] add_ln703_398_fu_2337_p2;
wire   [15:0] sub_ln703_299_fu_2070_p2;
wire   [15:0] add_ln703_412_fu_2357_p2;
wire   [15:0] add_ln703_411_fu_2352_p2;
wire   [15:0] sub_ln703_315_fu_2188_p2;
wire   [15:0] add_ln703_414_fu_2367_p2;
wire   [15:0] sub_ln703_244_fu_1827_p2;
wire   [15:0] add_ln703_426_fu_2378_p2;
wire   [15:0] sub_ln703_313_fu_2413_p2;
wire   [15:0] sub_ln703_314_fu_2417_p2;
wire   [15:0] sub_ln703_316_fu_2421_p2;
wire   [15:0] add_ln703_368_fu_2429_p2;
wire   [15:0] add_ln703_370_fu_2437_p2;
wire   [15:0] sub_ln703_326_fu_2441_p2;
wire   [15:0] sub_ln703_312_fu_2409_p2;
wire   [15:0] add_ln703_373_fu_2445_p2;
wire   [15:0] sub_ln703_329_fu_2450_p2;
wire   [15:0] sub_ln703_317_fu_2425_p2;
wire   [15:0] sub_ln703_334_fu_2464_p2;
wire   [15:0] sub_ln703_336_fu_2469_p2;
wire   [15:0] sub_ln703_337_fu_2473_p2;
wire   [15:0] sub_ln703_338_fu_2478_p2;
wire   [15:0] sub_ln703_294_fu_2405_p2;
wire   [15:0] add_ln703_395_fu_2564_p2;
wire   [15:0] add_ln703_393_fu_2559_p2;
wire   [15:0] sub_ln703_339_fu_2482_p2;
wire   [15:0] add_ln703_382_fu_2486_p2;
wire   [15:0] add_ln703_383_fu_2490_p2;
wire   [15:0] sub_ln703_340_fu_2495_p2;
wire   [15:0] add_ln703_385_fu_2499_p2;
wire   [15:0] sub_ln703_341_fu_2504_p2;
wire   [15:0] sub_ln703_342_fu_2509_p2;
wire   [15:0] add_ln703_386_fu_2514_p2;
wire   [15:0] add_ln703_387_fu_2518_p2;
wire   [15:0] sub_ln703_344_fu_2523_p2;
wire   [15:0] add_ln703_391_fu_2527_p2;
wire   [15:0] sub_ln703_320_fu_2433_p2;
wire   [15:0] add_ln703_403_fu_2645_p2;
wire   [15:0] sub_ln703_347_fu_2536_p2;
wire   [15:0] add_ln703_392_fu_2540_p2;
wire   [15:0] sub_ln703_348_fu_2545_p2;
wire   [15:0] sub_ln703_350_fu_2554_p2;
wire   [15:0] add_ln703_407_fu_2675_p2;
wire   [15:0] add_ln703_396_fu_2568_p2;
wire   [15:0] sub_ln703_351_fu_2574_p2;
wire   [15:0] sub_ln703_352_fu_2579_p2;
wire   [15:0] sub_ln703_353_fu_2584_p2;
wire   [15:0] sub_ln703_354_fu_2589_p2;
wire   [15:0] sub_ln703_355_fu_2594_p2;
wire   [15:0] add_ln703_397_fu_2599_p2;
wire   [15:0] sub_ln703_358_fu_2613_p2;
wire   [15:0] sub_ln703_359_fu_2618_p2;
wire   [15:0] add_ln703_417_fu_2737_p2;
wire   [15:0] add_ln703_416_fu_2733_p2;
wire   [15:0] add_ln703_401_fu_2623_p2;
wire   [15:0] sub_ln703_360_fu_2627_p2;
wire   [15:0] add_ln703_419_fu_2757_p2;
wire   [15:0] sub_ln703_333_fu_2460_p2;
wire   [15:0] add_ln703_421_fu_2766_p2;
wire   [15:0] sub_ln703_362_fu_2641_p2;
wire   [15:0] add_ln703_405_fu_2650_p2;
wire   [15:0] add_ln703_406_fu_2655_p2;
wire   [15:0] sub_ln703_363_fu_2660_p2;
wire   [15:0] sub_ln703_364_fu_2665_p2;
wire   [15:0] add_ln703_408_fu_2679_p2;
wire   [15:0] sub_ln703_367_fu_2689_p2;
wire   [15:0] sub_ln703_368_fu_2694_p2;
wire   [15:0] add_ln703_409_fu_2704_p2;
wire   [15:0] add_ln703_429_fu_2825_p2;
wire   [15:0] add_ln703_430_fu_2829_p2;
wire   [15:0] sub_ln703_371_fu_2719_p2;
wire   [15:0] sub_ln703_373_fu_2723_p2;
wire   [15:0] sub_ln703_376_fu_2752_p2;
wire   [15:0] add_ln703_420_fu_2761_p2;
wire   [15:0] add_ln703_422_fu_2771_p2;
wire   [15:0] sub_ln703_378_fu_2776_p2;
wire   [15:0] sub_ln703_380_fu_2786_p2;
wire   [15:0] sub_ln703_382_fu_2796_p2;
wire   [15:0] sub_ln703_365_fu_2670_p2;
wire   [15:0] sub_ln703_370_fu_2714_p2;
wire   [15:0] sub_ln703_388_fu_2821_p2;
wire   [15:0] add_ln703_431_fu_2834_p2;
wire   [15:0] sub_ln703_391_fu_2844_p2;
wire   [15:0] sub_ln703_330_fu_2455_p2;
wire   [15:0] add_ln703_441_fu_2913_p2;
wire   [15:0] add_ln703_440_fu_2908_p2;
wire   [15:0] sub_ln703_396_fu_2858_p2;
wire   [15:0] sub_ln703_400_fu_2868_p2;
wire   [15:0] sub_ln703_383_fu_2801_p2;
wire   [15:0] add_ln703_438_fu_2888_p2;
wire   [15:0] sub_ln703_345_fu_2532_p2;
wire   [15:0] add_ln703_477_fu_2947_p2;
wire   [15:0] add_ln703_479_fu_2957_p2;
wire   [15:0] add_ln703_478_fu_2952_p2;
wire   [15:0] sub_ln703_395_fu_2853_p2;
wire   [15:0] sub_ln703_349_fu_2549_p2;
wire   [15:0] sub_ln703_372_fu_2985_p2;
wire   [15:0] sub_ln703_377_fu_2989_p2;
wire   [15:0] add_ln703_423_fu_2993_p2;
wire   [15:0] sub_ln703_384_fu_2997_p2;
wire   [15:0] add_ln703_425_fu_3001_p2;
wire   [15:0] sub_ln703_387_fu_3005_p2;
wire   [15:0] sub_ln703_390_fu_3009_p2;
wire   [15:0] add_ln703_432_fu_3014_p2;
wire   [15:0] sub_ln703_393_fu_3018_p2;
wire   [15:0] sub_ln703_394_fu_3022_p2;
wire   [15:0] sub_ln703_399_fu_3031_p2;
wire   [15:0] add_ln703_433_fu_3036_p2;
wire   [15:0] sub_ln703_401_fu_3040_p2;
wire   [15:0] sub_ln703_403_fu_3044_p2;
wire   [15:0] sub_ln703_404_fu_3049_p2;
wire   [15:0] add_ln703_437_fu_3053_p2;
wire   [15:0] sub_ln703_406_fu_3062_p2;
wire   [15:0] sub_ln703_410_fu_3071_p2;
wire   [15:0] add_ln703_439_fu_3075_p2;
wire   [15:0] add_ln703_450_fu_3168_p2;
wire   [15:0] sub_ln703_412_fu_3080_p2;
wire   [15:0] add_ln703_443_fu_3099_p2;
wire   [15:0] sub_ln703_417_fu_3103_p2;
wire   [15:0] sub_ln703_418_fu_3108_p2;
wire   [15:0] sub_ln703_419_fu_3113_p2;
wire   [15:0] sub_ln703_420_fu_3117_p2;
wire   [15:0] add_ln703_445_fu_3122_p2;
wire   [15:0] sub_ln703_424_fu_3140_p2;
wire   [15:0] add_ln703_455_fu_3237_p2;
wire   [15:0] sub_ln703_405_fu_3057_p2;
wire   [15:0] sub_ln703_425_fu_3145_p2;
wire   [15:0] add_ln703_448_fu_3150_p2;
wire   [15:0] sub_ln703_427_fu_3154_p2;
wire   [15:0] add_ln703_449_fu_3158_p2;
wire   [15:0] add_ln703_452_fu_3172_p2;
wire   [15:0] sub_ln703_429_fu_3177_p2;
wire   [15:0] sub_ln703_431_fu_3185_p2;
wire   [15:0] sub_ln703_413_fu_3084_p2;
wire   [15:0] sub_ln703_415_fu_3094_p2;
wire   [15:0] sub_ln703_432_fu_3190_p2;
wire   [15:0] sub_ln703_433_fu_3194_p2;
wire   [15:0] sub_ln703_436_fu_3208_p2;
wire   [15:0] sub_ln703_437_fu_3213_p2;
wire   [15:0] add_ln703_453_fu_3218_p2;
wire   [15:0] sub_ln703_438_fu_3223_p2;
wire   [15:0] sub_ln703_421_fu_3126_p2;
wire   [15:0] sub_ln703_439_fu_3228_p2;
wire   [15:0] sub_ln703_422_fu_3130_p2;
wire   [15:0] add_ln703_454_fu_3232_p2;
wire   [15:0] add_ln703_456_fu_3241_p2;
wire   [15:0] sub_ln703_440_fu_3247_p2;
wire   [15:0] sub_ln703_407_fu_3066_p2;
wire   [15:0] add_ln703_466_fu_3358_p2;
wire   [15:0] sub_ln703_441_fu_3252_p2;
wire   [15:0] sub_ln703_444_fu_3266_p2;
wire   [15:0] sub_ln703_445_fu_3271_p2;
wire   [15:0] sub_ln703_446_fu_3276_p2;
wire   [15:0] add_ln703_457_fu_3281_p2;
wire   [15:0] add_ln703_458_fu_3286_p2;
wire   [15:0] sub_ln703_414_fu_3089_p2;
wire   [15:0] add_ln703_470_fu_3398_p2;
wire   [15:0] add_ln703_459_fu_3292_p2;
wire   [15:0] sub_ln703_447_fu_3298_p2;
wire   [15:0] add_ln703_460_fu_3303_p2;
wire   [15:0] sub_ln703_398_fu_3026_p2;
wire   [15:0] add_ln703_474_fu_3428_p2;
wire   [15:0] add_ln703_473_fu_3423_p2;
wire   [15:0] add_ln703_461_fu_3323_p2;
wire   [15:0] sub_ln703_423_fu_3135_p2;
wire   [15:0] add_ln703_481_fu_3443_p2;
wire   [15:0] sub_ln703_442_fu_3256_p2;
wire   [15:0] sub_ln703_443_fu_3261_p2;
wire   [15:0] add_ln703_469_fu_3383_p2;
wire   [15:0] sub_ln703_430_fu_3181_p2;
wire   [15:0] add_ln703_489_fu_3468_p2;
wire   [15:0] add_ln703_472_fu_3413_p2;
wire   [15:0] sub_ln703_435_fu_3204_p2;
wire   [15:0] add_ln703_494_fu_3487_p2;
wire   [15:0] sub_ln703_449_fu_3313_p2;
wire   [15:0] add_ln703_486_fu_3453_p2;
wire   [15:0] add_ln703_487_fu_3458_p2;
wire   [15:0] add_ln703_490_fu_3473_p2;
wire   [15:0] add_ln703_495_fu_3492_p2;
wire   [15:0] add_ln703_476_fu_3531_p2;
wire   [15:0] sub_ln703_460_fu_3535_p2;
wire   [15:0] sub_ln703_462_fu_3539_p2;
wire   [15:0] sub_ln703_463_fu_3543_p2;
wire   [15:0] sub_ln703_464_fu_3547_p2;
wire   [15:0] sub_ln703_465_fu_3551_p2;
wire   [15:0] add_ln703_484_fu_3555_p2;
wire   [15:0] add_ln703_485_fu_3559_p2;
wire   [15:0] sub_ln703_466_fu_3563_p2;
wire   [15:0] sub_ln703_467_fu_3567_p2;
wire   [15:0] add_ln703_488_fu_3571_p2;
wire   [15:0] sub_ln703_468_fu_3575_p2;
wire   [15:0] sub_ln703_470_fu_3579_p2;
wire   [15:0] sub_ln703_471_fu_3583_p2;
wire   [15:0] sub_ln703_472_fu_3587_p2;
wire   [15:0] sub_ln703_473_fu_3591_p2;
wire   [15:0] add_ln703_493_fu_3595_p2;
wire   [15:0] sub_ln703_475_fu_3599_p2;
wire   [15:0] sub_ln703_476_fu_3603_p2;
wire   [15:0] sub_ln703_477_fu_3607_p2;
wire   [15:0] sub_ln703_478_fu_3612_p2;
wire   [15:0] add_ln703_498_fu_3616_p2;
wire   [15:0] sub_ln703_479_fu_3621_p2;
wire   [15:0] sub_ln703_480_fu_3626_p2;
wire   [15:0] add_ln703_499_fu_3631_p2;
wire   [15:0] sub_ln703_482_fu_3640_p2;
wire   [15:0] sub_ln703_483_fu_3645_p2;
wire   [15:0] sub_ln703_484_fu_3650_p2;
wire   [15:0] add_ln703_500_fu_3655_p2;
wire   [15:0] sub_ln703_485_fu_3660_p2;
wire   [15:0] sub_ln703_488_fu_3665_p2;
wire   [15:0] sub_ln703_489_fu_3670_p2;
wire   [15:0] sub_ln703_492_fu_3679_p2;
wire   [15:0] sub_ln703_493_fu_3684_p2;
wire   [15:0] sub_ln703_494_fu_3689_p2;
wire   [15:0] sub_ln703_495_fu_3694_p2;
wire   [15:0] sub_ln703_496_fu_3699_p2;
wire   [15:0] add_ln703_501_fu_3708_p2;
wire   [15:0] add_ln703_502_fu_3713_p2;
wire   [15:0] sub_ln703_499_fu_3723_p2;
wire   [15:0] add_ln703_508_fu_3843_p2;
wire   [15:0] sub_ln703_501_fu_3728_p2;
wire   [15:0] sub_ln703_502_fu_3732_p2;
wire   [15:0] add_ln703_514_fu_3862_p2;
wire   [15:0] add_ln703_518_fu_3875_p2;
wire   [15:0] add_ln703_517_fu_3871_p2;
wire   [15:0] sub_ln703_503_fu_3737_p2;
wire   [15:0] sub_ln703_504_fu_3742_p2;
wire   [15:0] sub_ln703_505_fu_3747_p2;
wire   [15:0] sub_ln703_481_fu_3636_p2;
wire   [15:0] sub_ln703_506_fu_3752_p2;
wire   [15:0] add_ln703_503_fu_3757_p2;
wire   [15:0] sub_ln703_507_fu_3762_p2;
wire   [15:0] sub_ln703_508_fu_3767_p2;
wire   [15:0] sub_ln703_509_fu_3772_p2;
wire   [15:0] add_ln703_504_fu_3777_p2;
wire   [15:0] sub_ln703_510_fu_3781_p2;
wire   [15:0] add_ln703_505_fu_3785_p2;
wire   [15:0] add_ln703_527_fu_3949_p2;
wire   [15:0] add_ln703_526_fu_3945_p2;
wire   [15:0] sub_ln703_511_fu_3790_p2;
wire   [15:0] sub_ln703_490_fu_3675_p2;
wire   [15:0] add_ln703_506_fu_3795_p2;
wire   [15:0] add_ln703_507_fu_3799_p2;
wire   [15:0] sub_ln703_512_fu_3804_p2;
wire   [15:0] sub_ln703_513_fu_3809_p2;
wire   [15:0] sub_ln703_514_fu_3814_p2;
wire   [15:0] sub_ln703_515_fu_3819_p2;
wire   [15:0] sub_ln703_497_fu_3704_p2;
wire   [15:0] sub_ln703_516_fu_3824_p2;
wire   [15:0] sub_ln703_517_fu_3829_p2;
wire   [15:0] sub_ln703_498_fu_3718_p2;
wire   [15:0] sub_ln703_518_fu_3834_p2;
wire   [15:0] sub_ln703_519_fu_3839_p2;
wire   [15:0] add_ln703_511_fu_3847_p2;
wire   [15:0] acc_1_V_fu_3852_p2;
wire   [15:0] acc_2_V_fu_3857_p2;
wire   [15:0] acc_3_V_fu_3866_p2;
wire   [15:0] acc_4_V_fu_3879_p2;
wire   [15:0] acc_5_V_fu_3885_p2;
wire   [15:0] acc_6_V_fu_3890_p2;
wire   [15:0] acc_7_V_fu_3895_p2;
wire   [15:0] acc_8_V_fu_3900_p2;
wire   [15:0] acc_9_V_fu_3905_p2;
wire   [15:0] acc_10_V_fu_3910_p2;
wire   [15:0] acc_11_V_fu_3915_p2;
wire   [15:0] acc_12_V_fu_3920_p2;
wire   [15:0] acc_13_V_fu_3925_p2;
wire   [15:0] acc_14_V_fu_3930_p2;
wire   [15:0] acc_15_V_fu_3935_p2;
wire   [15:0] acc_16_V_fu_3940_p2;
wire   [15:0] acc_17_V_fu_3953_p2;
wire   [15:0] acc_18_V_fu_3959_p2;
wire   [15:0] acc_19_V_fu_3964_p2;
wire   [15:0] acc_20_V_fu_3969_p2;
wire   [15:0] acc_21_V_fu_3974_p2;
wire   [15:0] acc_22_V_fu_3979_p2;
wire   [15:0] acc_23_V_fu_3984_p2;
wire   [15:0] acc_24_V_fu_3989_p2;
wire   [15:0] acc_25_V_fu_3994_p2;
wire   [15:0] acc_26_V_fu_3999_p2;
wire   [15:0] acc_27_V_fu_4004_p2;
wire   [15:0] acc_28_V_fu_4009_p2;
wire   [15:0] acc_29_V_fu_4014_p2;
wire   [15:0] acc_30_V_fu_4019_p2;
wire   [15:0] acc_31_V_fu_4024_p2;
reg    ap_ce_reg;
reg   [15:0] data_0_V_read_int_reg;
reg   [15:0] data_1_V_read_int_reg;
reg   [15:0] data_2_V_read_int_reg;
reg   [15:0] data_3_V_read_int_reg;
reg   [15:0] data_4_V_read_int_reg;
reg   [15:0] data_5_V_read_int_reg;
reg   [15:0] data_6_V_read_int_reg;
reg   [15:0] data_7_V_read_int_reg;
reg   [15:0] data_8_V_read_int_reg;
reg   [15:0] data_9_V_read_int_reg;
reg   [15:0] data_10_V_read_int_reg;
reg   [15:0] data_11_V_read_int_reg;
reg   [15:0] data_12_V_read_int_reg;
reg   [15:0] data_13_V_read_int_reg;
reg   [15:0] data_14_V_read_int_reg;
reg   [15:0] data_15_V_read_int_reg;
reg   [15:0] data_16_V_read_int_reg;
reg   [15:0] data_17_V_read_int_reg;
reg   [15:0] data_18_V_read_int_reg;
reg   [15:0] data_19_V_read_int_reg;
reg   [15:0] data_20_V_read_int_reg;
reg   [15:0] data_21_V_read_int_reg;
reg   [15:0] data_22_V_read_int_reg;
reg   [15:0] data_23_V_read_int_reg;
reg   [15:0] data_24_V_read_int_reg;
reg   [15:0] data_25_V_read_int_reg;
reg   [15:0] data_26_V_read_int_reg;
reg   [15:0] data_27_V_read_int_reg;
reg   [15:0] data_28_V_read_int_reg;
reg   [15:0] data_29_V_read_int_reg;
reg   [15:0] data_30_V_read_int_reg;
reg   [15:0] data_31_V_read_int_reg;
reg   [15:0] ap_return_0_int_reg;
reg   [15:0] ap_return_1_int_reg;
reg   [15:0] ap_return_2_int_reg;
reg   [15:0] ap_return_3_int_reg;
reg   [15:0] ap_return_4_int_reg;
reg   [15:0] ap_return_5_int_reg;
reg   [15:0] ap_return_6_int_reg;
reg   [15:0] ap_return_7_int_reg;
reg   [15:0] ap_return_8_int_reg;
reg   [15:0] ap_return_9_int_reg;
reg   [15:0] ap_return_10_int_reg;
reg   [15:0] ap_return_11_int_reg;
reg   [15:0] ap_return_12_int_reg;
reg   [15:0] ap_return_13_int_reg;
reg   [15:0] ap_return_14_int_reg;
reg   [15:0] ap_return_15_int_reg;
reg   [15:0] ap_return_16_int_reg;
reg   [15:0] ap_return_17_int_reg;
reg   [15:0] ap_return_18_int_reg;
reg   [15:0] ap_return_19_int_reg;
reg   [15:0] ap_return_20_int_reg;
reg   [15:0] ap_return_21_int_reg;
reg   [15:0] ap_return_22_int_reg;
reg   [15:0] ap_return_23_int_reg;
reg   [15:0] ap_return_24_int_reg;
reg   [15:0] ap_return_25_int_reg;
reg   [15:0] ap_return_26_int_reg;
reg   [15:0] ap_return_27_int_reg;
reg   [15:0] ap_return_28_int_reg;
reg   [15:0] ap_return_29_int_reg;
reg   [15:0] ap_return_30_int_reg;
reg   [15:0] ap_return_31_int_reg;

always @ (posedge ap_clk) begin
    ap_ce_reg <= ap_ce;
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_ce_reg))) begin
        add_ln703_200_reg_5077 <= add_ln703_200_fu_304_p2;
        add_ln703_200_reg_5077_pp0_iter2_reg <= add_ln703_200_reg_5077;
        add_ln703_201_reg_5090 <= add_ln703_201_fu_312_p2;
        add_ln703_201_reg_5090_pp0_iter2_reg <= add_ln703_201_reg_5090;
        add_ln703_202_reg_5096 <= add_ln703_202_fu_316_p2;
        add_ln703_202_reg_5096_pp0_iter2_reg <= add_ln703_202_reg_5096;
        add_ln703_203_reg_5113 <= add_ln703_203_fu_329_p2;
        add_ln703_204_reg_5101 <= add_ln703_204_fu_320_p2;
        add_ln703_204_reg_5101_pp0_iter2_reg <= add_ln703_204_reg_5101;
        add_ln703_205_reg_5119 <= add_ln703_205_fu_333_p2;
        add_ln703_206_reg_5131 <= add_ln703_206_fu_341_p2;
        add_ln703_207_reg_5107 <= add_ln703_207_fu_325_p2;
        add_ln703_207_reg_5107_pp0_iter2_reg <= add_ln703_207_reg_5107;
        add_ln703_208_reg_5137 <= add_ln703_208_fu_345_p2;
        add_ln703_209_reg_5178 <= add_ln703_209_fu_416_p2;
        add_ln703_210_reg_5143 <= add_ln703_210_fu_349_p2;
        add_ln703_210_reg_5143_pp0_iter3_reg <= add_ln703_210_reg_5143;
        add_ln703_211_reg_5184 <= add_ln703_211_fu_420_p2;
        add_ln703_213_reg_5189 <= add_ln703_213_fu_429_p2;
        add_ln703_214_reg_5194 <= add_ln703_214_fu_433_p2;
        add_ln703_216_reg_5215 <= add_ln703_216_fu_461_p2;
        add_ln703_220_reg_5221 <= add_ln703_220_fu_484_p2;
        add_ln703_223_reg_5231 <= add_ln703_223_fu_507_p2;
        add_ln703_225_reg_5237 <= add_ln703_225_fu_513_p2;
        add_ln703_227_reg_5242 <= add_ln703_227_fu_522_p2;
        add_ln703_233_reg_5149 <= add_ln703_233_fu_353_p2;
        add_ln703_233_reg_5149_pp0_iter3_reg <= add_ln703_233_reg_5149;
        add_ln703_234_reg_5264 <= add_ln703_234_fu_564_p2;
        add_ln703_238_reg_5269 <= add_ln703_238_fu_569_p2;
        add_ln703_246_reg_5320 <= add_ln703_246_fu_787_p2;
        add_ln703_247_reg_5159 <= add_ln703_247_fu_357_p2;
        add_ln703_247_reg_5159_pp0_iter3_reg <= add_ln703_247_reg_5159;
        add_ln703_251_reg_5289 <= add_ln703_251_fu_589_p2;
        add_ln703_258_reg_5295 <= add_ln703_258_fu_593_p2;
        add_ln703_261_reg_5360 <= add_ln703_261_fu_955_p2;
        add_ln703_267_reg_5405 <= add_ln703_267_fu_1055_p2;
        add_ln703_268_reg_5415 <= add_ln703_268_fu_1065_p2;
        add_ln703_272_reg_5304 <= add_ln703_272_fu_597_p2;
        add_ln703_272_reg_5304_pp0_iter4_reg <= add_ln703_272_reg_5304;
        add_ln703_274_reg_5420 <= add_ln703_274_fu_1089_p2;
        add_ln703_276_reg_5430 <= add_ln703_276_fu_1100_p2;
        add_ln703_278_reg_5435 <= add_ln703_278_fu_1105_p2;
        add_ln703_281_reg_5455 <= add_ln703_281_fu_1129_p2;
        add_ln703_283_reg_5460 <= add_ln703_283_fu_1140_p2;
        add_ln703_287_reg_5525 <= add_ln703_287_fu_1354_p2;
        add_ln703_288_reg_5475 <= add_ln703_288_fu_1156_p2;
        add_ln703_291_reg_5530 <= add_ln703_291_fu_1371_p2;
        add_ln703_301_reg_5550 <= add_ln703_301_fu_1494_p2;
        add_ln703_304_reg_5314 <= add_ln703_304_fu_601_p2;
        add_ln703_307_reg_5555 <= add_ln703_307_fu_1504_p2;
        add_ln703_309_reg_5484 <= add_ln703_309_fu_1179_p2;
        add_ln703_314_reg_5490 <= add_ln703_314_fu_1183_p2;
        add_ln703_316_reg_5496 <= add_ln703_316_fu_1187_p2;
        add_ln703_321_reg_5590 <= add_ln703_321_fu_1636_p2;
        add_ln703_323_reg_5506 <= add_ln703_323_fu_1198_p2;
        add_ln703_326_reg_5625 <= add_ln703_326_fu_1686_p2;
        add_ln703_330_reg_5640 <= add_ln703_330_fu_1710_p2;
        add_ln703_335_reg_5645 <= add_ln703_335_fu_1730_p2;
        add_ln703_339_reg_5655 <= add_ln703_339_fu_1740_p2;
        add_ln703_343_reg_5660 <= add_ln703_343_fu_1745_p2;
        add_ln703_347_reg_5675 <= add_ln703_347_fu_1760_p2;
        add_ln703_353_reg_5743 <= add_ln703_353_fu_2060_p2;
        add_ln703_354_reg_5753 <= add_ln703_354_fu_2080_p2;
        add_ln703_357_reg_5683 <= add_ln703_357_fu_1764_p2;
        add_ln703_357_reg_5683_pp0_iter6_reg <= add_ln703_357_reg_5683;
        add_ln703_359_reg_5768 <= add_ln703_359_fu_2127_p2;
        add_ln703_371_reg_5691 <= add_ln703_371_fu_1768_p2;
        add_ln703_372_reg_5793 <= add_ln703_372_fu_2228_p2;
        add_ln703_377_reg_5833 <= add_ln703_377_fu_2283_p2;
        add_ln703_379_reg_5838 <= add_ln703_379_fu_2292_p2;
        add_ln703_381_reg_5848 <= add_ln703_381_fu_2307_p2;
        add_ln703_384_reg_5701 <= add_ln703_384_fu_1772_p2;
        add_ln703_384_reg_5701_pp0_iter6_reg <= add_ln703_384_reg_5701;
        add_ln703_390_reg_5858 <= add_ln703_390_fu_2326_p2;
        add_ln703_394_reg_5710 <= add_ln703_394_fu_1776_p2;
        add_ln703_394_reg_5710_pp0_iter6_reg <= add_ln703_394_reg_5710;
        add_ln703_400_reg_5868 <= add_ln703_400_fu_2346_p2;
        add_ln703_402_reg_5931 <= add_ln703_402_fu_2631_p2;
        add_ln703_404_reg_5718 <= add_ln703_404_fu_1780_p2;
        add_ln703_404_reg_5718_pp0_iter6_reg <= add_ln703_404_reg_5718;
        add_ln703_410_reg_5951 <= add_ln703_410_fu_2709_p2;
        add_ln703_413_reg_5873 <= add_ln703_413_fu_2361_p2;
        add_ln703_415_reg_5878 <= add_ln703_415_fu_2372_p2;
        add_ln703_418_reg_5961 <= add_ln703_418_fu_2741_p2;
        add_ln703_424_reg_5981 <= add_ln703_424_fu_2806_p2;
        add_ln703_427_reg_5883 <= add_ln703_427_fu_2383_p2;
        add_ln703_428_reg_5888 <= add_ln703_428_fu_2389_p2;
        add_ln703_434_reg_6011 <= add_ln703_434_fu_2873_p2;
        add_ln703_435_reg_5894 <= add_ln703_435_fu_2393_p2;
        add_ln703_436_reg_6021 <= add_ln703_436_fu_2883_p2;
        add_ln703_442_reg_6041 <= add_ln703_442_fu_2917_p2;
        add_ln703_444_reg_6051 <= add_ln703_444_fu_2928_p2;
        add_ln703_446_reg_5901 <= add_ln703_446_fu_2397_p2;
        add_ln703_447_reg_6056 <= add_ln703_447_fu_2933_p2;
        add_ln703_451_reg_6066 <= add_ln703_451_fu_2943_p2;
        add_ln703_451_reg_6066_pp0_iter8_reg <= add_ln703_451_reg_6066;
        add_ln703_462_reg_5909 <= add_ln703_462_fu_2401_p2;
        add_ln703_462_reg_5909_pp0_iter7_reg <= add_ln703_462_reg_5909;
        add_ln703_462_reg_5909_pp0_iter8_reg <= add_ln703_462_reg_5909_pp0_iter7_reg;
        add_ln703_463_reg_6128 <= add_ln703_463_fu_3328_p2;
        add_ln703_464_reg_6133 <= add_ln703_464_fu_3333_p2;
        add_ln703_465_reg_6138 <= add_ln703_465_fu_3338_p2;
        add_ln703_467_reg_6158 <= add_ln703_467_fu_3363_p2;
        add_ln703_468_reg_6173 <= add_ln703_468_fu_3378_p2;
        add_ln703_471_reg_6188 <= add_ln703_471_fu_3403_p2;
        add_ln703_475_reg_6203 <= add_ln703_475_fu_3432_p2;
        add_ln703_480_reg_6072 <= add_ln703_480_fu_2961_p2;
        add_ln703_480_reg_6072_pp0_iter8_reg <= add_ln703_480_reg_6072;
        add_ln703_482_reg_6077 <= add_ln703_482_fu_2967_p2;
        add_ln703_483_reg_6213 <= add_ln703_483_fu_3448_p2;
        add_ln703_491_reg_6087 <= add_ln703_491_fu_2971_p2;
        add_ln703_491_reg_6087_pp0_iter8_reg <= add_ln703_491_reg_6087;
        add_ln703_492_reg_6223 <= add_ln703_492_fu_3478_p2;
        add_ln703_496_reg_6234 <= add_ln703_496_fu_3497_p2;
        add_ln703_497_reg_6239 <= add_ln703_497_fu_3501_p2;
        add_ln703_509_reg_6092 <= add_ln703_509_fu_2976_p2;
        add_ln703_509_reg_6092_pp0_iter8_reg <= add_ln703_509_reg_6092;
        add_ln703_510_reg_6264 <= add_ln703_510_fu_3527_p2;
        add_ln703_516_reg_6103 <= add_ln703_516_fu_2980_p2;
        add_ln703_516_reg_6103_pp0_iter8_reg <= add_ln703_516_reg_6103;
        add_ln703_reg_5052 <= add_ln703_fu_280_p2;
        data_10_V_read11_reg_4832 <= data_10_V_read_int_reg;
        data_10_V_read11_reg_4832_pp0_iter1_reg <= data_10_V_read11_reg_4832;
        data_10_V_read11_reg_4832_pp0_iter2_reg <= data_10_V_read11_reg_4832_pp0_iter1_reg;
        data_10_V_read11_reg_4832_pp0_iter3_reg <= data_10_V_read11_reg_4832_pp0_iter2_reg;
        data_10_V_read11_reg_4832_pp0_iter4_reg <= data_10_V_read11_reg_4832_pp0_iter3_reg;
        data_11_V_read12_reg_4808 <= data_11_V_read_int_reg;
        data_11_V_read12_reg_4808_pp0_iter1_reg <= data_11_V_read12_reg_4808;
        data_11_V_read12_reg_4808_pp0_iter2_reg <= data_11_V_read12_reg_4808_pp0_iter1_reg;
        data_11_V_read12_reg_4808_pp0_iter3_reg <= data_11_V_read12_reg_4808_pp0_iter2_reg;
        data_11_V_read12_reg_4808_pp0_iter4_reg <= data_11_V_read12_reg_4808_pp0_iter3_reg;
        data_12_V_read13_reg_4778 <= data_12_V_read_int_reg;
        data_12_V_read13_reg_4778_pp0_iter1_reg <= data_12_V_read13_reg_4778;
        data_12_V_read13_reg_4778_pp0_iter2_reg <= data_12_V_read13_reg_4778_pp0_iter1_reg;
        data_12_V_read13_reg_4778_pp0_iter3_reg <= data_12_V_read13_reg_4778_pp0_iter2_reg;
        data_12_V_read13_reg_4778_pp0_iter4_reg <= data_12_V_read13_reg_4778_pp0_iter3_reg;
        data_13_V_read14_reg_4745 <= data_13_V_read_int_reg;
        data_13_V_read14_reg_4745_pp0_iter1_reg <= data_13_V_read14_reg_4745;
        data_13_V_read14_reg_4745_pp0_iter2_reg <= data_13_V_read14_reg_4745_pp0_iter1_reg;
        data_13_V_read14_reg_4745_pp0_iter3_reg <= data_13_V_read14_reg_4745_pp0_iter2_reg;
        data_13_V_read14_reg_4745_pp0_iter4_reg <= data_13_V_read14_reg_4745_pp0_iter3_reg;
        data_13_V_read14_reg_4745_pp0_iter5_reg <= data_13_V_read14_reg_4745_pp0_iter4_reg;
        data_14_V_read15_reg_4714 <= data_14_V_read_int_reg;
        data_14_V_read15_reg_4714_pp0_iter1_reg <= data_14_V_read15_reg_4714;
        data_14_V_read15_reg_4714_pp0_iter2_reg <= data_14_V_read15_reg_4714_pp0_iter1_reg;
        data_14_V_read15_reg_4714_pp0_iter3_reg <= data_14_V_read15_reg_4714_pp0_iter2_reg;
        data_14_V_read15_reg_4714_pp0_iter4_reg <= data_14_V_read15_reg_4714_pp0_iter3_reg;
        data_14_V_read15_reg_4714_pp0_iter5_reg <= data_14_V_read15_reg_4714_pp0_iter4_reg;
        data_15_V_read16_reg_4682 <= data_15_V_read_int_reg;
        data_15_V_read16_reg_4682_pp0_iter1_reg <= data_15_V_read16_reg_4682;
        data_15_V_read16_reg_4682_pp0_iter2_reg <= data_15_V_read16_reg_4682_pp0_iter1_reg;
        data_15_V_read16_reg_4682_pp0_iter3_reg <= data_15_V_read16_reg_4682_pp0_iter2_reg;
        data_15_V_read16_reg_4682_pp0_iter4_reg <= data_15_V_read16_reg_4682_pp0_iter3_reg;
        data_15_V_read16_reg_4682_pp0_iter5_reg <= data_15_V_read16_reg_4682_pp0_iter4_reg;
        data_16_V_read17_reg_4650 <= data_16_V_read_int_reg;
        data_16_V_read17_reg_4650_pp0_iter1_reg <= data_16_V_read17_reg_4650;
        data_16_V_read17_reg_4650_pp0_iter2_reg <= data_16_V_read17_reg_4650_pp0_iter1_reg;
        data_16_V_read17_reg_4650_pp0_iter3_reg <= data_16_V_read17_reg_4650_pp0_iter2_reg;
        data_16_V_read17_reg_4650_pp0_iter4_reg <= data_16_V_read17_reg_4650_pp0_iter3_reg;
        data_16_V_read17_reg_4650_pp0_iter5_reg <= data_16_V_read17_reg_4650_pp0_iter4_reg;
        data_17_V_read_8_reg_4621 <= data_17_V_read_int_reg;
        data_17_V_read_8_reg_4621_pp0_iter1_reg <= data_17_V_read_8_reg_4621;
        data_17_V_read_8_reg_4621_pp0_iter2_reg <= data_17_V_read_8_reg_4621_pp0_iter1_reg;
        data_17_V_read_8_reg_4621_pp0_iter3_reg <= data_17_V_read_8_reg_4621_pp0_iter2_reg;
        data_17_V_read_8_reg_4621_pp0_iter4_reg <= data_17_V_read_8_reg_4621_pp0_iter3_reg;
        data_17_V_read_8_reg_4621_pp0_iter5_reg <= data_17_V_read_8_reg_4621_pp0_iter4_reg;
        data_17_V_read_8_reg_4621_pp0_iter6_reg <= data_17_V_read_8_reg_4621_pp0_iter5_reg;
        data_18_V_read_7_reg_4594 <= data_18_V_read_int_reg;
        data_18_V_read_7_reg_4594_pp0_iter1_reg <= data_18_V_read_7_reg_4594;
        data_18_V_read_7_reg_4594_pp0_iter2_reg <= data_18_V_read_7_reg_4594_pp0_iter1_reg;
        data_18_V_read_7_reg_4594_pp0_iter3_reg <= data_18_V_read_7_reg_4594_pp0_iter2_reg;
        data_18_V_read_7_reg_4594_pp0_iter4_reg <= data_18_V_read_7_reg_4594_pp0_iter3_reg;
        data_18_V_read_7_reg_4594_pp0_iter5_reg <= data_18_V_read_7_reg_4594_pp0_iter4_reg;
        data_18_V_read_7_reg_4594_pp0_iter6_reg <= data_18_V_read_7_reg_4594_pp0_iter5_reg;
        data_19_V_read_7_reg_4567 <= data_19_V_read_int_reg;
        data_19_V_read_7_reg_4567_pp0_iter1_reg <= data_19_V_read_7_reg_4567;
        data_19_V_read_7_reg_4567_pp0_iter2_reg <= data_19_V_read_7_reg_4567_pp0_iter1_reg;
        data_19_V_read_7_reg_4567_pp0_iter3_reg <= data_19_V_read_7_reg_4567_pp0_iter2_reg;
        data_19_V_read_7_reg_4567_pp0_iter4_reg <= data_19_V_read_7_reg_4567_pp0_iter3_reg;
        data_19_V_read_7_reg_4567_pp0_iter5_reg <= data_19_V_read_7_reg_4567_pp0_iter4_reg;
        data_19_V_read_7_reg_4567_pp0_iter6_reg <= data_19_V_read_7_reg_4567_pp0_iter5_reg;
        data_20_V_read21_reg_4539 <= data_20_V_read_int_reg;
        data_20_V_read21_reg_4539_pp0_iter1_reg <= data_20_V_read21_reg_4539;
        data_20_V_read21_reg_4539_pp0_iter2_reg <= data_20_V_read21_reg_4539_pp0_iter1_reg;
        data_20_V_read21_reg_4539_pp0_iter3_reg <= data_20_V_read21_reg_4539_pp0_iter2_reg;
        data_20_V_read21_reg_4539_pp0_iter4_reg <= data_20_V_read21_reg_4539_pp0_iter3_reg;
        data_20_V_read21_reg_4539_pp0_iter5_reg <= data_20_V_read21_reg_4539_pp0_iter4_reg;
        data_20_V_read21_reg_4539_pp0_iter6_reg <= data_20_V_read21_reg_4539_pp0_iter5_reg;
        data_21_V_read22_reg_4512 <= data_21_V_read_int_reg;
        data_21_V_read22_reg_4512_pp0_iter1_reg <= data_21_V_read22_reg_4512;
        data_21_V_read22_reg_4512_pp0_iter2_reg <= data_21_V_read22_reg_4512_pp0_iter1_reg;
        data_21_V_read22_reg_4512_pp0_iter3_reg <= data_21_V_read22_reg_4512_pp0_iter2_reg;
        data_21_V_read22_reg_4512_pp0_iter4_reg <= data_21_V_read22_reg_4512_pp0_iter3_reg;
        data_21_V_read22_reg_4512_pp0_iter5_reg <= data_21_V_read22_reg_4512_pp0_iter4_reg;
        data_21_V_read22_reg_4512_pp0_iter6_reg <= data_21_V_read22_reg_4512_pp0_iter5_reg;
        data_22_V_read23_reg_4483 <= data_22_V_read_int_reg;
        data_22_V_read23_reg_4483_pp0_iter1_reg <= data_22_V_read23_reg_4483;
        data_22_V_read23_reg_4483_pp0_iter2_reg <= data_22_V_read23_reg_4483_pp0_iter1_reg;
        data_22_V_read23_reg_4483_pp0_iter3_reg <= data_22_V_read23_reg_4483_pp0_iter2_reg;
        data_22_V_read23_reg_4483_pp0_iter4_reg <= data_22_V_read23_reg_4483_pp0_iter3_reg;
        data_22_V_read23_reg_4483_pp0_iter5_reg <= data_22_V_read23_reg_4483_pp0_iter4_reg;
        data_22_V_read23_reg_4483_pp0_iter6_reg <= data_22_V_read23_reg_4483_pp0_iter5_reg;
        data_22_V_read23_reg_4483_pp0_iter7_reg <= data_22_V_read23_reg_4483_pp0_iter6_reg;
        data_23_V_read24_reg_4451 <= data_23_V_read_int_reg;
        data_23_V_read24_reg_4451_pp0_iter1_reg <= data_23_V_read24_reg_4451;
        data_23_V_read24_reg_4451_pp0_iter2_reg <= data_23_V_read24_reg_4451_pp0_iter1_reg;
        data_23_V_read24_reg_4451_pp0_iter3_reg <= data_23_V_read24_reg_4451_pp0_iter2_reg;
        data_23_V_read24_reg_4451_pp0_iter4_reg <= data_23_V_read24_reg_4451_pp0_iter3_reg;
        data_23_V_read24_reg_4451_pp0_iter5_reg <= data_23_V_read24_reg_4451_pp0_iter4_reg;
        data_23_V_read24_reg_4451_pp0_iter6_reg <= data_23_V_read24_reg_4451_pp0_iter5_reg;
        data_23_V_read24_reg_4451_pp0_iter7_reg <= data_23_V_read24_reg_4451_pp0_iter6_reg;
        data_24_V_read25_reg_4421 <= data_24_V_read_int_reg;
        data_24_V_read25_reg_4421_pp0_iter1_reg <= data_24_V_read25_reg_4421;
        data_24_V_read25_reg_4421_pp0_iter2_reg <= data_24_V_read25_reg_4421_pp0_iter1_reg;
        data_24_V_read25_reg_4421_pp0_iter3_reg <= data_24_V_read25_reg_4421_pp0_iter2_reg;
        data_24_V_read25_reg_4421_pp0_iter4_reg <= data_24_V_read25_reg_4421_pp0_iter3_reg;
        data_24_V_read25_reg_4421_pp0_iter5_reg <= data_24_V_read25_reg_4421_pp0_iter4_reg;
        data_24_V_read25_reg_4421_pp0_iter6_reg <= data_24_V_read25_reg_4421_pp0_iter5_reg;
        data_24_V_read25_reg_4421_pp0_iter7_reg <= data_24_V_read25_reg_4421_pp0_iter6_reg;
        data_25_V_read26_reg_4391 <= data_25_V_read_int_reg;
        data_25_V_read26_reg_4391_pp0_iter1_reg <= data_25_V_read26_reg_4391;
        data_25_V_read26_reg_4391_pp0_iter2_reg <= data_25_V_read26_reg_4391_pp0_iter1_reg;
        data_25_V_read26_reg_4391_pp0_iter3_reg <= data_25_V_read26_reg_4391_pp0_iter2_reg;
        data_25_V_read26_reg_4391_pp0_iter4_reg <= data_25_V_read26_reg_4391_pp0_iter3_reg;
        data_25_V_read26_reg_4391_pp0_iter5_reg <= data_25_V_read26_reg_4391_pp0_iter4_reg;
        data_25_V_read26_reg_4391_pp0_iter6_reg <= data_25_V_read26_reg_4391_pp0_iter5_reg;
        data_25_V_read26_reg_4391_pp0_iter7_reg <= data_25_V_read26_reg_4391_pp0_iter6_reg;
        data_26_V_read27_reg_4365 <= data_26_V_read_int_reg;
        data_26_V_read27_reg_4365_pp0_iter1_reg <= data_26_V_read27_reg_4365;
        data_26_V_read27_reg_4365_pp0_iter2_reg <= data_26_V_read27_reg_4365_pp0_iter1_reg;
        data_26_V_read27_reg_4365_pp0_iter3_reg <= data_26_V_read27_reg_4365_pp0_iter2_reg;
        data_26_V_read27_reg_4365_pp0_iter4_reg <= data_26_V_read27_reg_4365_pp0_iter3_reg;
        data_26_V_read27_reg_4365_pp0_iter5_reg <= data_26_V_read27_reg_4365_pp0_iter4_reg;
        data_26_V_read27_reg_4365_pp0_iter6_reg <= data_26_V_read27_reg_4365_pp0_iter5_reg;
        data_26_V_read27_reg_4365_pp0_iter7_reg <= data_26_V_read27_reg_4365_pp0_iter6_reg;
        data_27_V_read_8_reg_4342 <= data_27_V_read_int_reg;
        data_27_V_read_8_reg_4342_pp0_iter1_reg <= data_27_V_read_8_reg_4342;
        data_27_V_read_8_reg_4342_pp0_iter2_reg <= data_27_V_read_8_reg_4342_pp0_iter1_reg;
        data_27_V_read_8_reg_4342_pp0_iter3_reg <= data_27_V_read_8_reg_4342_pp0_iter2_reg;
        data_27_V_read_8_reg_4342_pp0_iter4_reg <= data_27_V_read_8_reg_4342_pp0_iter3_reg;
        data_27_V_read_8_reg_4342_pp0_iter5_reg <= data_27_V_read_8_reg_4342_pp0_iter4_reg;
        data_27_V_read_8_reg_4342_pp0_iter6_reg <= data_27_V_read_8_reg_4342_pp0_iter5_reg;
        data_27_V_read_8_reg_4342_pp0_iter7_reg <= data_27_V_read_8_reg_4342_pp0_iter6_reg;
        data_28_V_read_7_reg_4313 <= data_28_V_read_int_reg;
        data_28_V_read_7_reg_4313_pp0_iter1_reg <= data_28_V_read_7_reg_4313;
        data_28_V_read_7_reg_4313_pp0_iter2_reg <= data_28_V_read_7_reg_4313_pp0_iter1_reg;
        data_28_V_read_7_reg_4313_pp0_iter3_reg <= data_28_V_read_7_reg_4313_pp0_iter2_reg;
        data_28_V_read_7_reg_4313_pp0_iter4_reg <= data_28_V_read_7_reg_4313_pp0_iter3_reg;
        data_28_V_read_7_reg_4313_pp0_iter5_reg <= data_28_V_read_7_reg_4313_pp0_iter4_reg;
        data_28_V_read_7_reg_4313_pp0_iter6_reg <= data_28_V_read_7_reg_4313_pp0_iter5_reg;
        data_28_V_read_7_reg_4313_pp0_iter7_reg <= data_28_V_read_7_reg_4313_pp0_iter6_reg;
        data_28_V_read_7_reg_4313_pp0_iter8_reg <= data_28_V_read_7_reg_4313_pp0_iter7_reg;
        data_29_V_read_7_reg_4279 <= data_29_V_read_int_reg;
        data_29_V_read_7_reg_4279_pp0_iter1_reg <= data_29_V_read_7_reg_4279;
        data_29_V_read_7_reg_4279_pp0_iter2_reg <= data_29_V_read_7_reg_4279_pp0_iter1_reg;
        data_29_V_read_7_reg_4279_pp0_iter3_reg <= data_29_V_read_7_reg_4279_pp0_iter2_reg;
        data_29_V_read_7_reg_4279_pp0_iter4_reg <= data_29_V_read_7_reg_4279_pp0_iter3_reg;
        data_29_V_read_7_reg_4279_pp0_iter5_reg <= data_29_V_read_7_reg_4279_pp0_iter4_reg;
        data_29_V_read_7_reg_4279_pp0_iter6_reg <= data_29_V_read_7_reg_4279_pp0_iter5_reg;
        data_29_V_read_7_reg_4279_pp0_iter7_reg <= data_29_V_read_7_reg_4279_pp0_iter6_reg;
        data_29_V_read_7_reg_4279_pp0_iter8_reg <= data_29_V_read_7_reg_4279_pp0_iter7_reg;
        data_2_V_read_9_reg_5035 <= data_2_V_read_int_reg;
        data_30_V_read31_reg_4250 <= data_30_V_read_int_reg;
        data_30_V_read31_reg_4250_pp0_iter1_reg <= data_30_V_read31_reg_4250;
        data_30_V_read31_reg_4250_pp0_iter2_reg <= data_30_V_read31_reg_4250_pp0_iter1_reg;
        data_30_V_read31_reg_4250_pp0_iter3_reg <= data_30_V_read31_reg_4250_pp0_iter2_reg;
        data_30_V_read31_reg_4250_pp0_iter4_reg <= data_30_V_read31_reg_4250_pp0_iter3_reg;
        data_30_V_read31_reg_4250_pp0_iter5_reg <= data_30_V_read31_reg_4250_pp0_iter4_reg;
        data_30_V_read31_reg_4250_pp0_iter6_reg <= data_30_V_read31_reg_4250_pp0_iter5_reg;
        data_30_V_read31_reg_4250_pp0_iter7_reg <= data_30_V_read31_reg_4250_pp0_iter6_reg;
        data_30_V_read31_reg_4250_pp0_iter8_reg <= data_30_V_read31_reg_4250_pp0_iter7_reg;
        data_31_V_read32_reg_4221 <= data_31_V_read_int_reg;
        data_31_V_read32_reg_4221_pp0_iter1_reg <= data_31_V_read32_reg_4221;
        data_31_V_read32_reg_4221_pp0_iter2_reg <= data_31_V_read32_reg_4221_pp0_iter1_reg;
        data_31_V_read32_reg_4221_pp0_iter3_reg <= data_31_V_read32_reg_4221_pp0_iter2_reg;
        data_31_V_read32_reg_4221_pp0_iter4_reg <= data_31_V_read32_reg_4221_pp0_iter3_reg;
        data_31_V_read32_reg_4221_pp0_iter5_reg <= data_31_V_read32_reg_4221_pp0_iter4_reg;
        data_31_V_read32_reg_4221_pp0_iter6_reg <= data_31_V_read32_reg_4221_pp0_iter5_reg;
        data_31_V_read32_reg_4221_pp0_iter7_reg <= data_31_V_read32_reg_4221_pp0_iter6_reg;
        data_31_V_read32_reg_4221_pp0_iter8_reg <= data_31_V_read32_reg_4221_pp0_iter7_reg;
        data_3_V_read_9_reg_5019 <= data_3_V_read_int_reg;
        data_3_V_read_9_reg_5019_pp0_iter1_reg <= data_3_V_read_9_reg_5019;
        data_3_V_read_9_reg_5019_pp0_iter2_reg <= data_3_V_read_9_reg_5019_pp0_iter1_reg;
        data_4_V_read_9_reg_4998 <= data_4_V_read_int_reg;
        data_4_V_read_9_reg_4998_pp0_iter1_reg <= data_4_V_read_9_reg_4998;
        data_4_V_read_9_reg_4998_pp0_iter2_reg <= data_4_V_read_9_reg_4998_pp0_iter1_reg;
        data_5_V_read_8_reg_4969 <= data_5_V_read_int_reg;
        data_5_V_read_8_reg_4969_pp0_iter1_reg <= data_5_V_read_8_reg_4969;
        data_5_V_read_8_reg_4969_pp0_iter2_reg <= data_5_V_read_8_reg_4969_pp0_iter1_reg;
        data_5_V_read_8_reg_4969_pp0_iter3_reg <= data_5_V_read_8_reg_4969_pp0_iter2_reg;
        data_6_V_read_8_reg_4944 <= data_6_V_read_int_reg;
        data_6_V_read_8_reg_4944_pp0_iter1_reg <= data_6_V_read_8_reg_4944;
        data_6_V_read_8_reg_4944_pp0_iter2_reg <= data_6_V_read_8_reg_4944_pp0_iter1_reg;
        data_6_V_read_8_reg_4944_pp0_iter3_reg <= data_6_V_read_8_reg_4944_pp0_iter2_reg;
        data_7_V_read_8_reg_4916 <= data_7_V_read_int_reg;
        data_7_V_read_8_reg_4916_pp0_iter1_reg <= data_7_V_read_8_reg_4916;
        data_7_V_read_8_reg_4916_pp0_iter2_reg <= data_7_V_read_8_reg_4916_pp0_iter1_reg;
        data_7_V_read_8_reg_4916_pp0_iter3_reg <= data_7_V_read_8_reg_4916_pp0_iter2_reg;
        data_8_V_read_7_reg_4887 <= data_8_V_read_int_reg;
        data_8_V_read_7_reg_4887_pp0_iter1_reg <= data_8_V_read_7_reg_4887;
        data_8_V_read_7_reg_4887_pp0_iter2_reg <= data_8_V_read_7_reg_4887_pp0_iter1_reg;
        data_8_V_read_7_reg_4887_pp0_iter3_reg <= data_8_V_read_7_reg_4887_pp0_iter2_reg;
        data_9_V_read_7_reg_4859 <= data_9_V_read_int_reg;
        data_9_V_read_7_reg_4859_pp0_iter1_reg <= data_9_V_read_7_reg_4859;
        data_9_V_read_7_reg_4859_pp0_iter2_reg <= data_9_V_read_7_reg_4859_pp0_iter1_reg;
        data_9_V_read_7_reg_4859_pp0_iter3_reg <= data_9_V_read_7_reg_4859_pp0_iter2_reg;
        data_9_V_read_7_reg_4859_pp0_iter4_reg <= data_9_V_read_7_reg_4859_pp0_iter3_reg;
        sub_ln703_105_reg_5226 <= sub_ln703_105_fu_489_p2;
        sub_ln703_113_reg_5247 <= sub_ln703_113_fu_533_p2;
        sub_ln703_114_reg_5253 <= sub_ln703_114_fu_549_p2;
        sub_ln703_117_reg_5259 <= sub_ln703_117_fu_554_p2;
        sub_ln703_126_reg_5274 <= sub_ln703_126_fu_574_p2;
        sub_ln703_129_reg_5279 <= sub_ln703_129_fu_579_p2;
        sub_ln703_133_reg_5284 <= sub_ln703_133_fu_584_p2;
        sub_ln703_138_reg_5325 <= sub_ln703_138_fu_816_p2;
        sub_ln703_141_reg_5330 <= sub_ln703_141_fu_835_p2;
        sub_ln703_143_reg_5335 <= sub_ln703_143_fu_844_p2;
        sub_ln703_144_reg_5340 <= sub_ln703_144_fu_858_p2;
        sub_ln703_145_reg_5345 <= sub_ln703_145_fu_863_p2;
        sub_ln703_149_reg_5350 <= sub_ln703_149_fu_901_p2;
        sub_ln703_154_reg_5355 <= sub_ln703_154_fu_920_p2;
        sub_ln703_161_reg_5365 <= sub_ln703_161_fu_960_p2;
        sub_ln703_162_reg_5370 <= sub_ln703_162_fu_980_p2;
        sub_ln703_166_reg_5375 <= sub_ln703_166_fu_1000_p2;
        sub_ln703_171_reg_5380 <= sub_ln703_171_fu_1015_p2;
        sub_ln703_173_reg_5385 <= sub_ln703_173_fu_1025_p2;
        sub_ln703_176_reg_5390 <= sub_ln703_176_fu_1040_p2;
        sub_ln703_180_reg_5395 <= sub_ln703_180_fu_1045_p2;
        sub_ln703_181_reg_5400 <= sub_ln703_181_fu_1050_p2;
        sub_ln703_182_reg_5410 <= sub_ln703_182_fu_1060_p2;
        sub_ln703_185_reg_5425 <= sub_ln703_185_fu_1095_p2;
        sub_ln703_187_reg_5440 <= sub_ln703_187_fu_1110_p2;
        sub_ln703_189_reg_5445 <= sub_ln703_189_fu_1115_p2;
        sub_ln703_191_reg_5450 <= sub_ln703_191_fu_1120_p2;
        sub_ln703_198_reg_5465 <= sub_ln703_198_fu_1146_p2;
        sub_ln703_199_reg_5470 <= sub_ln703_199_fu_1151_p2;
        sub_ln703_200_reg_5515 <= sub_ln703_200_fu_1326_p2;
        sub_ln703_203_reg_5520 <= sub_ln703_203_fu_1339_p2;
        sub_ln703_207_reg_5535 <= sub_ln703_207_fu_1384_p2;
        sub_ln703_212_reg_5540 <= sub_ln703_212_fu_1412_p2;
        sub_ln703_215_reg_5545 <= sub_ln703_215_fu_1441_p2;
        sub_ln703_229_reg_5560 <= sub_ln703_229_fu_1518_p2;
        sub_ln703_237_reg_5565 <= sub_ln703_237_fu_1571_p2;
        sub_ln703_238_reg_5570 <= sub_ln703_238_fu_1576_p2;
        sub_ln703_246_reg_5501 <= sub_ln703_246_fu_1193_p2;
        sub_ln703_252_reg_5575 <= sub_ln703_252_fu_1616_p2;
        sub_ln703_253_reg_5580 <= sub_ln703_253_fu_1621_p2;
        sub_ln703_254_reg_5585 <= sub_ln703_254_fu_1626_p2;
        sub_ln703_257_reg_5595 <= sub_ln703_257_fu_1641_p2;
        sub_ln703_261_reg_5600 <= sub_ln703_261_fu_1646_p2;
        sub_ln703_262_reg_5605 <= sub_ln703_262_fu_1651_p2;
        sub_ln703_263_reg_5610 <= sub_ln703_263_fu_1671_p2;
        sub_ln703_265_reg_5615 <= sub_ln703_265_fu_1676_p2;
        sub_ln703_266_reg_5620 <= sub_ln703_266_fu_1681_p2;
        sub_ln703_270_reg_5630 <= sub_ln703_270_fu_1695_p2;
        sub_ln703_272_reg_5635 <= sub_ln703_272_fu_1700_p2;
        sub_ln703_276_reg_5728 <= sub_ln703_276_fu_1918_p2;
        sub_ln703_278_reg_5650 <= sub_ln703_278_fu_1735_p2;
        sub_ln703_283_reg_5733 <= sub_ln703_283_fu_1975_p2;
        sub_ln703_288_reg_5738 <= sub_ln703_288_fu_2003_p2;
        sub_ln703_289_reg_5665 <= sub_ln703_289_fu_1750_p2;
        sub_ln703_290_reg_5670 <= sub_ln703_290_fu_1755_p2;
        sub_ln703_300_reg_5748 <= sub_ln703_300_fu_2075_p2;
        sub_ln703_302_reg_5758 <= sub_ln703_302_fu_2089_p2;
        sub_ln703_304_reg_5763 <= sub_ln703_304_fu_2099_p2;
        sub_ln703_309_reg_5773 <= sub_ln703_309_fu_2148_p2;
        sub_ln703_311_reg_5778 <= sub_ln703_311_fu_2173_p2;
        sub_ln703_318_reg_5783 <= sub_ln703_318_fu_2203_p2;
        sub_ln703_321_reg_5788 <= sub_ln703_321_fu_2218_p2;
        sub_ln703_323_reg_5798 <= sub_ln703_323_fu_2233_p2;
        sub_ln703_324_reg_5803 <= sub_ln703_324_fu_2238_p2;
        sub_ln703_325_reg_5808 <= sub_ln703_325_fu_2243_p2;
        sub_ln703_327_reg_5813 <= sub_ln703_327_fu_2248_p2;
        sub_ln703_328_reg_5818 <= sub_ln703_328_fu_2253_p2;
        sub_ln703_331_reg_5823 <= sub_ln703_331_fu_2258_p2;
        sub_ln703_332_reg_5828 <= sub_ln703_332_fu_2273_p2;
        sub_ln703_335_reg_5843 <= sub_ln703_335_fu_2302_p2;
        sub_ln703_343_reg_5853 <= sub_ln703_343_fu_2312_p2;
        sub_ln703_346_reg_5863 <= sub_ln703_346_fu_2332_p2;
        sub_ln703_356_reg_5921 <= sub_ln703_356_fu_2603_p2;
        sub_ln703_357_reg_5926 <= sub_ln703_357_fu_2608_p2;
        sub_ln703_361_reg_5936 <= sub_ln703_361_fu_2636_p2;
        sub_ln703_366_reg_5941 <= sub_ln703_366_fu_2684_p2;
        sub_ln703_369_reg_5946 <= sub_ln703_369_fu_2699_p2;
        sub_ln703_374_reg_5956 <= sub_ln703_374_fu_2728_p2;
        sub_ln703_375_reg_5966 <= sub_ln703_375_fu_2747_p2;
        sub_ln703_379_reg_5971 <= sub_ln703_379_fu_2781_p2;
        sub_ln703_381_reg_5976 <= sub_ln703_381_fu_2791_p2;
        sub_ln703_385_reg_5986 <= sub_ln703_385_fu_2811_p2;
        sub_ln703_386_reg_5991 <= sub_ln703_386_fu_2816_p2;
        sub_ln703_389_reg_5996 <= sub_ln703_389_fu_2839_p2;
        sub_ln703_392_reg_6001 <= sub_ln703_392_fu_2848_p2;
        sub_ln703_397_reg_6006 <= sub_ln703_397_fu_2863_p2;
        sub_ln703_402_reg_6016 <= sub_ln703_402_fu_2878_p2;
        sub_ln703_408_reg_6026 <= sub_ln703_408_fu_2893_p2;
        sub_ln703_409_reg_6031 <= sub_ln703_409_fu_2898_p2;
        sub_ln703_411_reg_6036 <= sub_ln703_411_fu_2903_p2;
        sub_ln703_416_reg_6046 <= sub_ln703_416_fu_2923_p2;
        sub_ln703_426_reg_6061 <= sub_ln703_426_fu_2938_p2;
        sub_ln703_428_reg_6108 <= sub_ln703_428_fu_3163_p2;
        sub_ln703_434_reg_6113 <= sub_ln703_434_fu_3199_p2;
        sub_ln703_448_reg_6118 <= sub_ln703_448_fu_3308_p2;
        sub_ln703_450_reg_6123 <= sub_ln703_450_fu_3318_p2;
        sub_ln703_451_reg_6143 <= sub_ln703_451_fu_3343_p2;
        sub_ln703_452_reg_6148 <= sub_ln703_452_fu_3348_p2;
        sub_ln703_453_reg_6153 <= sub_ln703_453_fu_3353_p2;
        sub_ln703_454_reg_6163 <= sub_ln703_454_fu_3368_p2;
        sub_ln703_455_reg_6168 <= sub_ln703_455_fu_3373_p2;
        sub_ln703_456_reg_6178 <= sub_ln703_456_fu_3388_p2;
        sub_ln703_457_reg_6183 <= sub_ln703_457_fu_3393_p2;
        sub_ln703_458_reg_6193 <= sub_ln703_458_fu_3408_p2;
        sub_ln703_459_reg_6198 <= sub_ln703_459_fu_3418_p2;
        sub_ln703_461_reg_6208 <= sub_ln703_461_fu_3438_p2;
        sub_ln703_469_reg_6218 <= sub_ln703_469_fu_3463_p2;
        sub_ln703_474_reg_6229 <= sub_ln703_474_fu_3482_p2;
        sub_ln703_486_reg_6244 <= sub_ln703_486_fu_3507_p2;
        sub_ln703_487_reg_6249 <= sub_ln703_487_fu_3512_p2;
        sub_ln703_491_reg_6254 <= sub_ln703_491_fu_3517_p2;
        sub_ln703_500_reg_6259 <= sub_ln703_500_fu_3522_p2;
        sub_ln703_73_reg_5059 <= sub_ln703_73_fu_286_p2;
        sub_ln703_74_reg_5065 <= sub_ln703_74_fu_292_p2;
        sub_ln703_74_reg_5065_pp0_iter2_reg <= sub_ln703_74_reg_5065;
        sub_ln703_76_reg_5071 <= sub_ln703_76_fu_300_p2;
        sub_ln703_76_reg_5071_pp0_iter2_reg <= sub_ln703_76_reg_5071;
        sub_ln703_77_reg_5084 <= sub_ln703_77_fu_308_p2;
        sub_ln703_79_reg_5125 <= sub_ln703_79_fu_337_p2;
        sub_ln703_89_reg_5166 <= sub_ln703_89_fu_402_p2;
        sub_ln703_91_reg_5172 <= sub_ln703_91_fu_411_p2;
        sub_ln703_93_reg_5200 <= sub_ln703_93_fu_442_p2;
        sub_ln703_94_reg_5205 <= sub_ln703_94_fu_446_p2;
        sub_ln703_96_reg_5210 <= sub_ln703_96_fu_456_p2;
        sub_ln703_reg_5046 <= sub_ln703_fu_274_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_ce_reg)) begin
        ap_return_0_int_reg <= add_ln703_511_fu_3847_p2;
        ap_return_10_int_reg <= acc_10_V_fu_3910_p2;
        ap_return_11_int_reg <= acc_11_V_fu_3915_p2;
        ap_return_12_int_reg <= acc_12_V_fu_3920_p2;
        ap_return_13_int_reg <= acc_13_V_fu_3925_p2;
        ap_return_14_int_reg <= acc_14_V_fu_3930_p2;
        ap_return_15_int_reg <= acc_15_V_fu_3935_p2;
        ap_return_16_int_reg <= acc_16_V_fu_3940_p2;
        ap_return_17_int_reg <= acc_17_V_fu_3953_p2;
        ap_return_18_int_reg <= acc_18_V_fu_3959_p2;
        ap_return_19_int_reg <= acc_19_V_fu_3964_p2;
        ap_return_1_int_reg <= acc_1_V_fu_3852_p2;
        ap_return_20_int_reg <= acc_20_V_fu_3969_p2;
        ap_return_21_int_reg <= acc_21_V_fu_3974_p2;
        ap_return_22_int_reg <= acc_22_V_fu_3979_p2;
        ap_return_23_int_reg <= acc_23_V_fu_3984_p2;
        ap_return_24_int_reg <= acc_24_V_fu_3989_p2;
        ap_return_25_int_reg <= acc_25_V_fu_3994_p2;
        ap_return_26_int_reg <= acc_26_V_fu_3999_p2;
        ap_return_27_int_reg <= acc_27_V_fu_4004_p2;
        ap_return_28_int_reg <= acc_28_V_fu_4009_p2;
        ap_return_29_int_reg <= acc_29_V_fu_4014_p2;
        ap_return_2_int_reg <= acc_2_V_fu_3857_p2;
        ap_return_30_int_reg <= acc_30_V_fu_4019_p2;
        ap_return_31_int_reg <= acc_31_V_fu_4024_p2;
        ap_return_3_int_reg <= acc_3_V_fu_3866_p2;
        ap_return_4_int_reg <= acc_4_V_fu_3879_p2;
        ap_return_5_int_reg <= acc_5_V_fu_3885_p2;
        ap_return_6_int_reg <= acc_6_V_fu_3890_p2;
        ap_return_7_int_reg <= acc_7_V_fu_3895_p2;
        ap_return_8_int_reg <= acc_8_V_fu_3900_p2;
        ap_return_9_int_reg <= acc_9_V_fu_3905_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_ce)) begin
        data_0_V_read_int_reg <= data_0_V_read;
        data_10_V_read_int_reg <= data_10_V_read;
        data_11_V_read_int_reg <= data_11_V_read;
        data_12_V_read_int_reg <= data_12_V_read;
        data_13_V_read_int_reg <= data_13_V_read;
        data_14_V_read_int_reg <= data_14_V_read;
        data_15_V_read_int_reg <= data_15_V_read;
        data_16_V_read_int_reg <= data_16_V_read;
        data_17_V_read_int_reg <= data_17_V_read;
        data_18_V_read_int_reg <= data_18_V_read;
        data_19_V_read_int_reg <= data_19_V_read;
        data_1_V_read_int_reg <= data_1_V_read;
        data_20_V_read_int_reg <= data_20_V_read;
        data_21_V_read_int_reg <= data_21_V_read;
        data_22_V_read_int_reg <= data_22_V_read;
        data_23_V_read_int_reg <= data_23_V_read;
        data_24_V_read_int_reg <= data_24_V_read;
        data_25_V_read_int_reg <= data_25_V_read;
        data_26_V_read_int_reg <= data_26_V_read;
        data_27_V_read_int_reg <= data_27_V_read;
        data_28_V_read_int_reg <= data_28_V_read;
        data_29_V_read_int_reg <= data_29_V_read;
        data_2_V_read_int_reg <= data_2_V_read;
        data_30_V_read_int_reg <= data_30_V_read;
        data_31_V_read_int_reg <= data_31_V_read;
        data_3_V_read_int_reg <= data_3_V_read;
        data_4_V_read_int_reg <= data_4_V_read;
        data_5_V_read_int_reg <= data_5_V_read;
        data_6_V_read_int_reg <= data_6_V_read;
        data_7_V_read_int_reg <= data_7_V_read;
        data_8_V_read_int_reg <= data_8_V_read;
        data_9_V_read_int_reg <= data_9_V_read;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_0 = ap_return_0_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_0 = add_ln703_511_fu_3847_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_1 = ap_return_1_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_1 = acc_1_V_fu_3852_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_10 = ap_return_10_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_10 = acc_10_V_fu_3910_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_11 = ap_return_11_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_11 = acc_11_V_fu_3915_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_12 = ap_return_12_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_12 = acc_12_V_fu_3920_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_13 = ap_return_13_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_13 = acc_13_V_fu_3925_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_14 = ap_return_14_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_14 = acc_14_V_fu_3930_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_15 = ap_return_15_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_15 = acc_15_V_fu_3935_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_16 = ap_return_16_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_16 = acc_16_V_fu_3940_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_17 = ap_return_17_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_17 = acc_17_V_fu_3953_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_18 = ap_return_18_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_18 = acc_18_V_fu_3959_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_19 = ap_return_19_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_19 = acc_19_V_fu_3964_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_2 = ap_return_2_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_2 = acc_2_V_fu_3857_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_20 = ap_return_20_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_20 = acc_20_V_fu_3969_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_21 = ap_return_21_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_21 = acc_21_V_fu_3974_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_22 = ap_return_22_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_22 = acc_22_V_fu_3979_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_23 = ap_return_23_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_23 = acc_23_V_fu_3984_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_24 = ap_return_24_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_24 = acc_24_V_fu_3989_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_25 = ap_return_25_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_25 = acc_25_V_fu_3994_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_26 = ap_return_26_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_26 = acc_26_V_fu_3999_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_27 = ap_return_27_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_27 = acc_27_V_fu_4004_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_28 = ap_return_28_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_28 = acc_28_V_fu_4009_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_29 = ap_return_29_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_29 = acc_29_V_fu_4014_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_3 = ap_return_3_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_3 = acc_3_V_fu_3866_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_30 = ap_return_30_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_30 = acc_30_V_fu_4019_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_31 = ap_return_31_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_31 = acc_31_V_fu_4024_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_4 = ap_return_4_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_4 = acc_4_V_fu_3879_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_5 = ap_return_5_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_5 = acc_5_V_fu_3885_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_6 = ap_return_6_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_6 = acc_6_V_fu_3890_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_7 = ap_return_7_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_7 = acc_7_V_fu_3895_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_8 = ap_return_8_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_8 = acc_8_V_fu_3900_p2;
    end
end

always @ (*) begin
    if ((1'b0 == ap_ce_reg)) begin
        ap_return_9 = ap_return_9_int_reg;
    end else if ((1'b1 == ap_ce_reg)) begin
        ap_return_9 = acc_9_V_fu_3905_p2;
    end
end

assign acc_10_V_fu_3910_p2 = (add_ln703_503_fu_3757_p2 - data_31_V_read32_reg_4221_pp0_iter8_reg);

assign acc_11_V_fu_3915_p2 = (sub_ln703_507_fu_3762_p2 - data_31_V_read32_reg_4221_pp0_iter8_reg);

assign acc_12_V_fu_3920_p2 = (sub_ln703_508_fu_3767_p2 + data_31_V_read32_reg_4221_pp0_iter8_reg);

assign acc_13_V_fu_3925_p2 = (sub_ln703_509_fu_3772_p2 - data_31_V_read32_reg_4221_pp0_iter8_reg);

assign acc_14_V_fu_3930_p2 = (add_ln703_504_fu_3777_p2 - data_31_V_read32_reg_4221_pp0_iter8_reg);

assign acc_15_V_fu_3935_p2 = (sub_ln703_510_fu_3781_p2 + data_31_V_read32_reg_4221_pp0_iter8_reg);

assign acc_16_V_fu_3940_p2 = (add_ln703_505_fu_3785_p2 - data_31_V_read32_reg_4221_pp0_iter8_reg);

assign acc_17_V_fu_3953_p2 = (add_ln703_527_fu_3949_p2 + add_ln703_526_fu_3945_p2);

assign acc_18_V_fu_3959_p2 = (sub_ln703_511_fu_3790_p2 + data_31_V_read32_reg_4221_pp0_iter8_reg);

assign acc_19_V_fu_3964_p2 = (add_ln703_509_reg_6092_pp0_iter8_reg + sub_ln703_490_fu_3675_p2);

assign acc_1_V_fu_3852_p2 = (sub_ln703_501_fu_3728_p2 + data_31_V_read32_reg_4221_pp0_iter8_reg);

assign acc_20_V_fu_3969_p2 = (add_ln703_506_fu_3795_p2 - data_31_V_read32_reg_4221_pp0_iter8_reg);

assign acc_21_V_fu_3974_p2 = (add_ln703_507_fu_3799_p2 - data_31_V_read32_reg_4221_pp0_iter8_reg);

assign acc_22_V_fu_3979_p2 = (sub_ln703_512_fu_3804_p2 + data_31_V_read32_reg_4221_pp0_iter8_reg);

assign acc_23_V_fu_3984_p2 = (sub_ln703_513_fu_3809_p2 + data_31_V_read32_reg_4221_pp0_iter8_reg);

assign acc_24_V_fu_3989_p2 = (sub_ln703_514_fu_3814_p2 + data_31_V_read32_reg_4221_pp0_iter8_reg);

assign acc_25_V_fu_3994_p2 = (sub_ln703_515_fu_3819_p2 + data_31_V_read32_reg_4221_pp0_iter8_reg);

assign acc_26_V_fu_3999_p2 = (add_ln703_509_reg_6092_pp0_iter8_reg + sub_ln703_497_fu_3704_p2);

assign acc_27_V_fu_4004_p2 = (sub_ln703_516_fu_3824_p2 - data_31_V_read32_reg_4221_pp0_iter8_reg);

assign acc_28_V_fu_4009_p2 = (sub_ln703_517_fu_3829_p2 + data_31_V_read32_reg_4221_pp0_iter8_reg);

assign acc_29_V_fu_4014_p2 = (add_ln703_509_reg_6092_pp0_iter8_reg + sub_ln703_498_fu_3718_p2);

assign acc_2_V_fu_3857_p2 = (sub_ln703_502_fu_3732_p2 + data_31_V_read32_reg_4221_pp0_iter8_reg);

assign acc_30_V_fu_4019_p2 = (sub_ln703_518_fu_3834_p2 - data_31_V_read32_reg_4221_pp0_iter8_reg);

assign acc_31_V_fu_4024_p2 = (sub_ln703_519_fu_3839_p2 - data_31_V_read32_reg_4221_pp0_iter8_reg);

assign acc_3_V_fu_3866_p2 = (add_ln703_509_reg_6092_pp0_iter8_reg + add_ln703_514_fu_3862_p2);

assign acc_4_V_fu_3879_p2 = (add_ln703_518_fu_3875_p2 + add_ln703_517_fu_3871_p2);

assign acc_5_V_fu_3885_p2 = (sub_ln703_503_fu_3737_p2 + data_31_V_read32_reg_4221_pp0_iter8_reg);

assign acc_6_V_fu_3890_p2 = (sub_ln703_504_fu_3742_p2 - data_31_V_read32_reg_4221_pp0_iter8_reg);

assign acc_7_V_fu_3895_p2 = (sub_ln703_505_fu_3747_p2 + data_31_V_read32_reg_4221_pp0_iter8_reg);

assign acc_8_V_fu_3900_p2 = (add_ln703_509_reg_6092_pp0_iter8_reg + sub_ln703_481_fu_3636_p2);

assign acc_9_V_fu_3905_p2 = (sub_ln703_506_fu_3752_p2 + data_31_V_read32_reg_4221_pp0_iter8_reg);

assign add_ln703_200_fu_304_p2 = (add_ln703_reg_5052 + data_2_V_read_9_reg_5035);

assign add_ln703_201_fu_312_p2 = (sub_ln703_reg_5046 + data_2_V_read_9_reg_5035);

assign add_ln703_202_fu_316_p2 = (sub_ln703_73_reg_5059 + data_2_V_read_9_reg_5035);

assign add_ln703_203_fu_329_p2 = (sub_ln703_74_reg_5065 + data_3_V_read_9_reg_5019_pp0_iter1_reg);

assign add_ln703_204_fu_320_p2 = (sub_ln703_75_fu_296_p2 + data_3_V_read_9_reg_5019);

assign add_ln703_205_fu_333_p2 = (add_ln703_200_reg_5077 + data_3_V_read_9_reg_5019_pp0_iter1_reg);

assign add_ln703_206_fu_341_p2 = (sub_ln703_76_reg_5071 + data_3_V_read_9_reg_5019_pp0_iter1_reg);

assign add_ln703_207_fu_325_p2 = (data_3_V_read_9_reg_5019 + data_4_V_read_9_reg_4998);

assign add_ln703_208_fu_345_p2 = (add_ln703_207_reg_5107 + sub_ln703_77_reg_5084);

assign add_ln703_209_fu_416_p2 = (add_ln703_205_reg_5119 + data_4_V_read_9_reg_4998_pp0_iter2_reg);

assign add_ln703_210_fu_349_p2 = (add_ln703_204_reg_5101 + data_4_V_read_9_reg_4998_pp0_iter1_reg);

assign add_ln703_211_fu_420_p2 = (sub_ln703_82_fu_373_p2 + data_4_V_read_9_reg_4998_pp0_iter2_reg);

assign add_ln703_212_fu_425_p2 = (add_ln703_203_reg_5113 + data_4_V_read_9_reg_4998_pp0_iter2_reg);

assign add_ln703_213_fu_429_p2 = (add_ln703_207_reg_5107_pp0_iter2_reg + add_ln703_201_reg_5090_pp0_iter2_reg);

assign add_ln703_214_fu_433_p2 = (add_ln703_206_reg_5131 + data_4_V_read_9_reg_4998_pp0_iter2_reg);

assign add_ln703_215_fu_605_p2 = (sub_ln703_89_reg_5166 + data_5_V_read_8_reg_4969_pp0_iter3_reg);

assign add_ln703_216_fu_461_p2 = (sub_ln703_90_fu_406_p2 + data_5_V_read_8_reg_4969_pp0_iter2_reg);

assign add_ln703_217_fu_470_p2 = (add_ln703_210_reg_5143 + data_5_V_read_8_reg_4969_pp0_iter2_reg);

assign add_ln703_218_fu_474_p2 = (add_ln703_211_fu_420_p2 + data_5_V_read_8_reg_4969_pp0_iter2_reg);

assign add_ln703_219_fu_479_p2 = (add_ln703_212_fu_425_p2 + data_5_V_read_8_reg_4969_pp0_iter2_reg);

assign add_ln703_220_fu_484_p2 = (sub_ln703_87_fu_393_p2 + data_5_V_read_8_reg_4969_pp0_iter2_reg);

assign add_ln703_221_fu_499_p2 = (add_ln703_208_reg_5137 + data_5_V_read_8_reg_4969_pp0_iter2_reg);

assign add_ln703_222_fu_503_p2 = (data_5_V_read_8_reg_4969_pp0_iter2_reg + data_6_V_read_8_reg_4944_pp0_iter2_reg);

assign add_ln703_223_fu_507_p2 = (add_ln703_222_fu_503_p2 + sub_ln703_85_fu_385_p2);

assign add_ln703_224_fu_645_p2 = (sub_ln703_96_reg_5210 + data_6_V_read_8_reg_4944_pp0_iter3_reg);

assign add_ln703_225_fu_513_p2 = (sub_ln703_98_fu_466_p2 + data_6_V_read_8_reg_4944_pp0_iter2_reg);

assign add_ln703_226_fu_518_p2 = (sub_ln703_79_reg_5125 + data_4_V_read_9_reg_4998_pp0_iter2_reg);

assign add_ln703_227_fu_522_p2 = (add_ln703_222_fu_503_p2 + add_ln703_226_fu_518_p2);

assign add_ln703_228_fu_663_p2 = (sub_ln703_99_fu_613_p2 + data_6_V_read_8_reg_4944_pp0_iter3_reg);

assign add_ln703_229_fu_668_p2 = (sub_ln703_100_fu_617_p2 + data_6_V_read_8_reg_4944_pp0_iter3_reg);

assign add_ln703_230_fu_538_p2 = (sub_ln703_83_fu_377_p2 + data_4_V_read_9_reg_4998_pp0_iter2_reg);

assign add_ln703_231_fu_543_p2 = (add_ln703_222_fu_503_p2 + add_ln703_230_fu_538_p2);

assign add_ln703_232_fu_673_p2 = (sub_ln703_101_fu_621_p2 + data_6_V_read_8_reg_4944_pp0_iter3_reg);

assign add_ln703_233_fu_353_p2 = (data_6_V_read_8_reg_4944_pp0_iter1_reg + data_7_V_read_8_reg_4916_pp0_iter1_reg);

assign add_ln703_234_fu_564_p2 = (add_ln703_233_reg_5149 + sub_ln703_95_fu_451_p2);

assign add_ln703_235_fu_701_p2 = (add_ln703_223_reg_5231 + data_7_V_read_8_reg_4916_pp0_iter3_reg);

assign add_ln703_236_fu_710_p2 = (sub_ln703_111_fu_658_p2 + data_7_V_read_8_reg_4916_pp0_iter3_reg);

assign add_ln703_237_fu_715_p2 = (add_ln703_233_reg_5149_pp0_iter3_reg + add_ln703_216_reg_5215);

assign add_ln703_238_fu_569_p2 = (add_ln703_233_reg_5149 + sub_ln703_94_fu_446_p2);

assign add_ln703_239_fu_750_p2 = (add_ln703_233_reg_5149_pp0_iter3_reg + sub_ln703_102_fu_625_p2);

assign add_ln703_240_fu_755_p2 = (sub_ln703_115_fu_678_p2 + data_7_V_read_8_reg_4916_pp0_iter3_reg);

assign add_ln703_241_fu_765_p2 = (sub_ln703_117_reg_5259 + data_7_V_read_8_reg_4916_pp0_iter3_reg);

assign add_ln703_242_fu_769_p2 = (add_ln703_233_reg_5149_pp0_iter3_reg + sub_ln703_107_fu_637_p2);

assign add_ln703_243_fu_774_p2 = (add_ln703_209_reg_5178 + data_5_V_read_8_reg_4969_pp0_iter3_reg);

assign add_ln703_244_fu_778_p2 = (add_ln703_233_reg_5149_pp0_iter3_reg + add_ln703_243_fu_774_p2);

assign add_ln703_245_fu_783_p2 = (sub_ln703_114_reg_5253 + data_7_V_read_8_reg_4916_pp0_iter3_reg);

assign add_ln703_246_fu_787_p2 = (sub_ln703_119_fu_687_p2 + data_8_V_read_7_reg_4887_pp0_iter3_reg);

assign add_ln703_247_fu_357_p2 = (data_7_V_read_8_reg_4916_pp0_iter1_reg + data_8_V_read_7_reg_4887_pp0_iter1_reg);

assign add_ln703_248_fu_801_p2 = (add_ln703_247_reg_5159_pp0_iter3_reg + sub_ln703_109_fu_649_p2);

assign add_ln703_249_fu_830_p2 = (sub_ln703_123_fu_719_p2 + data_8_V_read_7_reg_4887_pp0_iter3_reg);

assign add_ln703_250_fu_849_p2 = (sub_ln703_91_reg_5172 + data_5_V_read_8_reg_4969_pp0_iter3_reg);

assign add_ln703_251_fu_589_p2 = (add_ln703_247_reg_5159 + data_6_V_read_8_reg_4944_pp0_iter2_reg);

assign add_ln703_252_fu_853_p2 = (add_ln703_251_reg_5289 + add_ln703_250_fu_849_p2);

assign add_ln703_253_fu_873_p2 = (sub_ln703_105_reg_5226 + data_6_V_read_8_reg_4944_pp0_iter3_reg);

assign add_ln703_254_fu_877_p2 = (add_ln703_247_reg_5159_pp0_iter3_reg + add_ln703_253_fu_873_p2);

assign add_ln703_255_fu_887_p2 = (add_ln703_214_reg_5194 + data_5_V_read_8_reg_4969_pp0_iter3_reg);

assign add_ln703_256_fu_891_p2 = (add_ln703_251_reg_5289 + add_ln703_255_fu_887_p2);

assign add_ln703_257_fu_925_p2 = (sub_ln703_139_fu_821_p2 + data_9_V_read_7_reg_4859_pp0_iter3_reg);

assign add_ln703_258_fu_593_p2 = (data_8_V_read_7_reg_4887_pp0_iter2_reg + data_9_V_read_7_reg_4859_pp0_iter2_reg);

assign add_ln703_259_fu_940_p2 = (add_ln703_258_reg_5295 + sub_ln703_124_fu_723_p2);

assign add_ln703_260_fu_950_p2 = (add_ln703_258_reg_5295 + sub_ln703_127_fu_732_p2);

assign add_ln703_261_fu_955_p2 = (add_ln703_258_reg_5295 + sub_ln703_131_fu_745_p2);

assign add_ln703_262_fu_965_p2 = (sub_ln703_104_fu_633_p2 + data_6_V_read_8_reg_4944_pp0_iter3_reg);

assign add_ln703_263_fu_970_p2 = (add_ln703_258_reg_5295 + data_7_V_read_8_reg_4916_pp0_iter3_reg);

assign add_ln703_264_fu_974_p2 = (add_ln703_263_fu_970_p2 + add_ln703_262_fu_965_p2);

assign add_ln703_265_fu_1010_p2 = (sub_ln703_153_fu_915_p2 + data_10_V_read11_reg_4832_pp0_iter3_reg);

assign add_ln703_266_fu_1232_p2 = (sub_ln703_158_fu_1210_p2 + data_10_V_read11_reg_4832_pp0_iter4_reg);

assign add_ln703_267_fu_1055_p2 = (sub_ln703_164_fu_990_p2 + data_10_V_read11_reg_4832_pp0_iter3_reg);

assign add_ln703_268_fu_1065_p2 = (data_9_V_read_7_reg_4859_pp0_iter3_reg + data_10_V_read11_reg_4832_pp0_iter3_reg);

assign add_ln703_269_fu_1069_p2 = (add_ln703_268_fu_1065_p2 + sub_ln703_150_fu_906_p2);

assign add_ln703_270_fu_1255_p2 = (sub_ln703_169_fu_1222_p2 + data_11_V_read12_reg_4808_pp0_iter4_reg);

assign add_ln703_271_fu_1080_p2 = (sub_ln703_120_fu_691_p2 + data_8_V_read_7_reg_4887_pp0_iter3_reg);

assign add_ln703_272_fu_597_p2 = (data_10_V_read11_reg_4832_pp0_iter2_reg + data_11_V_read12_reg_4808_pp0_iter2_reg);

assign add_ln703_273_fu_1085_p2 = (add_ln703_272_reg_5304 + data_9_V_read_7_reg_4859_pp0_iter3_reg);

assign add_ln703_274_fu_1089_p2 = (add_ln703_273_fu_1085_p2 + add_ln703_271_fu_1080_p2);

assign add_ln703_275_fu_1260_p2 = (add_ln703_272_reg_5304_pp0_iter4_reg + sub_ln703_154_reg_5355);

assign add_ln703_276_fu_1100_p2 = (sub_ln703_136_fu_806_p2 + data_9_V_read_7_reg_4859_pp0_iter3_reg);

assign add_ln703_277_fu_1264_p2 = (add_ln703_272_reg_5304_pp0_iter4_reg + add_ln703_276_reg_5430);

assign add_ln703_278_fu_1105_p2 = (sub_ln703_137_fu_811_p2 + data_9_V_read_7_reg_4859_pp0_iter3_reg);

assign add_ln703_279_fu_1268_p2 = (add_ln703_272_reg_5304_pp0_iter4_reg + add_ln703_278_reg_5435);

assign add_ln703_280_fu_1125_p2 = (sub_ln703_129_reg_5279 + data_8_V_read_7_reg_4887_pp0_iter3_reg);

assign add_ln703_281_fu_1129_p2 = (add_ln703_273_fu_1085_p2 + add_ln703_280_fu_1125_p2);

assign add_ln703_282_fu_1135_p2 = (sub_ln703_130_fu_741_p2 + data_8_V_read_7_reg_4887_pp0_iter3_reg);

assign add_ln703_283_fu_1140_p2 = (add_ln703_273_fu_1085_p2 + add_ln703_282_fu_1135_p2);

assign add_ln703_284_fu_1296_p2 = (sub_ln703_145_reg_5345 + data_9_V_read_7_reg_4859_pp0_iter4_reg);

assign add_ln703_285_fu_1300_p2 = (add_ln703_272_reg_5304_pp0_iter4_reg + add_ln703_284_fu_1296_p2);

assign add_ln703_286_fu_1305_p2 = (sub_ln703_180_reg_5395 + data_11_V_read12_reg_4808_pp0_iter4_reg);

assign add_ln703_287_fu_1354_p2 = (sub_ln703_186_fu_1272_p2 + data_12_V_read13_reg_4778_pp0_iter4_reg);

assign add_ln703_288_fu_1156_p2 = (data_11_V_read12_reg_4808_pp0_iter3_reg + data_12_V_read13_reg_4778_pp0_iter3_reg);

assign add_ln703_289_fu_1359_p2 = (add_ln703_288_reg_5475 + sub_ln703_171_reg_5380);

assign add_ln703_290_fu_1367_p2 = (sub_ln703_189_reg_5445 + data_12_V_read13_reg_4778_pp0_iter4_reg);

assign add_ln703_291_fu_1371_p2 = (sub_ln703_190_fu_1281_p2 + data_12_V_read13_reg_4778_pp0_iter4_reg);

assign add_ln703_292_fu_1376_p2 = (sub_ln703_191_reg_5450 + data_12_V_read13_reg_4778_pp0_iter4_reg);

assign add_ln703_293_fu_1380_p2 = (add_ln703_288_reg_5475 + sub_ln703_176_reg_5390);

assign add_ln703_294_fu_1397_p2 = (add_ln703_288_reg_5475 + sub_ln703_178_fu_1242_p2);

assign add_ln703_295_fu_1427_p2 = (sub_ln703_196_fu_1317_p2 + data_12_V_read13_reg_4778_pp0_iter4_reg);

assign add_ln703_296_fu_1432_p2 = (sub_ln703_166_reg_5375 + data_10_V_read11_reg_4832_pp0_iter4_reg);

assign add_ln703_297_fu_1436_p2 = (add_ln703_288_reg_5475 + add_ln703_296_fu_1432_p2);

assign add_ln703_298_fu_1454_p2 = (sub_ln703_202_fu_1335_p2 + data_13_V_read14_reg_4745_pp0_iter4_reg);

assign add_ln703_299_fu_1464_p2 = (sub_ln703_205_fu_1349_p2 + data_13_V_read14_reg_4745_pp0_iter4_reg);

assign add_ln703_300_fu_1474_p2 = (sub_ln703_206_fu_1363_p2 + data_13_V_read14_reg_4745_pp0_iter4_reg);

assign add_ln703_301_fu_1494_p2 = (sub_ln703_208_fu_1389_p2 + data_13_V_read14_reg_4745_pp0_iter4_reg);

assign add_ln703_302_fu_1160_p2 = (sub_ln703_113_reg_5247 + data_7_V_read_8_reg_4916_pp0_iter3_reg);

assign add_ln703_303_fu_1164_p2 = (add_ln703_258_reg_5295 + add_ln703_302_fu_1160_p2);

assign add_ln703_304_fu_601_p2 = (data_12_V_read13_reg_4778_pp0_iter2_reg + data_13_V_read14_reg_4745_pp0_iter2_reg);

assign add_ln703_305_fu_1169_p2 = (add_ln703_304_reg_5314 + add_ln703_272_reg_5304);

assign add_ln703_306_fu_1173_p2 = (add_ln703_305_fu_1169_p2 + add_ln703_303_fu_1164_p2);

assign add_ln703_307_fu_1504_p2 = (sub_ln703_210_fu_1402_p2 + data_13_V_read14_reg_4745_pp0_iter4_reg);

assign add_ln703_308_fu_1509_p2 = (add_ln703_268_reg_5415 + sub_ln703_144_reg_5340);

assign add_ln703_309_fu_1179_p2 = (add_ln703_304_reg_5314 + data_11_V_read12_reg_4808_pp0_iter3_reg);

assign add_ln703_310_fu_1513_p2 = (add_ln703_309_reg_5484 + add_ln703_308_fu_1509_p2);

assign add_ln703_311_fu_1523_p2 = (sub_ln703_162_reg_5370 + data_10_V_read11_reg_4832_pp0_iter4_reg);

assign add_ln703_312_fu_1527_p2 = (add_ln703_309_reg_5484 + add_ln703_311_fu_1523_p2);

assign add_ln703_313_fu_1532_p2 = (sub_ln703_213_fu_1417_p2 + data_13_V_read14_reg_4745_pp0_iter4_reg);

assign add_ln703_314_fu_1183_p2 = (data_13_V_read14_reg_4745_pp0_iter3_reg + data_14_V_read15_reg_4714_pp0_iter3_reg);

assign add_ln703_315_fu_1552_p2 = (add_ln703_314_reg_5490 + sub_ln703_201_fu_1331_p2);

assign add_ln703_316_fu_1187_p2 = (add_ln703_268_fu_1065_p2 + sub_ln703_135_fu_796_p2);

assign add_ln703_317_fu_1562_p2 = (add_ln703_314_reg_5490 + add_ln703_288_reg_5475);

assign add_ln703_318_fu_1566_p2 = (add_ln703_317_fu_1562_p2 + add_ln703_316_reg_5496);

assign add_ln703_319_fu_1591_p2 = (sub_ln703_223_fu_1479_p2 + data_14_V_read15_reg_4714_pp0_iter4_reg);

assign add_ln703_320_fu_1822_p2 = (sub_ln703_224_fu_1796_p2 + data_14_V_read15_reg_4714_pp0_iter5_reg);

assign add_ln703_321_fu_1636_p2 = (sub_ln703_236_fu_1557_p2 + data_15_V_read16_reg_4682_pp0_iter4_reg);

assign add_ln703_322_fu_1656_p2 = (sub_ln703_188_fu_1277_p2 + data_12_V_read13_reg_4778_pp0_iter4_reg);

assign add_ln703_323_fu_1198_p2 = (data_14_V_read15_reg_4714_pp0_iter3_reg + data_15_V_read16_reg_4682_pp0_iter3_reg);

assign add_ln703_324_fu_1661_p2 = (add_ln703_323_reg_5506 + data_13_V_read14_reg_4745_pp0_iter4_reg);

assign add_ln703_325_fu_1665_p2 = (add_ln703_324_fu_1661_p2 + add_ln703_322_fu_1656_p2);

assign add_ln703_326_fu_1686_p2 = (add_ln703_323_reg_5506 + sub_ln703_228_fu_1499_p2);

assign add_ln703_327_fu_1887_p2 = (sub_ln703_250_fu_1844_p2 + data_15_V_read16_reg_4682_pp0_iter5_reg);

assign add_ln703_328_fu_1892_p2 = (sub_ln703_252_reg_5575 + data_15_V_read16_reg_4682_pp0_iter5_reg);

assign add_ln703_329_fu_1705_p2 = (sub_ln703_214_fu_1422_p2 + data_13_V_read14_reg_4745_pp0_iter4_reg);

assign add_ln703_330_fu_1710_p2 = (add_ln703_323_reg_5506 + add_ln703_329_fu_1705_p2);

assign add_ln703_331_fu_1900_p2 = (sub_ln703_254_reg_5585 + data_15_V_read16_reg_4682_pp0_iter5_reg);

assign add_ln703_332_fu_1715_p2 = (sub_ln703_216_fu_1446_p2 + data_13_V_read14_reg_4745_pp0_iter4_reg);

assign add_ln703_333_fu_1720_p2 = (add_ln703_323_reg_5506 + add_ln703_332_fu_1715_p2);

assign add_ln703_334_fu_1725_p2 = (add_ln703_323_reg_5506 + sub_ln703_234_fu_1547_p2);

assign add_ln703_335_fu_1730_p2 = (sub_ln703_256_fu_1631_p2 + data_16_V_read17_reg_4650_pp0_iter4_reg);

assign add_ln703_336_fu_1913_p2 = (sub_ln703_258_fu_1854_p2 + data_16_V_read17_reg_4650_pp0_iter5_reg);

assign add_ln703_337_fu_1923_p2 = (sub_ln703_261_reg_5600 + data_16_V_read17_reg_4650_pp0_iter5_reg);

assign add_ln703_338_fu_1939_p2 = (sub_ln703_266_reg_5620 + data_16_V_read17_reg_4650_pp0_iter5_reg);

assign add_ln703_339_fu_1740_p2 = (sub_ln703_209_fu_1393_p2 + data_13_V_read14_reg_4745_pp0_iter4_reg);

assign add_ln703_340_fu_1943_p2 = (data_15_V_read16_reg_4682_pp0_iter5_reg + data_16_V_read17_reg_4650_pp0_iter5_reg);

assign add_ln703_341_fu_1947_p2 = (add_ln703_340_fu_1943_p2 + data_14_V_read15_reg_4714_pp0_iter5_reg);

assign add_ln703_342_fu_1952_p2 = (add_ln703_341_fu_1947_p2 + add_ln703_339_reg_5655);

assign add_ln703_343_fu_1745_p2 = (sub_ln703_268_fu_1691_p2 + data_16_V_read17_reg_4650_pp0_iter4_reg);

assign add_ln703_344_fu_1966_p2 = (sub_ln703_270_reg_5630 + data_16_V_read17_reg_4650_pp0_iter5_reg);

assign add_ln703_345_fu_1970_p2 = (sub_ln703_271_fu_1882_p2 + data_16_V_read17_reg_4650_pp0_iter5_reg);

assign add_ln703_346_fu_1993_p2 = (sub_ln703_273_fu_1896_p2 + data_16_V_read17_reg_4650_pp0_iter5_reg);

assign add_ln703_347_fu_1760_p2 = (data_16_V_read17_reg_4650_pp0_iter4_reg + data_17_V_read_8_reg_4621_pp0_iter4_reg);

assign add_ln703_348_fu_2017_p2 = (add_ln703_347_reg_5675 + sub_ln703_257_reg_5595);

assign add_ln703_349_fu_2021_p2 = (sub_ln703_219_fu_1788_p2 + data_14_V_read15_reg_4714_pp0_iter5_reg);

assign add_ln703_350_fu_2026_p2 = (add_ln703_347_reg_5675 + data_15_V_read16_reg_4682_pp0_iter5_reg);

assign add_ln703_351_fu_2030_p2 = (add_ln703_350_fu_2026_p2 + add_ln703_349_fu_2021_p2);

assign add_ln703_352_fu_2051_p2 = (sub_ln703_278_reg_5650 + data_17_V_read_8_reg_4621_pp0_iter5_reg);

assign add_ln703_353_fu_2060_p2 = (add_ln703_347_reg_5675 + sub_ln703_264_fu_1867_p2);

assign add_ln703_354_fu_2080_p2 = (sub_ln703_281_fu_1957_p2 + data_17_V_read_8_reg_4621_pp0_iter5_reg);

assign add_ln703_355_fu_2114_p2 = (sub_ln703_290_reg_5670 + data_17_V_read_8_reg_4621_pp0_iter5_reg);

assign add_ln703_356_fu_2118_p2 = (sub_ln703_235_fu_1812_p2 + data_15_V_read16_reg_4682_pp0_iter5_reg);

assign add_ln703_357_fu_1764_p2 = (data_17_V_read_8_reg_4621_pp0_iter4_reg + data_18_V_read_7_reg_4594_pp0_iter4_reg);

assign add_ln703_358_fu_2123_p2 = (add_ln703_357_reg_5683 + data_16_V_read17_reg_4650_pp0_iter5_reg);

assign add_ln703_359_fu_2127_p2 = (add_ln703_358_fu_2123_p2 + add_ln703_356_fu_2118_p2);

assign add_ln703_360_fu_2138_p2 = (sub_ln703_292_fu_2012_p2 + data_18_V_read_7_reg_4594_pp0_iter5_reg);

assign add_ln703_361_fu_2153_p2 = (sub_ln703_259_fu_1858_p2 + data_16_V_read17_reg_4650_pp0_iter5_reg);

assign add_ln703_362_fu_2158_p2 = (add_ln703_357_reg_5683 + add_ln703_361_fu_2153_p2);

assign add_ln703_363_fu_2163_p2 = (sub_ln703_295_fu_2041_p2 + data_18_V_read_7_reg_4594_pp0_iter5_reg);

assign add_ln703_364_fu_2178_p2 = (sub_ln703_297_fu_2055_p2 + data_18_V_read_7_reg_4594_pp0_iter5_reg);

assign add_ln703_365_fu_2183_p2 = (sub_ln703_298_fu_2065_p2 + data_18_V_read_7_reg_4594_pp0_iter5_reg);

assign add_ln703_366_fu_2193_p2 = (sub_ln703_303_fu_2094_p2 + data_18_V_read_7_reg_4594_pp0_iter5_reg);

assign add_ln703_367_fu_2198_p2 = (sub_ln703_305_fu_2104_p2 + data_18_V_read_7_reg_4594_pp0_iter5_reg);

assign add_ln703_368_fu_2429_p2 = (add_ln703_357_reg_5683_pp0_iter6_reg + sub_ln703_288_reg_5738);

assign add_ln703_369_fu_2213_p2 = (sub_ln703_307_fu_2133_p2 + data_19_V_read_7_reg_4567_pp0_iter5_reg);

assign add_ln703_370_fu_2437_p2 = (sub_ln703_309_reg_5773 + data_19_V_read_7_reg_4567_pp0_iter6_reg);

assign add_ln703_371_fu_1768_p2 = (data_18_V_read_7_reg_4594_pp0_iter4_reg + data_19_V_read_7_reg_4567_pp0_iter4_reg);

assign add_ln703_372_fu_2228_p2 = (add_ln703_371_reg_5691 + sub_ln703_293_fu_2036_p2);

assign add_ln703_373_fu_2445_p2 = (sub_ln703_313_fu_2413_p2 + data_19_V_read_7_reg_4567_pp0_iter6_reg);

assign add_ln703_374_fu_2263_p2 = (sub_ln703_284_fu_1980_p2 + data_17_V_read_8_reg_4621_pp0_iter5_reg);

assign add_ln703_375_fu_2268_p2 = (add_ln703_371_reg_5691 + add_ln703_374_fu_2263_p2);

assign add_ln703_376_fu_2278_p2 = (sub_ln703_287_fu_1998_p2 + data_17_V_read_8_reg_4621_pp0_iter5_reg);

assign add_ln703_377_fu_2283_p2 = (add_ln703_371_reg_5691 + add_ln703_376_fu_2278_p2);

assign add_ln703_378_fu_2288_p2 = (sub_ln703_289_reg_5665 + data_17_V_read_8_reg_4621_pp0_iter5_reg);

assign add_ln703_379_fu_2292_p2 = (add_ln703_371_reg_5691 + add_ln703_378_fu_2288_p2);

assign add_ln703_380_fu_2297_p2 = (sub_ln703_319_fu_2208_p2 + data_19_V_read_7_reg_4567_pp0_iter5_reg);

assign add_ln703_381_fu_2307_p2 = (sub_ln703_322_fu_2223_p2 + data_20_V_read21_reg_4539_pp0_iter5_reg);

assign add_ln703_382_fu_2486_p2 = (sub_ln703_325_reg_5808 + data_20_V_read21_reg_4539_pp0_iter6_reg);

assign add_ln703_383_fu_2490_p2 = (sub_ln703_326_fu_2441_p2 + data_20_V_read21_reg_4539_pp0_iter6_reg);

assign add_ln703_384_fu_1772_p2 = (data_19_V_read_7_reg_4567_pp0_iter4_reg + data_20_V_read21_reg_4539_pp0_iter4_reg);

assign add_ln703_385_fu_2499_p2 = (add_ln703_384_reg_5701_pp0_iter6_reg + sub_ln703_312_fu_2409_p2);

assign add_ln703_386_fu_2514_p2 = (sub_ln703_331_reg_5823 + data_20_V_read21_reg_4539_pp0_iter6_reg);

assign add_ln703_387_fu_2518_p2 = (add_ln703_384_reg_5701_pp0_iter6_reg + sub_ln703_317_fu_2425_p2);

assign add_ln703_388_fu_2317_p2 = (sub_ln703_285_fu_1984_p2 + data_17_V_read_8_reg_4621_pp0_iter5_reg);

assign add_ln703_389_fu_2322_p2 = (add_ln703_384_reg_5701 + data_18_V_read_7_reg_4594_pp0_iter5_reg);

assign add_ln703_390_fu_2326_p2 = (add_ln703_389_fu_2322_p2 + add_ln703_388_fu_2317_p2);

assign add_ln703_391_fu_2527_p2 = (sub_ln703_334_fu_2464_p2 + data_20_V_read21_reg_4539_pp0_iter6_reg);

assign add_ln703_392_fu_2540_p2 = (sub_ln703_336_fu_2469_p2 + data_21_V_read22_reg_4512_pp0_iter6_reg);

assign add_ln703_393_fu_2559_p2 = (sub_ln703_294_fu_2405_p2 + data_18_V_read_7_reg_4594_pp0_iter6_reg);

assign add_ln703_394_fu_1776_p2 = (data_20_V_read21_reg_4539_pp0_iter4_reg + data_21_V_read22_reg_4512_pp0_iter4_reg);

assign add_ln703_395_fu_2564_p2 = (add_ln703_394_reg_5710_pp0_iter6_reg + data_19_V_read_7_reg_4567_pp0_iter6_reg);

assign add_ln703_396_fu_2568_p2 = (add_ln703_395_fu_2564_p2 + add_ln703_393_fu_2559_p2);

assign add_ln703_397_fu_2599_p2 = (add_ln703_394_reg_5710_pp0_iter6_reg + sub_ln703_328_reg_5818);

assign add_ln703_398_fu_2337_p2 = (add_ln703_347_reg_5675 + sub_ln703_267_fu_1872_p2);

assign add_ln703_399_fu_2342_p2 = (add_ln703_394_reg_5710 + add_ln703_371_reg_5691);

assign add_ln703_400_fu_2346_p2 = (add_ln703_399_fu_2342_p2 + add_ln703_398_fu_2337_p2);

assign add_ln703_401_fu_2623_p2 = (sub_ln703_343_reg_5853 + data_21_V_read22_reg_4512_pp0_iter6_reg);

assign add_ln703_402_fu_2631_p2 = (sub_ln703_344_fu_2523_p2 + data_21_V_read22_reg_4512_pp0_iter6_reg);

assign add_ln703_403_fu_2645_p2 = (sub_ln703_320_fu_2433_p2 + data_20_V_read21_reg_4539_pp0_iter6_reg);

assign add_ln703_404_fu_1780_p2 = (data_21_V_read22_reg_4512_pp0_iter4_reg + data_22_V_read23_reg_4483_pp0_iter4_reg);

assign add_ln703_405_fu_2650_p2 = (add_ln703_404_reg_5718_pp0_iter6_reg + add_ln703_403_fu_2645_p2);

assign add_ln703_406_fu_2655_p2 = (sub_ln703_347_fu_2536_p2 + data_22_V_read23_reg_4483_pp0_iter6_reg);

assign add_ln703_407_fu_2675_p2 = (sub_ln703_323_reg_5798 + data_20_V_read21_reg_4539_pp0_iter6_reg);

assign add_ln703_408_fu_2679_p2 = (add_ln703_404_reg_5718_pp0_iter6_reg + add_ln703_407_fu_2675_p2);

assign add_ln703_409_fu_2704_p2 = (sub_ln703_354_fu_2589_p2 + data_22_V_read23_reg_4483_pp0_iter6_reg);

assign add_ln703_410_fu_2709_p2 = (sub_ln703_355_fu_2594_p2 + data_22_V_read23_reg_4483_pp0_iter6_reg);

assign add_ln703_411_fu_2352_p2 = (add_ln703_371_reg_5691 + sub_ln703_299_fu_2070_p2);

assign add_ln703_412_fu_2357_p2 = (add_ln703_404_reg_5718 + data_20_V_read21_reg_4539_pp0_iter5_reg);

assign add_ln703_413_fu_2361_p2 = (add_ln703_412_fu_2357_p2 + add_ln703_411_fu_2352_p2);

assign add_ln703_414_fu_2367_p2 = (sub_ln703_315_fu_2188_p2 + data_19_V_read_7_reg_4567_pp0_iter5_reg);

assign add_ln703_415_fu_2372_p2 = (add_ln703_412_fu_2357_p2 + add_ln703_414_fu_2367_p2);

assign add_ln703_416_fu_2733_p2 = (add_ln703_357_reg_5683_pp0_iter6_reg + sub_ln703_283_reg_5733);

assign add_ln703_417_fu_2737_p2 = (add_ln703_404_reg_5718_pp0_iter6_reg + add_ln703_384_reg_5701_pp0_iter6_reg);

assign add_ln703_418_fu_2741_p2 = (add_ln703_417_fu_2737_p2 + add_ln703_416_fu_2733_p2);

assign add_ln703_419_fu_2757_p2 = (sub_ln703_332_reg_5828 + data_20_V_read21_reg_4539_pp0_iter6_reg);

assign add_ln703_420_fu_2761_p2 = (add_ln703_404_reg_5718_pp0_iter6_reg + add_ln703_419_fu_2757_p2);

assign add_ln703_421_fu_2766_p2 = (sub_ln703_333_fu_2460_p2 + data_20_V_read21_reg_4539_pp0_iter6_reg);

assign add_ln703_422_fu_2771_p2 = (add_ln703_404_reg_5718_pp0_iter6_reg + add_ln703_421_fu_2766_p2);

assign add_ln703_423_fu_2993_p2 = (sub_ln703_361_reg_5936 + data_22_V_read23_reg_4483_pp0_iter7_reg);

assign add_ln703_424_fu_2806_p2 = (sub_ln703_367_fu_2689_p2 + data_23_V_read24_reg_4451_pp0_iter6_reg);

assign add_ln703_425_fu_3001_p2 = (sub_ln703_369_reg_5946 + data_23_V_read24_reg_4451_pp0_iter7_reg);

assign add_ln703_426_fu_2378_p2 = (sub_ln703_244_fu_1827_p2 + data_15_V_read16_reg_4682_pp0_iter5_reg);

assign add_ln703_427_fu_2383_p2 = (add_ln703_358_fu_2123_p2 + add_ln703_426_fu_2378_p2);

assign add_ln703_428_fu_2389_p2 = (data_22_V_read23_reg_4483_pp0_iter5_reg + data_23_V_read24_reg_4451_pp0_iter5_reg);

assign add_ln703_429_fu_2825_p2 = (add_ln703_428_reg_5888 + data_21_V_read22_reg_4512_pp0_iter6_reg);

assign add_ln703_430_fu_2829_p2 = (add_ln703_429_fu_2825_p2 + add_ln703_384_reg_5701_pp0_iter6_reg);

assign add_ln703_431_fu_2834_p2 = (add_ln703_430_fu_2829_p2 + add_ln703_427_reg_5883);

assign add_ln703_432_fu_3014_p2 = (sub_ln703_374_reg_5956 + data_23_V_read24_reg_4451_pp0_iter7_reg);

assign add_ln703_433_fu_3036_p2 = (sub_ln703_379_reg_5971 + data_24_V_read25_reg_4421_pp0_iter7_reg);

assign add_ln703_434_fu_2873_p2 = (sub_ln703_380_fu_2786_p2 + data_24_V_read25_reg_4421_pp0_iter6_reg);

assign add_ln703_435_fu_2393_p2 = (data_23_V_read24_reg_4451_pp0_iter5_reg + data_24_V_read25_reg_4421_pp0_iter5_reg);

assign add_ln703_436_fu_2883_p2 = (add_ln703_435_reg_5894 + sub_ln703_365_fu_2670_p2);

assign add_ln703_437_fu_3053_p2 = (sub_ln703_385_reg_5986 + data_24_V_read25_reg_4421_pp0_iter7_reg);

assign add_ln703_438_fu_2888_p2 = (add_ln703_435_reg_5894 + sub_ln703_370_fu_2714_p2);

assign add_ln703_439_fu_3075_p2 = (sub_ln703_390_fu_3009_p2 + data_24_V_read25_reg_4421_pp0_iter7_reg);

assign add_ln703_440_fu_2908_p2 = (add_ln703_394_reg_5710_pp0_iter6_reg + sub_ln703_330_fu_2455_p2);

assign add_ln703_441_fu_2913_p2 = (add_ln703_435_reg_5894 + data_22_V_read23_reg_4483_pp0_iter6_reg);

assign add_ln703_442_fu_2917_p2 = (add_ln703_441_fu_2913_p2 + add_ln703_440_fu_2908_p2);

assign add_ln703_443_fu_3099_p2 = (sub_ln703_397_reg_6006 + data_24_V_read25_reg_4421_pp0_iter7_reg);

assign add_ln703_444_fu_2928_p2 = (sub_ln703_400_fu_2868_p2 + data_24_V_read25_reg_4421_pp0_iter6_reg);

assign add_ln703_445_fu_3122_p2 = (sub_ln703_402_reg_6016 + data_25_V_read26_reg_4391_pp0_iter7_reg);

assign add_ln703_446_fu_2397_p2 = (data_24_V_read25_reg_4421_pp0_iter5_reg + data_25_V_read26_reg_4391_pp0_iter5_reg);

assign add_ln703_447_fu_2933_p2 = (add_ln703_446_reg_5901 + sub_ln703_383_fu_2801_p2);

assign add_ln703_448_fu_3150_p2 = (sub_ln703_408_reg_6026 + data_25_V_read26_reg_4391_pp0_iter7_reg);

assign add_ln703_449_fu_3158_p2 = (sub_ln703_410_fu_3071_p2 + data_25_V_read26_reg_4391_pp0_iter7_reg);

assign add_ln703_450_fu_3168_p2 = (sub_ln703_357_reg_5926 + data_22_V_read23_reg_4483_pp0_iter7_reg);

assign add_ln703_451_fu_2943_p2 = (add_ln703_446_reg_5901 + data_23_V_read24_reg_4451_pp0_iter6_reg);

assign add_ln703_452_fu_3172_p2 = (add_ln703_451_reg_6066 + add_ln703_450_fu_3168_p2);

assign add_ln703_453_fu_3218_p2 = (sub_ln703_420_fu_3117_p2 + data_26_V_read27_reg_4365_pp0_iter7_reg);

assign add_ln703_454_fu_3232_p2 = (sub_ln703_424_fu_3140_p2 + data_26_V_read27_reg_4365_pp0_iter7_reg);

assign add_ln703_455_fu_3237_p2 = (data_25_V_read26_reg_4391_pp0_iter7_reg + data_26_V_read27_reg_4365_pp0_iter7_reg);

assign add_ln703_456_fu_3241_p2 = (add_ln703_455_fu_3237_p2 + sub_ln703_405_fu_3057_p2);

assign add_ln703_457_fu_3281_p2 = (sub_ln703_431_fu_3185_p2 + data_26_V_read27_reg_4365_pp0_iter7_reg);

assign add_ln703_458_fu_3286_p2 = (add_ln703_455_fu_3237_p2 + sub_ln703_413_fu_3084_p2);

assign add_ln703_459_fu_3292_p2 = (add_ln703_455_fu_3237_p2 + sub_ln703_415_fu_3094_p2);

assign add_ln703_460_fu_3303_p2 = (sub_ln703_433_fu_3194_p2 + data_26_V_read27_reg_4365_pp0_iter7_reg);

assign add_ln703_461_fu_3323_p2 = (sub_ln703_438_fu_3223_p2 + data_27_V_read_8_reg_4342_pp0_iter7_reg);

assign add_ln703_462_fu_2401_p2 = (data_26_V_read27_reg_4365_pp0_iter5_reg + data_27_V_read_8_reg_4342_pp0_iter5_reg);

assign add_ln703_463_fu_3328_p2 = (add_ln703_462_reg_5909_pp0_iter7_reg + sub_ln703_421_fu_3126_p2);

assign add_ln703_464_fu_3333_p2 = (sub_ln703_439_fu_3228_p2 + data_27_V_read_8_reg_4342_pp0_iter7_reg);

assign add_ln703_465_fu_3338_p2 = (add_ln703_462_reg_5909_pp0_iter7_reg + sub_ln703_422_fu_3130_p2);

assign add_ln703_466_fu_3358_p2 = (sub_ln703_407_fu_3066_p2 + data_25_V_read26_reg_4391_pp0_iter7_reg);

assign add_ln703_467_fu_3363_p2 = (add_ln703_462_reg_5909_pp0_iter7_reg + add_ln703_466_fu_3358_p2);

assign add_ln703_468_fu_3378_p2 = (sub_ln703_445_fu_3271_p2 + data_27_V_read_8_reg_4342_pp0_iter7_reg);

assign add_ln703_469_fu_3383_p2 = (sub_ln703_446_fu_3276_p2 + data_27_V_read_8_reg_4342_pp0_iter7_reg);

assign add_ln703_470_fu_3398_p2 = (sub_ln703_414_fu_3089_p2 + data_25_V_read26_reg_4391_pp0_iter7_reg);

assign add_ln703_471_fu_3403_p2 = (add_ln703_462_reg_5909_pp0_iter7_reg + add_ln703_470_fu_3398_p2);

assign add_ln703_472_fu_3413_p2 = (sub_ln703_447_fu_3298_p2 + data_27_V_read_8_reg_4342_pp0_iter7_reg);

assign add_ln703_473_fu_3423_p2 = (sub_ln703_398_fu_3026_p2 + data_24_V_read25_reg_4421_pp0_iter7_reg);

assign add_ln703_474_fu_3428_p2 = (add_ln703_462_reg_5909_pp0_iter7_reg + data_25_V_read26_reg_4391_pp0_iter7_reg);

assign add_ln703_475_fu_3432_p2 = (add_ln703_474_fu_3428_p2 + add_ln703_473_fu_3423_p2);

assign add_ln703_476_fu_3531_p2 = (add_ln703_462_reg_5909_pp0_iter8_reg + sub_ln703_434_reg_6113);

assign add_ln703_477_fu_2947_p2 = (sub_ln703_345_fu_2532_p2 + data_21_V_read22_reg_4512_pp0_iter6_reg);

assign add_ln703_478_fu_2952_p2 = (add_ln703_428_reg_5888 + add_ln703_477_fu_2947_p2);

assign add_ln703_479_fu_2957_p2 = (add_ln703_462_reg_5909 + add_ln703_446_reg_5901);

assign add_ln703_480_fu_2961_p2 = (add_ln703_479_fu_2957_p2 + add_ln703_478_fu_2952_p2);

assign add_ln703_481_fu_3443_p2 = (sub_ln703_423_fu_3135_p2 + data_26_V_read27_reg_4365_pp0_iter7_reg);

assign add_ln703_482_fu_2967_p2 = (data_27_V_read_8_reg_4342_pp0_iter6_reg + data_28_V_read_7_reg_4313_pp0_iter6_reg);

assign add_ln703_483_fu_3448_p2 = (add_ln703_482_reg_6077 + add_ln703_481_fu_3443_p2);

assign add_ln703_484_fu_3555_p2 = (sub_ln703_452_reg_6148 + data_28_V_read_7_reg_4313_pp0_iter8_reg);

assign add_ln703_485_fu_3559_p2 = (sub_ln703_453_reg_6153 + data_28_V_read_7_reg_4313_pp0_iter8_reg);

assign add_ln703_486_fu_3453_p2 = (add_ln703_482_reg_6077 + sub_ln703_442_fu_3256_p2);

assign add_ln703_487_fu_3458_p2 = (add_ln703_482_reg_6077 + sub_ln703_443_fu_3261_p2);

assign add_ln703_488_fu_3571_p2 = (sub_ln703_455_reg_6168 + data_28_V_read_7_reg_4313_pp0_iter8_reg);

assign add_ln703_489_fu_3468_p2 = (sub_ln703_430_fu_3181_p2 + data_26_V_read27_reg_4365_pp0_iter7_reg);

assign add_ln703_490_fu_3473_p2 = (add_ln703_482_reg_6077 + add_ln703_489_fu_3468_p2);

assign add_ln703_491_fu_2971_p2 = (add_ln703_446_reg_5901 + sub_ln703_395_fu_2853_p2);

assign add_ln703_492_fu_3478_p2 = (add_ln703_482_reg_6077 + data_26_V_read27_reg_4365_pp0_iter7_reg);

assign add_ln703_493_fu_3595_p2 = (add_ln703_492_reg_6223 + add_ln703_491_reg_6087_pp0_iter8_reg);

assign add_ln703_494_fu_3487_p2 = (sub_ln703_435_fu_3204_p2 + data_26_V_read27_reg_4365_pp0_iter7_reg);

assign add_ln703_495_fu_3492_p2 = (add_ln703_482_reg_6077 + add_ln703_494_fu_3487_p2);

assign add_ln703_496_fu_3497_p2 = (data_28_V_read_7_reg_4313_pp0_iter7_reg + data_29_V_read_7_reg_4279_pp0_iter7_reg);

assign add_ln703_497_fu_3501_p2 = (add_ln703_496_fu_3497_p2 + sub_ln703_449_fu_3313_p2);

assign add_ln703_498_fu_3616_p2 = (sub_ln703_460_fu_3535_p2 + data_29_V_read_7_reg_4279_pp0_iter8_reg);

assign add_ln703_499_fu_3631_p2 = (sub_ln703_464_fu_3547_p2 + data_29_V_read_7_reg_4279_pp0_iter8_reg);

assign add_ln703_500_fu_3655_p2 = (sub_ln703_466_fu_3563_p2 + data_29_V_read_7_reg_4279_pp0_iter8_reg);

assign add_ln703_501_fu_3708_p2 = (sub_ln703_475_fu_3599_p2 + data_29_V_read_7_reg_4279_pp0_iter8_reg);

assign add_ln703_502_fu_3713_p2 = (sub_ln703_476_fu_3603_p2 + data_29_V_read_7_reg_4279_pp0_iter8_reg);

assign add_ln703_503_fu_3757_p2 = (sub_ln703_483_fu_3645_p2 + data_30_V_read31_reg_4250_pp0_iter8_reg);

assign add_ln703_504_fu_3777_p2 = (sub_ln703_486_reg_6244 + data_30_V_read31_reg_4250_pp0_iter8_reg);

assign add_ln703_505_fu_3785_p2 = (sub_ln703_488_fu_3665_p2 + data_30_V_read31_reg_4250_pp0_iter8_reg);

assign add_ln703_506_fu_3795_p2 = (sub_ln703_491_reg_6254 + data_30_V_read31_reg_4250_pp0_iter8_reg);

assign add_ln703_507_fu_3799_p2 = (sub_ln703_492_fu_3679_p2 + data_30_V_read31_reg_4250_pp0_iter8_reg);

assign add_ln703_508_fu_3843_p2 = (sub_ln703_448_reg_6118 + data_28_V_read_7_reg_4313_pp0_iter8_reg);

assign add_ln703_509_fu_2976_p2 = (data_30_V_read31_reg_4250_pp0_iter6_reg + data_31_V_read32_reg_4221_pp0_iter6_reg);

assign add_ln703_510_fu_3527_p2 = (add_ln703_509_reg_6092 + data_29_V_read_7_reg_4279_pp0_iter7_reg);

assign add_ln703_511_fu_3847_p2 = (add_ln703_510_reg_6264 + add_ln703_508_fu_3843_p2);

assign add_ln703_514_fu_3862_p2 = (sub_ln703_461_reg_6208 + data_29_V_read_7_reg_4279_pp0_iter8_reg);

assign add_ln703_516_fu_2980_p2 = (sub_ln703_349_fu_2549_p2 + data_22_V_read23_reg_4483_pp0_iter6_reg);

assign add_ln703_517_fu_3871_p2 = (add_ln703_451_reg_6066_pp0_iter8_reg + add_ln703_516_reg_6103_pp0_iter8_reg);

assign add_ln703_518_fu_3875_p2 = (add_ln703_510_reg_6264 + add_ln703_492_reg_6223);

assign add_ln703_526_fu_3945_p2 = (add_ln703_462_reg_5909_pp0_iter8_reg + sub_ln703_428_reg_6108);

assign add_ln703_527_fu_3949_p2 = (add_ln703_509_reg_6092_pp0_iter8_reg + add_ln703_496_reg_6234);

assign add_ln703_fu_280_p2 = (data_0_V_read_int_reg + data_1_V_read_int_reg);

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_state10_pp0_stage0_iter9 = ~(1'b1 == 1'b1);

assign ap_block_state1_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter4 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage0_iter5 = ~(1'b1 == 1'b1);

assign ap_block_state7_pp0_stage0_iter6 = ~(1'b1 == 1'b1);

assign ap_block_state8_pp0_stage0_iter7 = ~(1'b1 == 1'b1);

assign ap_block_state9_pp0_stage0_iter8 = ~(1'b1 == 1'b1);

assign sub_ln703_100_fu_617_p2 = (add_ln703_210_reg_5143_pp0_iter3_reg - data_5_V_read_8_reg_4969_pp0_iter3_reg);

assign sub_ln703_101_fu_621_p2 = (add_ln703_213_reg_5189 - data_5_V_read_8_reg_4969_pp0_iter3_reg);

assign sub_ln703_102_fu_625_p2 = (sub_ln703_89_reg_5166 - data_5_V_read_8_reg_4969_pp0_iter3_reg);

assign sub_ln703_103_fu_629_p2 = (add_ln703_214_reg_5194 - data_5_V_read_8_reg_4969_pp0_iter3_reg);

assign sub_ln703_104_fu_633_p2 = (add_ln703_211_reg_5184 - data_5_V_read_8_reg_4969_pp0_iter3_reg);

assign sub_ln703_105_fu_489_p2 = (sub_ln703_92_fu_437_p2 - data_5_V_read_8_reg_4969_pp0_iter2_reg);

assign sub_ln703_106_fu_494_p2 = (add_ln703_212_fu_425_p2 - data_5_V_read_8_reg_4969_pp0_iter2_reg);

assign sub_ln703_107_fu_637_p2 = (sub_ln703_93_reg_5200 - data_5_V_read_8_reg_4969_pp0_iter3_reg);

assign sub_ln703_108_fu_641_p2 = (sub_ln703_94_reg_5205 - data_6_V_read_8_reg_4944_pp0_iter3_reg);

assign sub_ln703_109_fu_649_p2 = (add_ln703_215_fu_605_p2 - data_6_V_read_8_reg_4944_pp0_iter3_reg);

assign sub_ln703_110_fu_654_p2 = (add_ln703_216_reg_5215 - data_6_V_read_8_reg_4944_pp0_iter3_reg);

assign sub_ln703_111_fu_658_p2 = (sub_ln703_97_fu_609_p2 - data_6_V_read_8_reg_4944_pp0_iter3_reg);

assign sub_ln703_112_fu_528_p2 = (add_ln703_217_fu_470_p2 - data_6_V_read_8_reg_4944_pp0_iter2_reg);

assign sub_ln703_113_fu_533_p2 = (add_ln703_218_fu_474_p2 - data_6_V_read_8_reg_4944_pp0_iter2_reg);

assign sub_ln703_114_fu_549_p2 = (add_ln703_219_fu_479_p2 - data_6_V_read_8_reg_4944_pp0_iter2_reg);

assign sub_ln703_115_fu_678_p2 = (sub_ln703_103_fu_629_p2 - data_6_V_read_8_reg_4944_pp0_iter3_reg);

assign sub_ln703_116_fu_683_p2 = (add_ln703_220_reg_5221 - data_6_V_read_8_reg_4944_pp0_iter3_reg);

assign sub_ln703_117_fu_554_p2 = (sub_ln703_106_fu_494_p2 - data_6_V_read_8_reg_4944_pp0_iter2_reg);

assign sub_ln703_118_fu_559_p2 = (add_ln703_221_fu_499_p2 - data_6_V_read_8_reg_4944_pp0_iter2_reg);

assign sub_ln703_119_fu_687_p2 = (add_ln703_223_reg_5231 - data_7_V_read_8_reg_4916_pp0_iter3_reg);

assign sub_ln703_120_fu_691_p2 = (sub_ln703_108_fu_641_p2 - data_7_V_read_8_reg_4916_pp0_iter3_reg);

assign sub_ln703_121_fu_696_p2 = (add_ln703_224_fu_645_p2 - data_7_V_read_8_reg_4916_pp0_iter3_reg);

assign sub_ln703_122_fu_705_p2 = (sub_ln703_110_fu_654_p2 - data_7_V_read_8_reg_4916_pp0_iter3_reg);

assign sub_ln703_123_fu_719_p2 = (add_ln703_225_reg_5237 - data_7_V_read_8_reg_4916_pp0_iter3_reg);

assign sub_ln703_124_fu_723_p2 = (add_ln703_227_reg_5242 - data_7_V_read_8_reg_4916_pp0_iter3_reg);

assign sub_ln703_125_fu_727_p2 = (add_ln703_228_fu_663_p2 - data_7_V_read_8_reg_4916_pp0_iter3_reg);

assign sub_ln703_126_fu_574_p2 = (sub_ln703_112_fu_528_p2 - data_7_V_read_8_reg_4916_pp0_iter2_reg);

assign sub_ln703_127_fu_732_p2 = (sub_ln703_113_reg_5247 - data_7_V_read_8_reg_4916_pp0_iter3_reg);

assign sub_ln703_128_fu_736_p2 = (add_ln703_229_fu_668_p2 - data_7_V_read_8_reg_4916_pp0_iter3_reg);

assign sub_ln703_129_fu_579_p2 = (add_ln703_231_fu_543_p2 - data_7_V_read_8_reg_4916_pp0_iter2_reg);

assign sub_ln703_130_fu_741_p2 = (sub_ln703_114_reg_5253 - data_7_V_read_8_reg_4916_pp0_iter3_reg);

assign sub_ln703_131_fu_745_p2 = (add_ln703_232_fu_673_p2 - data_7_V_read_8_reg_4916_pp0_iter3_reg);

assign sub_ln703_132_fu_760_p2 = (sub_ln703_116_fu_683_p2 - data_7_V_read_8_reg_4916_pp0_iter3_reg);

assign sub_ln703_133_fu_584_p2 = (sub_ln703_118_fu_559_p2 - data_7_V_read_8_reg_4916_pp0_iter2_reg);

assign sub_ln703_134_fu_792_p2 = (add_ln703_234_reg_5264 - data_8_V_read_7_reg_4887_pp0_iter3_reg);

assign sub_ln703_135_fu_796_p2 = (sub_ln703_121_fu_696_p2 - data_8_V_read_7_reg_4887_pp0_iter3_reg);

assign sub_ln703_136_fu_806_p2 = (add_ln703_235_fu_701_p2 - data_8_V_read_7_reg_4887_pp0_iter3_reg);

assign sub_ln703_137_fu_811_p2 = (sub_ln703_122_fu_705_p2 - data_8_V_read_7_reg_4887_pp0_iter3_reg);

assign sub_ln703_138_fu_816_p2 = (add_ln703_236_fu_710_p2 - data_8_V_read_7_reg_4887_pp0_iter3_reg);

assign sub_ln703_139_fu_821_p2 = (add_ln703_237_fu_715_p2 - data_8_V_read_7_reg_4887_pp0_iter3_reg);

assign sub_ln703_140_fu_826_p2 = (add_ln703_238_reg_5269 - data_8_V_read_7_reg_4887_pp0_iter3_reg);

assign sub_ln703_141_fu_835_p2 = (sub_ln703_125_fu_727_p2 - data_8_V_read_7_reg_4887_pp0_iter3_reg);

assign sub_ln703_142_fu_840_p2 = (sub_ln703_126_reg_5274 - data_8_V_read_7_reg_4887_pp0_iter3_reg);

assign sub_ln703_143_fu_844_p2 = (sub_ln703_128_fu_736_p2 - data_8_V_read_7_reg_4887_pp0_iter3_reg);

assign sub_ln703_144_fu_858_p2 = (add_ln703_239_fu_750_p2 - data_8_V_read_7_reg_4887_pp0_iter3_reg);

assign sub_ln703_145_fu_863_p2 = (add_ln703_240_fu_755_p2 - data_8_V_read_7_reg_4887_pp0_iter3_reg);

assign sub_ln703_146_fu_868_p2 = (sub_ln703_132_fu_760_p2 - data_8_V_read_7_reg_4887_pp0_iter3_reg);

assign sub_ln703_147_fu_882_p2 = (add_ln703_241_fu_765_p2 - data_8_V_read_7_reg_4887_pp0_iter3_reg);

assign sub_ln703_148_fu_896_p2 = (add_ln703_242_fu_769_p2 - data_8_V_read_7_reg_4887_pp0_iter3_reg);

assign sub_ln703_149_fu_901_p2 = (add_ln703_244_fu_778_p2 - data_8_V_read_7_reg_4887_pp0_iter3_reg);

assign sub_ln703_150_fu_906_p2 = (add_ln703_245_fu_783_p2 - data_8_V_read_7_reg_4887_pp0_iter3_reg);

assign sub_ln703_151_fu_911_p2 = (sub_ln703_133_reg_5284 - data_8_V_read_7_reg_4887_pp0_iter3_reg);

assign sub_ln703_152_fu_1202_p2 = (add_ln703_246_reg_5320 - data_9_V_read_7_reg_4859_pp0_iter4_reg);

assign sub_ln703_153_fu_915_p2 = (sub_ln703_134_fu_792_p2 - data_9_V_read_7_reg_4859_pp0_iter3_reg);

assign sub_ln703_154_fu_920_p2 = (add_ln703_248_fu_801_p2 - data_9_V_read_7_reg_4859_pp0_iter3_reg);

assign sub_ln703_155_fu_1206_p2 = (sub_ln703_138_reg_5325 - data_9_V_read_7_reg_4859_pp0_iter4_reg);

assign sub_ln703_156_fu_930_p2 = (sub_ln703_140_fu_826_p2 - data_9_V_read_7_reg_4859_pp0_iter3_reg);

assign sub_ln703_157_fu_935_p2 = (add_ln703_249_fu_830_p2 - data_9_V_read_7_reg_4859_pp0_iter3_reg);

assign sub_ln703_158_fu_1210_p2 = (sub_ln703_141_reg_5330 - data_9_V_read_7_reg_4859_pp0_iter4_reg);

assign sub_ln703_159_fu_945_p2 = (sub_ln703_142_fu_840_p2 - data_9_V_read_7_reg_4859_pp0_iter3_reg);

assign sub_ln703_160_fu_1214_p2 = (sub_ln703_143_reg_5335 - data_9_V_read_7_reg_4859_pp0_iter4_reg);

assign sub_ln703_161_fu_960_p2 = (add_ln703_252_fu_853_p2 - data_9_V_read_7_reg_4859_pp0_iter3_reg);

assign sub_ln703_162_fu_980_p2 = (sub_ln703_146_fu_868_p2 - data_9_V_read_7_reg_4859_pp0_iter3_reg);

assign sub_ln703_163_fu_985_p2 = (add_ln703_254_fu_877_p2 - data_9_V_read_7_reg_4859_pp0_iter3_reg);

assign sub_ln703_164_fu_990_p2 = (sub_ln703_147_fu_882_p2 - data_9_V_read_7_reg_4859_pp0_iter3_reg);

assign sub_ln703_165_fu_995_p2 = (add_ln703_256_fu_891_p2 - data_9_V_read_7_reg_4859_pp0_iter3_reg);

assign sub_ln703_166_fu_1000_p2 = (sub_ln703_148_fu_896_p2 - data_9_V_read_7_reg_4859_pp0_iter3_reg);

assign sub_ln703_167_fu_1218_p2 = (sub_ln703_149_reg_5350 - data_9_V_read_7_reg_4859_pp0_iter4_reg);

assign sub_ln703_168_fu_1005_p2 = (sub_ln703_151_fu_911_p2 - data_9_V_read_7_reg_4859_pp0_iter3_reg);

assign sub_ln703_169_fu_1222_p2 = (sub_ln703_152_fu_1202_p2 - data_10_V_read11_reg_4832_pp0_iter4_reg);

assign sub_ln703_170_fu_1227_p2 = (sub_ln703_155_fu_1206_p2 - data_10_V_read11_reg_4832_pp0_iter4_reg);

assign sub_ln703_171_fu_1015_p2 = (add_ln703_257_fu_925_p2 - data_10_V_read11_reg_4832_pp0_iter3_reg);

assign sub_ln703_172_fu_1020_p2 = (sub_ln703_156_fu_930_p2 - data_10_V_read11_reg_4832_pp0_iter3_reg);

assign sub_ln703_173_fu_1025_p2 = (sub_ln703_157_fu_935_p2 - data_10_V_read11_reg_4832_pp0_iter3_reg);

assign sub_ln703_174_fu_1030_p2 = (add_ln703_259_fu_940_p2 - data_10_V_read11_reg_4832_pp0_iter3_reg);

assign sub_ln703_175_fu_1035_p2 = (sub_ln703_159_fu_945_p2 - data_10_V_read11_reg_4832_pp0_iter3_reg);

assign sub_ln703_176_fu_1040_p2 = (add_ln703_260_fu_950_p2 - data_10_V_read11_reg_4832_pp0_iter3_reg);

assign sub_ln703_177_fu_1237_p2 = (sub_ln703_160_fu_1214_p2 - data_10_V_read11_reg_4832_pp0_iter4_reg);

assign sub_ln703_178_fu_1242_p2 = (add_ln703_261_reg_5360 - data_10_V_read11_reg_4832_pp0_iter4_reg);

assign sub_ln703_179_fu_1246_p2 = (sub_ln703_161_reg_5365 - data_10_V_read11_reg_4832_pp0_iter4_reg);

assign sub_ln703_180_fu_1045_p2 = (add_ln703_264_fu_974_p2 - data_10_V_read11_reg_4832_pp0_iter3_reg);

assign sub_ln703_181_fu_1050_p2 = (sub_ln703_163_fu_985_p2 - data_10_V_read11_reg_4832_pp0_iter3_reg);

assign sub_ln703_182_fu_1060_p2 = (sub_ln703_165_fu_995_p2 - data_10_V_read11_reg_4832_pp0_iter3_reg);

assign sub_ln703_183_fu_1250_p2 = (sub_ln703_167_fu_1218_p2 - data_10_V_read11_reg_4832_pp0_iter4_reg);

assign sub_ln703_184_fu_1075_p2 = (sub_ln703_168_fu_1005_p2 - data_10_V_read11_reg_4832_pp0_iter3_reg);

assign sub_ln703_185_fu_1095_p2 = (add_ln703_265_fu_1010_p2 - data_11_V_read12_reg_4808_pp0_iter3_reg);

assign sub_ln703_186_fu_1272_p2 = (sub_ln703_170_fu_1227_p2 - data_11_V_read12_reg_4808_pp0_iter4_reg);

assign sub_ln703_187_fu_1110_p2 = (sub_ln703_172_fu_1020_p2 - data_11_V_read12_reg_4808_pp0_iter3_reg);

assign sub_ln703_188_fu_1277_p2 = (sub_ln703_173_reg_5385 - data_11_V_read12_reg_4808_pp0_iter4_reg);

assign sub_ln703_189_fu_1115_p2 = (sub_ln703_174_fu_1030_p2 - data_11_V_read12_reg_4808_pp0_iter3_reg);

assign sub_ln703_190_fu_1281_p2 = (add_ln703_266_fu_1232_p2 - data_11_V_read12_reg_4808_pp0_iter4_reg);

assign sub_ln703_191_fu_1120_p2 = (sub_ln703_175_fu_1035_p2 - data_11_V_read12_reg_4808_pp0_iter3_reg);

assign sub_ln703_192_fu_1286_p2 = (sub_ln703_177_fu_1237_p2 - data_11_V_read12_reg_4808_pp0_iter4_reg);

assign sub_ln703_193_fu_1291_p2 = (sub_ln703_179_fu_1246_p2 - data_11_V_read12_reg_4808_pp0_iter4_reg);

assign sub_ln703_194_fu_1309_p2 = (sub_ln703_181_reg_5400 - data_11_V_read12_reg_4808_pp0_iter4_reg);

assign sub_ln703_195_fu_1313_p2 = (add_ln703_267_reg_5405 - data_11_V_read12_reg_4808_pp0_iter4_reg);

assign sub_ln703_196_fu_1317_p2 = (sub_ln703_182_reg_5410 - data_11_V_read12_reg_4808_pp0_iter4_reg);

assign sub_ln703_197_fu_1321_p2 = (sub_ln703_183_fu_1250_p2 - data_11_V_read12_reg_4808_pp0_iter4_reg);

assign sub_ln703_198_fu_1146_p2 = (add_ln703_269_fu_1069_p2 - data_11_V_read12_reg_4808_pp0_iter3_reg);

assign sub_ln703_199_fu_1151_p2 = (sub_ln703_184_fu_1075_p2 - data_11_V_read12_reg_4808_pp0_iter3_reg);

assign sub_ln703_200_fu_1326_p2 = (add_ln703_270_fu_1255_p2 - data_12_V_read13_reg_4778_pp0_iter4_reg);

assign sub_ln703_201_fu_1331_p2 = (add_ln703_274_reg_5420 - data_12_V_read13_reg_4778_pp0_iter4_reg);

assign sub_ln703_202_fu_1335_p2 = (sub_ln703_185_reg_5425 - data_12_V_read13_reg_4778_pp0_iter4_reg);

assign sub_ln703_203_fu_1339_p2 = (add_ln703_275_fu_1260_p2 - data_12_V_read13_reg_4778_pp0_iter4_reg);

assign sub_ln703_204_fu_1344_p2 = (add_ln703_277_fu_1264_p2 - data_12_V_read13_reg_4778_pp0_iter4_reg);

assign sub_ln703_205_fu_1349_p2 = (add_ln703_279_fu_1268_p2 - data_12_V_read13_reg_4778_pp0_iter4_reg);

assign sub_ln703_206_fu_1363_p2 = (sub_ln703_187_reg_5440 - data_12_V_read13_reg_4778_pp0_iter4_reg);

assign sub_ln703_207_fu_1384_p2 = (sub_ln703_192_fu_1286_p2 - data_12_V_read13_reg_4778_pp0_iter4_reg);

assign sub_ln703_208_fu_1389_p2 = (add_ln703_281_reg_5455 - data_12_V_read13_reg_4778_pp0_iter4_reg);

assign sub_ln703_209_fu_1393_p2 = (add_ln703_283_reg_5460 - data_12_V_read13_reg_4778_pp0_iter4_reg);

assign sub_ln703_210_fu_1402_p2 = (sub_ln703_193_fu_1291_p2 - data_12_V_read13_reg_4778_pp0_iter4_reg);

assign sub_ln703_211_fu_1407_p2 = (add_ln703_285_fu_1300_p2 - data_12_V_read13_reg_4778_pp0_iter4_reg);

assign sub_ln703_212_fu_1412_p2 = (add_ln703_286_fu_1305_p2 - data_12_V_read13_reg_4778_pp0_iter4_reg);

assign sub_ln703_213_fu_1417_p2 = (sub_ln703_194_fu_1309_p2 - data_12_V_read13_reg_4778_pp0_iter4_reg);

assign sub_ln703_214_fu_1422_p2 = (sub_ln703_195_fu_1313_p2 - data_12_V_read13_reg_4778_pp0_iter4_reg);

assign sub_ln703_215_fu_1441_p2 = (sub_ln703_197_fu_1321_p2 - data_12_V_read13_reg_4778_pp0_iter4_reg);

assign sub_ln703_216_fu_1446_p2 = (sub_ln703_198_reg_5465 - data_12_V_read13_reg_4778_pp0_iter4_reg);

assign sub_ln703_217_fu_1450_p2 = (sub_ln703_199_reg_5470 - data_12_V_read13_reg_4778_pp0_iter4_reg);

assign sub_ln703_218_fu_1784_p2 = (sub_ln703_200_reg_5515 - data_13_V_read14_reg_4745_pp0_iter5_reg);

assign sub_ln703_219_fu_1788_p2 = (sub_ln703_203_reg_5520 - data_13_V_read14_reg_4745_pp0_iter5_reg);

assign sub_ln703_220_fu_1459_p2 = (sub_ln703_204_fu_1344_p2 - data_13_V_read14_reg_4745_pp0_iter4_reg);

assign sub_ln703_221_fu_1792_p2 = (add_ln703_287_reg_5525 - data_13_V_read14_reg_4745_pp0_iter5_reg);

assign sub_ln703_222_fu_1469_p2 = (add_ln703_289_fu_1359_p2 - data_13_V_read14_reg_4745_pp0_iter4_reg);

assign sub_ln703_223_fu_1479_p2 = (add_ln703_290_fu_1367_p2 - data_13_V_read14_reg_4745_pp0_iter4_reg);

assign sub_ln703_224_fu_1796_p2 = (add_ln703_291_reg_5530 - data_13_V_read14_reg_4745_pp0_iter5_reg);

assign sub_ln703_225_fu_1484_p2 = (add_ln703_292_fu_1376_p2 - data_13_V_read14_reg_4745_pp0_iter4_reg);

assign sub_ln703_226_fu_1489_p2 = (add_ln703_293_fu_1380_p2 - data_13_V_read14_reg_4745_pp0_iter4_reg);

assign sub_ln703_227_fu_1800_p2 = (sub_ln703_207_reg_5535 - data_13_V_read14_reg_4745_pp0_iter5_reg);

assign sub_ln703_228_fu_1499_p2 = (add_ln703_294_fu_1397_p2 - data_13_V_read14_reg_4745_pp0_iter4_reg);

assign sub_ln703_229_fu_1518_p2 = (sub_ln703_211_fu_1407_p2 - data_13_V_read14_reg_4745_pp0_iter4_reg);

assign sub_ln703_230_fu_1804_p2 = (sub_ln703_212_reg_5540 - data_13_V_read14_reg_4745_pp0_iter5_reg);

assign sub_ln703_231_fu_1537_p2 = (add_ln703_295_fu_1427_p2 - data_13_V_read14_reg_4745_pp0_iter4_reg);

assign sub_ln703_232_fu_1542_p2 = (add_ln703_297_fu_1436_p2 - data_13_V_read14_reg_4745_pp0_iter4_reg);

assign sub_ln703_233_fu_1808_p2 = (sub_ln703_215_reg_5545 - data_13_V_read14_reg_4745_pp0_iter5_reg);

assign sub_ln703_234_fu_1547_p2 = (sub_ln703_217_fu_1450_p2 - data_13_V_read14_reg_4745_pp0_iter4_reg);

assign sub_ln703_235_fu_1812_p2 = (sub_ln703_218_fu_1784_p2 - data_14_V_read15_reg_4714_pp0_iter5_reg);

assign sub_ln703_236_fu_1557_p2 = (add_ln703_298_fu_1454_p2 - data_14_V_read15_reg_4714_pp0_iter4_reg);

assign sub_ln703_237_fu_1571_p2 = (sub_ln703_220_fu_1459_p2 - data_14_V_read15_reg_4714_pp0_iter4_reg);

assign sub_ln703_238_fu_1576_p2 = (add_ln703_299_fu_1464_p2 - data_14_V_read15_reg_4714_pp0_iter4_reg);

assign sub_ln703_239_fu_1817_p2 = (sub_ln703_221_fu_1792_p2 - data_14_V_read15_reg_4714_pp0_iter5_reg);

assign sub_ln703_240_fu_1581_p2 = (sub_ln703_222_fu_1469_p2 - data_14_V_read15_reg_4714_pp0_iter4_reg);

assign sub_ln703_241_fu_1586_p2 = (add_ln703_300_fu_1474_p2 - data_14_V_read15_reg_4714_pp0_iter4_reg);

assign sub_ln703_242_fu_1596_p2 = (sub_ln703_225_fu_1484_p2 - data_14_V_read15_reg_4714_pp0_iter4_reg);

assign sub_ln703_243_fu_1601_p2 = (sub_ln703_226_fu_1489_p2 - data_14_V_read15_reg_4714_pp0_iter4_reg);

assign sub_ln703_244_fu_1827_p2 = (sub_ln703_227_fu_1800_p2 - data_14_V_read15_reg_4714_pp0_iter5_reg);

assign sub_ln703_245_fu_1832_p2 = (add_ln703_301_reg_5550 - data_14_V_read15_reg_4714_pp0_iter5_reg);

assign sub_ln703_246_fu_1193_p2 = (add_ln703_306_fu_1173_p2 - data_14_V_read15_reg_4714_pp0_iter3_reg);

assign sub_ln703_247_fu_1836_p2 = (add_ln703_307_reg_5555 - data_14_V_read15_reg_4714_pp0_iter5_reg);

assign sub_ln703_248_fu_1606_p2 = (add_ln703_310_fu_1513_p2 - data_14_V_read15_reg_4714_pp0_iter4_reg);

assign sub_ln703_249_fu_1840_p2 = (sub_ln703_229_reg_5560 - data_14_V_read15_reg_4714_pp0_iter5_reg);

assign sub_ln703_250_fu_1844_p2 = (sub_ln703_230_fu_1804_p2 - data_14_V_read15_reg_4714_pp0_iter5_reg);

assign sub_ln703_251_fu_1611_p2 = (add_ln703_312_fu_1527_p2 - data_14_V_read15_reg_4714_pp0_iter4_reg);

assign sub_ln703_252_fu_1616_p2 = (add_ln703_313_fu_1532_p2 - data_14_V_read15_reg_4714_pp0_iter4_reg);

assign sub_ln703_253_fu_1621_p2 = (sub_ln703_231_fu_1537_p2 - data_14_V_read15_reg_4714_pp0_iter4_reg);

assign sub_ln703_254_fu_1626_p2 = (sub_ln703_232_fu_1542_p2 - data_14_V_read15_reg_4714_pp0_iter4_reg);

assign sub_ln703_255_fu_1849_p2 = (sub_ln703_233_fu_1808_p2 - data_14_V_read15_reg_4714_pp0_iter5_reg);

assign sub_ln703_256_fu_1631_p2 = (add_ln703_315_fu_1552_p2 - data_15_V_read16_reg_4682_pp0_iter4_reg);

assign sub_ln703_257_fu_1641_p2 = (add_ln703_318_fu_1566_p2 - data_15_V_read16_reg_4682_pp0_iter4_reg);

assign sub_ln703_258_fu_1854_p2 = (sub_ln703_237_reg_5565 - data_15_V_read16_reg_4682_pp0_iter5_reg);

assign sub_ln703_259_fu_1858_p2 = (sub_ln703_238_reg_5570 - data_15_V_read16_reg_4682_pp0_iter5_reg);

assign sub_ln703_260_fu_1862_p2 = (sub_ln703_239_fu_1817_p2 - data_15_V_read16_reg_4682_pp0_iter5_reg);

assign sub_ln703_261_fu_1646_p2 = (sub_ln703_240_fu_1581_p2 - data_15_V_read16_reg_4682_pp0_iter4_reg);

assign sub_ln703_262_fu_1651_p2 = (sub_ln703_241_fu_1586_p2 - data_15_V_read16_reg_4682_pp0_iter4_reg);

assign sub_ln703_263_fu_1671_p2 = (add_ln703_319_fu_1591_p2 - data_15_V_read16_reg_4682_pp0_iter4_reg);

assign sub_ln703_264_fu_1867_p2 = (add_ln703_320_fu_1822_p2 - data_15_V_read16_reg_4682_pp0_iter5_reg);

assign sub_ln703_265_fu_1676_p2 = (sub_ln703_242_fu_1596_p2 - data_15_V_read16_reg_4682_pp0_iter4_reg);

assign sub_ln703_266_fu_1681_p2 = (sub_ln703_243_fu_1601_p2 - data_15_V_read16_reg_4682_pp0_iter4_reg);

assign sub_ln703_267_fu_1872_p2 = (sub_ln703_245_fu_1832_p2 - data_15_V_read16_reg_4682_pp0_iter5_reg);

assign sub_ln703_268_fu_1691_p2 = (sub_ln703_246_reg_5501 - data_15_V_read16_reg_4682_pp0_iter4_reg);

assign sub_ln703_269_fu_1877_p2 = (sub_ln703_247_fu_1836_p2 - data_15_V_read16_reg_4682_pp0_iter5_reg);

assign sub_ln703_270_fu_1695_p2 = (sub_ln703_248_fu_1606_p2 - data_15_V_read16_reg_4682_pp0_iter4_reg);

assign sub_ln703_271_fu_1882_p2 = (sub_ln703_249_fu_1840_p2 - data_15_V_read16_reg_4682_pp0_iter5_reg);

assign sub_ln703_272_fu_1700_p2 = (sub_ln703_251_fu_1611_p2 - data_15_V_read16_reg_4682_pp0_iter4_reg);

assign sub_ln703_273_fu_1896_p2 = (sub_ln703_253_reg_5580 - data_15_V_read16_reg_4682_pp0_iter5_reg);

assign sub_ln703_274_fu_1904_p2 = (sub_ln703_255_fu_1849_p2 - data_15_V_read16_reg_4682_pp0_iter5_reg);

assign sub_ln703_275_fu_1909_p2 = (add_ln703_321_reg_5590 - data_16_V_read17_reg_4650_pp0_iter5_reg);

assign sub_ln703_276_fu_1918_p2 = (sub_ln703_260_fu_1862_p2 - data_16_V_read17_reg_4650_pp0_iter5_reg);

assign sub_ln703_277_fu_1927_p2 = (sub_ln703_262_reg_5605 - data_16_V_read17_reg_4650_pp0_iter5_reg);

assign sub_ln703_278_fu_1735_p2 = (add_ln703_325_fu_1665_p2 - data_16_V_read17_reg_4650_pp0_iter4_reg);

assign sub_ln703_279_fu_1931_p2 = (sub_ln703_263_reg_5610 - data_16_V_read17_reg_4650_pp0_iter5_reg);

assign sub_ln703_280_fu_1935_p2 = (sub_ln703_265_reg_5615 - data_16_V_read17_reg_4650_pp0_iter5_reg);

assign sub_ln703_281_fu_1957_p2 = (add_ln703_326_reg_5625 - data_16_V_read17_reg_4650_pp0_iter5_reg);

assign sub_ln703_282_fu_1961_p2 = (sub_ln703_269_fu_1877_p2 - data_16_V_read17_reg_4650_pp0_iter5_reg);

assign sub_ln703_283_fu_1975_p2 = (add_ln703_327_fu_1887_p2 - data_16_V_read17_reg_4650_pp0_iter5_reg);

assign sub_ln703_284_fu_1980_p2 = (sub_ln703_272_reg_5635 - data_16_V_read17_reg_4650_pp0_iter5_reg);

assign sub_ln703_285_fu_1984_p2 = (add_ln703_328_fu_1892_p2 - data_16_V_read17_reg_4650_pp0_iter5_reg);

assign sub_ln703_286_fu_1989_p2 = (add_ln703_330_reg_5640 - data_16_V_read17_reg_4650_pp0_iter5_reg);

assign sub_ln703_287_fu_1998_p2 = (add_ln703_331_fu_1900_p2 - data_16_V_read17_reg_4650_pp0_iter5_reg);

assign sub_ln703_288_fu_2003_p2 = (sub_ln703_274_fu_1904_p2 - data_16_V_read17_reg_4650_pp0_iter5_reg);

assign sub_ln703_289_fu_1750_p2 = (add_ln703_333_fu_1720_p2 - data_16_V_read17_reg_4650_pp0_iter4_reg);

assign sub_ln703_290_fu_1755_p2 = (add_ln703_334_fu_1725_p2 - data_16_V_read17_reg_4650_pp0_iter4_reg);

assign sub_ln703_291_fu_2008_p2 = (add_ln703_335_reg_5645 - data_17_V_read_8_reg_4621_pp0_iter5_reg);

assign sub_ln703_292_fu_2012_p2 = (sub_ln703_275_fu_1909_p2 - data_17_V_read_8_reg_4621_pp0_iter5_reg);

assign sub_ln703_293_fu_2036_p2 = (add_ln703_336_fu_1913_p2 - data_17_V_read_8_reg_4621_pp0_iter5_reg);

assign sub_ln703_294_fu_2405_p2 = (sub_ln703_276_reg_5728 - data_17_V_read_8_reg_4621_pp0_iter6_reg);

assign sub_ln703_295_fu_2041_p2 = (add_ln703_337_fu_1923_p2 - data_17_V_read_8_reg_4621_pp0_iter5_reg);

assign sub_ln703_296_fu_2046_p2 = (sub_ln703_277_fu_1927_p2 - data_17_V_read_8_reg_4621_pp0_iter5_reg);

assign sub_ln703_297_fu_2055_p2 = (sub_ln703_279_fu_1931_p2 - data_17_V_read_8_reg_4621_pp0_iter5_reg);

assign sub_ln703_298_fu_2065_p2 = (sub_ln703_280_fu_1935_p2 - data_17_V_read_8_reg_4621_pp0_iter5_reg);

assign sub_ln703_299_fu_2070_p2 = (add_ln703_338_fu_1939_p2 - data_17_V_read_8_reg_4621_pp0_iter5_reg);

assign sub_ln703_300_fu_2075_p2 = (add_ln703_342_fu_1952_p2 - data_17_V_read_8_reg_4621_pp0_iter5_reg);

assign sub_ln703_301_fu_2085_p2 = (add_ln703_343_reg_5660 - data_17_V_read_8_reg_4621_pp0_iter5_reg);

assign sub_ln703_302_fu_2089_p2 = (sub_ln703_282_fu_1961_p2 - data_17_V_read_8_reg_4621_pp0_iter5_reg);

assign sub_ln703_303_fu_2094_p2 = (add_ln703_344_fu_1966_p2 - data_17_V_read_8_reg_4621_pp0_iter5_reg);

assign sub_ln703_304_fu_2099_p2 = (add_ln703_345_fu_1970_p2 - data_17_V_read_8_reg_4621_pp0_iter5_reg);

assign sub_ln703_305_fu_2104_p2 = (sub_ln703_286_fu_1989_p2 - data_17_V_read_8_reg_4621_pp0_iter5_reg);

assign sub_ln703_306_fu_2109_p2 = (add_ln703_346_fu_1993_p2 - data_17_V_read_8_reg_4621_pp0_iter5_reg);

assign sub_ln703_307_fu_2133_p2 = (sub_ln703_291_fu_2008_p2 - data_18_V_read_7_reg_4594_pp0_iter5_reg);

assign sub_ln703_308_fu_2143_p2 = (add_ln703_348_fu_2017_p2 - data_18_V_read_7_reg_4594_pp0_iter5_reg);

assign sub_ln703_309_fu_2148_p2 = (add_ln703_351_fu_2030_p2 - data_18_V_read_7_reg_4594_pp0_iter5_reg);

assign sub_ln703_310_fu_2168_p2 = (sub_ln703_296_fu_2046_p2 - data_18_V_read_7_reg_4594_pp0_iter5_reg);

assign sub_ln703_311_fu_2173_p2 = (add_ln703_352_fu_2051_p2 - data_18_V_read_7_reg_4594_pp0_iter5_reg);

assign sub_ln703_312_fu_2409_p2 = (add_ln703_353_reg_5743 - data_18_V_read_7_reg_4594_pp0_iter6_reg);

assign sub_ln703_313_fu_2413_p2 = (sub_ln703_300_reg_5748 - data_18_V_read_7_reg_4594_pp0_iter6_reg);

assign sub_ln703_314_fu_2417_p2 = (add_ln703_354_reg_5753 - data_18_V_read_7_reg_4594_pp0_iter6_reg);

assign sub_ln703_315_fu_2188_p2 = (sub_ln703_301_fu_2085_p2 - data_18_V_read_7_reg_4594_pp0_iter5_reg);

assign sub_ln703_316_fu_2421_p2 = (sub_ln703_302_reg_5758 - data_18_V_read_7_reg_4594_pp0_iter6_reg);

assign sub_ln703_317_fu_2425_p2 = (sub_ln703_304_reg_5763 - data_18_V_read_7_reg_4594_pp0_iter6_reg);

assign sub_ln703_318_fu_2203_p2 = (sub_ln703_306_fu_2109_p2 - data_18_V_read_7_reg_4594_pp0_iter5_reg);

assign sub_ln703_319_fu_2208_p2 = (add_ln703_355_fu_2114_p2 - data_18_V_read_7_reg_4594_pp0_iter5_reg);

assign sub_ln703_320_fu_2433_p2 = (add_ln703_359_reg_5768 - data_19_V_read_7_reg_4567_pp0_iter6_reg);

assign sub_ln703_321_fu_2218_p2 = (add_ln703_360_fu_2138_p2 - data_19_V_read_7_reg_4567_pp0_iter5_reg);

assign sub_ln703_322_fu_2223_p2 = (sub_ln703_308_fu_2143_p2 - data_19_V_read_7_reg_4567_pp0_iter5_reg);

assign sub_ln703_323_fu_2233_p2 = (add_ln703_362_fu_2158_p2 - data_19_V_read_7_reg_4567_pp0_iter5_reg);

assign sub_ln703_324_fu_2238_p2 = (add_ln703_363_fu_2163_p2 - data_19_V_read_7_reg_4567_pp0_iter5_reg);

assign sub_ln703_325_fu_2243_p2 = (sub_ln703_310_fu_2168_p2 - data_19_V_read_7_reg_4567_pp0_iter5_reg);

assign sub_ln703_326_fu_2441_p2 = (sub_ln703_311_reg_5778 - data_19_V_read_7_reg_4567_pp0_iter6_reg);

assign sub_ln703_327_fu_2248_p2 = (add_ln703_364_fu_2178_p2 - data_19_V_read_7_reg_4567_pp0_iter5_reg);

assign sub_ln703_328_fu_2253_p2 = (add_ln703_365_fu_2183_p2 - data_19_V_read_7_reg_4567_pp0_iter5_reg);

assign sub_ln703_329_fu_2450_p2 = (sub_ln703_314_fu_2417_p2 - data_19_V_read_7_reg_4567_pp0_iter6_reg);

assign sub_ln703_330_fu_2455_p2 = (sub_ln703_316_fu_2421_p2 - data_19_V_read_7_reg_4567_pp0_iter6_reg);

assign sub_ln703_331_fu_2258_p2 = (add_ln703_366_fu_2193_p2 - data_19_V_read_7_reg_4567_pp0_iter5_reg);

assign sub_ln703_332_fu_2273_p2 = (add_ln703_367_fu_2198_p2 - data_19_V_read_7_reg_4567_pp0_iter5_reg);

assign sub_ln703_333_fu_2460_p2 = (sub_ln703_318_reg_5783 - data_19_V_read_7_reg_4567_pp0_iter6_reg);

assign sub_ln703_334_fu_2464_p2 = (add_ln703_368_fu_2429_p2 - data_19_V_read_7_reg_4567_pp0_iter6_reg);

assign sub_ln703_335_fu_2302_p2 = (add_ln703_369_fu_2213_p2 - data_20_V_read21_reg_4539_pp0_iter5_reg);

assign sub_ln703_336_fu_2469_p2 = (sub_ln703_321_reg_5788 - data_20_V_read21_reg_4539_pp0_iter6_reg);

assign sub_ln703_337_fu_2473_p2 = (add_ln703_370_fu_2437_p2 - data_20_V_read21_reg_4539_pp0_iter6_reg);

assign sub_ln703_338_fu_2478_p2 = (add_ln703_372_reg_5793 - data_20_V_read21_reg_4539_pp0_iter6_reg);

assign sub_ln703_339_fu_2482_p2 = (sub_ln703_324_reg_5803 - data_20_V_read21_reg_4539_pp0_iter6_reg);

assign sub_ln703_340_fu_2495_p2 = (sub_ln703_327_reg_5813 - data_20_V_read21_reg_4539_pp0_iter6_reg);

assign sub_ln703_341_fu_2504_p2 = (add_ln703_373_fu_2445_p2 - data_20_V_read21_reg_4539_pp0_iter6_reg);

assign sub_ln703_342_fu_2509_p2 = (sub_ln703_329_fu_2450_p2 - data_20_V_read21_reg_4539_pp0_iter6_reg);

assign sub_ln703_343_fu_2312_p2 = (add_ln703_375_fu_2268_p2 - data_20_V_read21_reg_4539_pp0_iter5_reg);

assign sub_ln703_344_fu_2523_p2 = (add_ln703_377_reg_5833 - data_20_V_read21_reg_4539_pp0_iter6_reg);

assign sub_ln703_345_fu_2532_p2 = (add_ln703_379_reg_5838 - data_20_V_read21_reg_4539_pp0_iter6_reg);

assign sub_ln703_346_fu_2332_p2 = (add_ln703_380_fu_2297_p2 - data_20_V_read21_reg_4539_pp0_iter5_reg);

assign sub_ln703_347_fu_2536_p2 = (sub_ln703_335_reg_5843 - data_21_V_read22_reg_4512_pp0_iter6_reg);

assign sub_ln703_348_fu_2545_p2 = (add_ln703_381_reg_5848 - data_21_V_read22_reg_4512_pp0_iter6_reg);

assign sub_ln703_349_fu_2549_p2 = (sub_ln703_337_fu_2473_p2 - data_21_V_read22_reg_4512_pp0_iter6_reg);

assign sub_ln703_350_fu_2554_p2 = (sub_ln703_338_fu_2478_p2 - data_21_V_read22_reg_4512_pp0_iter6_reg);

assign sub_ln703_351_fu_2574_p2 = (sub_ln703_339_fu_2482_p2 - data_21_V_read22_reg_4512_pp0_iter6_reg);

assign sub_ln703_352_fu_2579_p2 = (add_ln703_382_fu_2486_p2 - data_21_V_read22_reg_4512_pp0_iter6_reg);

assign sub_ln703_353_fu_2584_p2 = (add_ln703_383_fu_2490_p2 - data_21_V_read22_reg_4512_pp0_iter6_reg);

assign sub_ln703_354_fu_2589_p2 = (sub_ln703_340_fu_2495_p2 - data_21_V_read22_reg_4512_pp0_iter6_reg);

assign sub_ln703_355_fu_2594_p2 = (add_ln703_385_fu_2499_p2 - data_21_V_read22_reg_4512_pp0_iter6_reg);

assign sub_ln703_356_fu_2603_p2 = (sub_ln703_341_fu_2504_p2 - data_21_V_read22_reg_4512_pp0_iter6_reg);

assign sub_ln703_357_fu_2608_p2 = (sub_ln703_342_fu_2509_p2 - data_21_V_read22_reg_4512_pp0_iter6_reg);

assign sub_ln703_358_fu_2613_p2 = (add_ln703_386_fu_2514_p2 - data_21_V_read22_reg_4512_pp0_iter6_reg);

assign sub_ln703_359_fu_2618_p2 = (add_ln703_387_fu_2518_p2 - data_21_V_read22_reg_4512_pp0_iter6_reg);

assign sub_ln703_360_fu_2627_p2 = (add_ln703_390_reg_5858 - data_21_V_read22_reg_4512_pp0_iter6_reg);

assign sub_ln703_361_fu_2636_p2 = (add_ln703_391_fu_2527_p2 - data_21_V_read22_reg_4512_pp0_iter6_reg);

assign sub_ln703_362_fu_2641_p2 = (sub_ln703_346_reg_5863 - data_21_V_read22_reg_4512_pp0_iter6_reg);

assign sub_ln703_363_fu_2660_p2 = (add_ln703_392_fu_2540_p2 - data_22_V_read23_reg_4483_pp0_iter6_reg);

assign sub_ln703_364_fu_2665_p2 = (sub_ln703_348_fu_2545_p2 - data_22_V_read23_reg_4483_pp0_iter6_reg);

assign sub_ln703_365_fu_2670_p2 = (sub_ln703_350_fu_2554_p2 - data_22_V_read23_reg_4483_pp0_iter6_reg);

assign sub_ln703_366_fu_2684_p2 = (add_ln703_396_fu_2568_p2 - data_22_V_read23_reg_4483_pp0_iter6_reg);

assign sub_ln703_367_fu_2689_p2 = (sub_ln703_351_fu_2574_p2 - data_22_V_read23_reg_4483_pp0_iter6_reg);

assign sub_ln703_368_fu_2694_p2 = (sub_ln703_352_fu_2579_p2 - data_22_V_read23_reg_4483_pp0_iter6_reg);

assign sub_ln703_369_fu_2699_p2 = (sub_ln703_353_fu_2584_p2 - data_22_V_read23_reg_4483_pp0_iter6_reg);

assign sub_ln703_370_fu_2714_p2 = (add_ln703_397_fu_2599_p2 - data_22_V_read23_reg_4483_pp0_iter6_reg);

assign sub_ln703_371_fu_2719_p2 = (add_ln703_400_reg_5868 - data_22_V_read23_reg_4483_pp0_iter6_reg);

assign sub_ln703_372_fu_2985_p2 = (sub_ln703_356_reg_5921 - data_22_V_read23_reg_4483_pp0_iter7_reg);

assign sub_ln703_373_fu_2723_p2 = (sub_ln703_358_fu_2613_p2 - data_22_V_read23_reg_4483_pp0_iter6_reg);

assign sub_ln703_374_fu_2728_p2 = (sub_ln703_359_fu_2618_p2 - data_22_V_read23_reg_4483_pp0_iter6_reg);

assign sub_ln703_375_fu_2747_p2 = (add_ln703_401_fu_2623_p2 - data_22_V_read23_reg_4483_pp0_iter6_reg);

assign sub_ln703_376_fu_2752_p2 = (sub_ln703_360_fu_2627_p2 - data_22_V_read23_reg_4483_pp0_iter6_reg);

assign sub_ln703_377_fu_2989_p2 = (add_ln703_402_reg_5931 - data_22_V_read23_reg_4483_pp0_iter7_reg);

assign sub_ln703_378_fu_2776_p2 = (sub_ln703_362_fu_2641_p2 - data_22_V_read23_reg_4483_pp0_iter6_reg);

assign sub_ln703_379_fu_2781_p2 = (add_ln703_405_fu_2650_p2 - data_23_V_read24_reg_4451_pp0_iter6_reg);

assign sub_ln703_380_fu_2786_p2 = (add_ln703_406_fu_2655_p2 - data_23_V_read24_reg_4451_pp0_iter6_reg);

assign sub_ln703_381_fu_2791_p2 = (sub_ln703_363_fu_2660_p2 - data_23_V_read24_reg_4451_pp0_iter6_reg);

assign sub_ln703_382_fu_2796_p2 = (sub_ln703_364_fu_2665_p2 - data_23_V_read24_reg_4451_pp0_iter6_reg);

assign sub_ln703_383_fu_2801_p2 = (add_ln703_408_fu_2679_p2 - data_23_V_read24_reg_4451_pp0_iter6_reg);

assign sub_ln703_384_fu_2997_p2 = (sub_ln703_366_reg_5941 - data_23_V_read24_reg_4451_pp0_iter7_reg);

assign sub_ln703_385_fu_2811_p2 = (sub_ln703_368_fu_2694_p2 - data_23_V_read24_reg_4451_pp0_iter6_reg);

assign sub_ln703_386_fu_2816_p2 = (add_ln703_409_fu_2704_p2 - data_23_V_read24_reg_4451_pp0_iter6_reg);

assign sub_ln703_387_fu_3005_p2 = (add_ln703_410_reg_5951 - data_23_V_read24_reg_4451_pp0_iter7_reg);

assign sub_ln703_388_fu_2821_p2 = (add_ln703_413_reg_5873 - data_23_V_read24_reg_4451_pp0_iter6_reg);

assign sub_ln703_389_fu_2839_p2 = (sub_ln703_371_fu_2719_p2 - data_23_V_read24_reg_4451_pp0_iter6_reg);

assign sub_ln703_390_fu_3009_p2 = (sub_ln703_372_fu_2985_p2 - data_23_V_read24_reg_4451_pp0_iter7_reg);

assign sub_ln703_391_fu_2844_p2 = (add_ln703_415_reg_5878 - data_23_V_read24_reg_4451_pp0_iter6_reg);

assign sub_ln703_392_fu_2848_p2 = (sub_ln703_373_fu_2723_p2 - data_23_V_read24_reg_4451_pp0_iter6_reg);

assign sub_ln703_393_fu_3018_p2 = (add_ln703_418_reg_5961 - data_23_V_read24_reg_4451_pp0_iter7_reg);

assign sub_ln703_394_fu_3022_p2 = (sub_ln703_375_reg_5966 - data_23_V_read24_reg_4451_pp0_iter7_reg);

assign sub_ln703_395_fu_2853_p2 = (sub_ln703_376_fu_2752_p2 - data_23_V_read24_reg_4451_pp0_iter6_reg);

assign sub_ln703_396_fu_2858_p2 = (add_ln703_420_fu_2761_p2 - data_23_V_read24_reg_4451_pp0_iter6_reg);

assign sub_ln703_397_fu_2863_p2 = (add_ln703_422_fu_2771_p2 - data_23_V_read24_reg_4451_pp0_iter6_reg);

assign sub_ln703_398_fu_3026_p2 = (sub_ln703_377_fu_2989_p2 - data_23_V_read24_reg_4451_pp0_iter7_reg);

assign sub_ln703_399_fu_3031_p2 = (add_ln703_423_fu_2993_p2 - data_23_V_read24_reg_4451_pp0_iter7_reg);

assign sub_ln703_400_fu_2868_p2 = (sub_ln703_378_fu_2776_p2 - data_23_V_read24_reg_4451_pp0_iter6_reg);

assign sub_ln703_401_fu_3040_p2 = (sub_ln703_381_reg_5976 - data_24_V_read25_reg_4421_pp0_iter7_reg);

assign sub_ln703_402_fu_2878_p2 = (sub_ln703_382_fu_2796_p2 - data_24_V_read25_reg_4421_pp0_iter6_reg);

assign sub_ln703_403_fu_3044_p2 = (sub_ln703_384_fu_2997_p2 - data_24_V_read25_reg_4421_pp0_iter7_reg);

assign sub_ln703_404_fu_3049_p2 = (add_ln703_424_reg_5981 - data_24_V_read25_reg_4421_pp0_iter7_reg);

assign sub_ln703_405_fu_3057_p2 = (add_ln703_425_fu_3001_p2 - data_24_V_read25_reg_4421_pp0_iter7_reg);

assign sub_ln703_406_fu_3062_p2 = (sub_ln703_386_reg_5991 - data_24_V_read25_reg_4421_pp0_iter7_reg);

assign sub_ln703_407_fu_3066_p2 = (sub_ln703_387_fu_3005_p2 - data_24_V_read25_reg_4421_pp0_iter7_reg);

assign sub_ln703_408_fu_2893_p2 = (sub_ln703_388_fu_2821_p2 - data_24_V_read25_reg_4421_pp0_iter6_reg);

assign sub_ln703_409_fu_2898_p2 = (add_ln703_431_fu_2834_p2 - data_24_V_read25_reg_4421_pp0_iter6_reg);

assign sub_ln703_410_fu_3071_p2 = (sub_ln703_389_reg_5996 - data_24_V_read25_reg_4421_pp0_iter7_reg);

assign sub_ln703_411_fu_2903_p2 = (sub_ln703_391_fu_2844_p2 - data_24_V_read25_reg_4421_pp0_iter6_reg);

assign sub_ln703_412_fu_3080_p2 = (sub_ln703_392_reg_6001 - data_24_V_read25_reg_4421_pp0_iter7_reg);

assign sub_ln703_413_fu_3084_p2 = (add_ln703_432_fu_3014_p2 - data_24_V_read25_reg_4421_pp0_iter7_reg);

assign sub_ln703_414_fu_3089_p2 = (sub_ln703_393_fu_3018_p2 - data_24_V_read25_reg_4421_pp0_iter7_reg);

assign sub_ln703_415_fu_3094_p2 = (sub_ln703_394_fu_3022_p2 - data_24_V_read25_reg_4421_pp0_iter7_reg);

assign sub_ln703_416_fu_2923_p2 = (sub_ln703_396_fu_2858_p2 - data_24_V_read25_reg_4421_pp0_iter6_reg);

assign sub_ln703_417_fu_3103_p2 = (sub_ln703_399_fu_3031_p2 - data_24_V_read25_reg_4421_pp0_iter7_reg);

assign sub_ln703_418_fu_3108_p2 = (add_ln703_433_fu_3036_p2 - data_25_V_read26_reg_4391_pp0_iter7_reg);

assign sub_ln703_419_fu_3113_p2 = (add_ln703_434_reg_6011 - data_25_V_read26_reg_4391_pp0_iter7_reg);

assign sub_ln703_420_fu_3117_p2 = (sub_ln703_401_fu_3040_p2 - data_25_V_read26_reg_4391_pp0_iter7_reg);

assign sub_ln703_421_fu_3126_p2 = (add_ln703_436_reg_6021 - data_25_V_read26_reg_4391_pp0_iter7_reg);

assign sub_ln703_422_fu_3130_p2 = (sub_ln703_403_fu_3044_p2 - data_25_V_read26_reg_4391_pp0_iter7_reg);

assign sub_ln703_423_fu_3135_p2 = (sub_ln703_404_fu_3049_p2 - data_25_V_read26_reg_4391_pp0_iter7_reg);

assign sub_ln703_424_fu_3140_p2 = (add_ln703_437_fu_3053_p2 - data_25_V_read26_reg_4391_pp0_iter7_reg);

assign sub_ln703_425_fu_3145_p2 = (sub_ln703_406_fu_3062_p2 - data_25_V_read26_reg_4391_pp0_iter7_reg);

assign sub_ln703_426_fu_2938_p2 = (add_ln703_438_fu_2888_p2 - data_25_V_read26_reg_4391_pp0_iter6_reg);

assign sub_ln703_427_fu_3154_p2 = (sub_ln703_409_reg_6031 - data_25_V_read26_reg_4391_pp0_iter7_reg);

assign sub_ln703_428_fu_3163_p2 = (add_ln703_439_fu_3075_p2 - data_25_V_read26_reg_4391_pp0_iter7_reg);

assign sub_ln703_429_fu_3177_p2 = (sub_ln703_411_reg_6036 - data_25_V_read26_reg_4391_pp0_iter7_reg);

assign sub_ln703_430_fu_3181_p2 = (add_ln703_442_reg_6041 - data_25_V_read26_reg_4391_pp0_iter7_reg);

assign sub_ln703_431_fu_3185_p2 = (sub_ln703_412_fu_3080_p2 - data_25_V_read26_reg_4391_pp0_iter7_reg);

assign sub_ln703_432_fu_3190_p2 = (sub_ln703_416_reg_6046 - data_25_V_read26_reg_4391_pp0_iter7_reg);

assign sub_ln703_433_fu_3194_p2 = (add_ln703_443_fu_3099_p2 - data_25_V_read26_reg_4391_pp0_iter7_reg);

assign sub_ln703_434_fu_3199_p2 = (sub_ln703_417_fu_3103_p2 - data_25_V_read26_reg_4391_pp0_iter7_reg);

assign sub_ln703_435_fu_3204_p2 = (add_ln703_444_reg_6051 - data_25_V_read26_reg_4391_pp0_iter7_reg);

assign sub_ln703_436_fu_3208_p2 = (sub_ln703_418_fu_3108_p2 - data_26_V_read27_reg_4365_pp0_iter7_reg);

assign sub_ln703_437_fu_3213_p2 = (sub_ln703_419_fu_3113_p2 - data_26_V_read27_reg_4365_pp0_iter7_reg);

assign sub_ln703_438_fu_3223_p2 = (add_ln703_445_fu_3122_p2 - data_26_V_read27_reg_4365_pp0_iter7_reg);

assign sub_ln703_439_fu_3228_p2 = (add_ln703_447_reg_6056 - data_26_V_read27_reg_4365_pp0_iter7_reg);

assign sub_ln703_440_fu_3247_p2 = (sub_ln703_425_fu_3145_p2 - data_26_V_read27_reg_4365_pp0_iter7_reg);

assign sub_ln703_441_fu_3252_p2 = (sub_ln703_426_reg_6061 - data_26_V_read27_reg_4365_pp0_iter7_reg);

assign sub_ln703_442_fu_3256_p2 = (add_ln703_448_fu_3150_p2 - data_26_V_read27_reg_4365_pp0_iter7_reg);

assign sub_ln703_443_fu_3261_p2 = (sub_ln703_427_fu_3154_p2 - data_26_V_read27_reg_4365_pp0_iter7_reg);

assign sub_ln703_444_fu_3266_p2 = (add_ln703_449_fu_3158_p2 - data_26_V_read27_reg_4365_pp0_iter7_reg);

assign sub_ln703_445_fu_3271_p2 = (add_ln703_452_fu_3172_p2 - data_26_V_read27_reg_4365_pp0_iter7_reg);

assign sub_ln703_446_fu_3276_p2 = (sub_ln703_429_fu_3177_p2 - data_26_V_read27_reg_4365_pp0_iter7_reg);

assign sub_ln703_447_fu_3298_p2 = (sub_ln703_432_fu_3190_p2 - data_26_V_read27_reg_4365_pp0_iter7_reg);

assign sub_ln703_448_fu_3308_p2 = (sub_ln703_436_fu_3208_p2 - data_27_V_read_8_reg_4342_pp0_iter7_reg);

assign sub_ln703_449_fu_3313_p2 = (sub_ln703_437_fu_3213_p2 - data_27_V_read_8_reg_4342_pp0_iter7_reg);

assign sub_ln703_450_fu_3318_p2 = (add_ln703_453_fu_3218_p2 - data_27_V_read_8_reg_4342_pp0_iter7_reg);

assign sub_ln703_451_fu_3343_p2 = (add_ln703_454_fu_3232_p2 - data_27_V_read_8_reg_4342_pp0_iter7_reg);

assign sub_ln703_452_fu_3348_p2 = (add_ln703_456_fu_3241_p2 - data_27_V_read_8_reg_4342_pp0_iter7_reg);

assign sub_ln703_453_fu_3353_p2 = (sub_ln703_440_fu_3247_p2 - data_27_V_read_8_reg_4342_pp0_iter7_reg);

assign sub_ln703_454_fu_3368_p2 = (sub_ln703_441_fu_3252_p2 - data_27_V_read_8_reg_4342_pp0_iter7_reg);

assign sub_ln703_455_fu_3373_p2 = (sub_ln703_444_fu_3266_p2 - data_27_V_read_8_reg_4342_pp0_iter7_reg);

assign sub_ln703_456_fu_3388_p2 = (add_ln703_457_fu_3281_p2 - data_27_V_read_8_reg_4342_pp0_iter7_reg);

assign sub_ln703_457_fu_3393_p2 = (add_ln703_458_fu_3286_p2 - data_27_V_read_8_reg_4342_pp0_iter7_reg);

assign sub_ln703_458_fu_3408_p2 = (add_ln703_459_fu_3292_p2 - data_27_V_read_8_reg_4342_pp0_iter7_reg);

assign sub_ln703_459_fu_3418_p2 = (add_ln703_460_fu_3303_p2 - data_27_V_read_8_reg_4342_pp0_iter7_reg);

assign sub_ln703_460_fu_3535_p2 = (sub_ln703_450_reg_6123 - data_28_V_read_7_reg_4313_pp0_iter8_reg);

assign sub_ln703_461_fu_3438_p2 = (add_ln703_461_fu_3323_p2 - data_28_V_read_7_reg_4313_pp0_iter7_reg);

assign sub_ln703_462_fu_3539_p2 = (add_ln703_463_reg_6128 - data_28_V_read_7_reg_4313_pp0_iter8_reg);

assign sub_ln703_463_fu_3543_p2 = (add_ln703_464_reg_6133 - data_28_V_read_7_reg_4313_pp0_iter8_reg);

assign sub_ln703_464_fu_3547_p2 = (add_ln703_465_reg_6138 - data_28_V_read_7_reg_4313_pp0_iter8_reg);

assign sub_ln703_465_fu_3551_p2 = (sub_ln703_451_reg_6143 - data_28_V_read_7_reg_4313_pp0_iter8_reg);

assign sub_ln703_466_fu_3563_p2 = (add_ln703_467_reg_6158 - data_28_V_read_7_reg_4313_pp0_iter8_reg);

assign sub_ln703_467_fu_3567_p2 = (sub_ln703_454_reg_6163 - data_28_V_read_7_reg_4313_pp0_iter8_reg);

assign sub_ln703_468_fu_3575_p2 = (add_ln703_468_reg_6173 - data_28_V_read_7_reg_4313_pp0_iter8_reg);

assign sub_ln703_469_fu_3463_p2 = (add_ln703_469_fu_3383_p2 - data_28_V_read_7_reg_4313_pp0_iter7_reg);

assign sub_ln703_470_fu_3579_p2 = (sub_ln703_456_reg_6178 - data_28_V_read_7_reg_4313_pp0_iter8_reg);

assign sub_ln703_471_fu_3583_p2 = (sub_ln703_457_reg_6183 - data_28_V_read_7_reg_4313_pp0_iter8_reg);

assign sub_ln703_472_fu_3587_p2 = (add_ln703_471_reg_6188 - data_28_V_read_7_reg_4313_pp0_iter8_reg);

assign sub_ln703_473_fu_3591_p2 = (sub_ln703_458_reg_6193 - data_28_V_read_7_reg_4313_pp0_iter8_reg);

assign sub_ln703_474_fu_3482_p2 = (add_ln703_472_fu_3413_p2 - data_28_V_read_7_reg_4313_pp0_iter7_reg);

assign sub_ln703_475_fu_3599_p2 = (sub_ln703_459_reg_6198 - data_28_V_read_7_reg_4313_pp0_iter8_reg);

assign sub_ln703_476_fu_3603_p2 = (add_ln703_475_reg_6203 - data_28_V_read_7_reg_4313_pp0_iter8_reg);

assign sub_ln703_477_fu_3607_p2 = (add_ln703_476_fu_3531_p2 - data_28_V_read_7_reg_4313_pp0_iter8_reg);

assign sub_ln703_478_fu_3612_p2 = (add_ln703_480_reg_6072_pp0_iter8_reg - data_28_V_read_7_reg_4313_pp0_iter8_reg);

assign sub_ln703_479_fu_3621_p2 = (sub_ln703_462_fu_3539_p2 - data_29_V_read_7_reg_4279_pp0_iter8_reg);

assign sub_ln703_480_fu_3626_p2 = (sub_ln703_463_fu_3543_p2 - data_29_V_read_7_reg_4279_pp0_iter8_reg);

assign sub_ln703_481_fu_3636_p2 = (add_ln703_483_reg_6213 - data_29_V_read_7_reg_4279_pp0_iter8_reg);

assign sub_ln703_482_fu_3640_p2 = (sub_ln703_465_fu_3551_p2 - data_29_V_read_7_reg_4279_pp0_iter8_reg);

assign sub_ln703_483_fu_3645_p2 = (add_ln703_484_fu_3555_p2 - data_29_V_read_7_reg_4279_pp0_iter8_reg);

assign sub_ln703_484_fu_3650_p2 = (add_ln703_485_fu_3559_p2 - data_29_V_read_7_reg_4279_pp0_iter8_reg);

assign sub_ln703_485_fu_3660_p2 = (sub_ln703_467_fu_3567_p2 - data_29_V_read_7_reg_4279_pp0_iter8_reg);

assign sub_ln703_486_fu_3507_p2 = (add_ln703_486_fu_3453_p2 - data_29_V_read_7_reg_4279_pp0_iter7_reg);

assign sub_ln703_487_fu_3512_p2 = (add_ln703_487_fu_3458_p2 - data_29_V_read_7_reg_4279_pp0_iter7_reg);

assign sub_ln703_488_fu_3665_p2 = (add_ln703_488_fu_3571_p2 - data_29_V_read_7_reg_4279_pp0_iter8_reg);

assign sub_ln703_489_fu_3670_p2 = (sub_ln703_468_fu_3575_p2 - data_29_V_read_7_reg_4279_pp0_iter8_reg);

assign sub_ln703_490_fu_3675_p2 = (sub_ln703_469_reg_6218 - data_29_V_read_7_reg_4279_pp0_iter8_reg);

assign sub_ln703_491_fu_3517_p2 = (add_ln703_490_fu_3473_p2 - data_29_V_read_7_reg_4279_pp0_iter7_reg);

assign sub_ln703_492_fu_3679_p2 = (sub_ln703_470_fu_3579_p2 - data_29_V_read_7_reg_4279_pp0_iter8_reg);

assign sub_ln703_493_fu_3684_p2 = (sub_ln703_471_fu_3583_p2 - data_29_V_read_7_reg_4279_pp0_iter8_reg);

assign sub_ln703_494_fu_3689_p2 = (sub_ln703_472_fu_3587_p2 - data_29_V_read_7_reg_4279_pp0_iter8_reg);

assign sub_ln703_495_fu_3694_p2 = (sub_ln703_473_fu_3591_p2 - data_29_V_read_7_reg_4279_pp0_iter8_reg);

assign sub_ln703_496_fu_3699_p2 = (add_ln703_493_fu_3595_p2 - data_29_V_read_7_reg_4279_pp0_iter8_reg);

assign sub_ln703_497_fu_3704_p2 = (sub_ln703_474_reg_6229 - data_29_V_read_7_reg_4279_pp0_iter8_reg);

assign sub_ln703_498_fu_3718_p2 = (sub_ln703_477_fu_3607_p2 - data_29_V_read_7_reg_4279_pp0_iter8_reg);

assign sub_ln703_499_fu_3723_p2 = (sub_ln703_478_fu_3612_p2 - data_29_V_read_7_reg_4279_pp0_iter8_reg);

assign sub_ln703_500_fu_3522_p2 = (add_ln703_495_fu_3492_p2 - data_29_V_read_7_reg_4279_pp0_iter7_reg);

assign sub_ln703_501_fu_3728_p2 = (add_ln703_497_reg_6239 - data_30_V_read31_reg_4250_pp0_iter8_reg);

assign sub_ln703_502_fu_3732_p2 = (add_ln703_498_fu_3616_p2 - data_30_V_read31_reg_4250_pp0_iter8_reg);

assign sub_ln703_503_fu_3737_p2 = (sub_ln703_479_fu_3621_p2 - data_30_V_read31_reg_4250_pp0_iter8_reg);

assign sub_ln703_504_fu_3742_p2 = (sub_ln703_480_fu_3626_p2 - data_30_V_read31_reg_4250_pp0_iter8_reg);

assign sub_ln703_505_fu_3747_p2 = (add_ln703_499_fu_3631_p2 - data_30_V_read31_reg_4250_pp0_iter8_reg);

assign sub_ln703_506_fu_3752_p2 = (sub_ln703_482_fu_3640_p2 - data_30_V_read31_reg_4250_pp0_iter8_reg);

assign sub_ln703_507_fu_3762_p2 = (sub_ln703_484_fu_3650_p2 - data_30_V_read31_reg_4250_pp0_iter8_reg);

assign sub_ln703_508_fu_3767_p2 = (add_ln703_500_fu_3655_p2 - data_30_V_read31_reg_4250_pp0_iter8_reg);

assign sub_ln703_509_fu_3772_p2 = (sub_ln703_485_fu_3660_p2 - data_30_V_read31_reg_4250_pp0_iter8_reg);

assign sub_ln703_510_fu_3781_p2 = (sub_ln703_487_reg_6249 - data_30_V_read31_reg_4250_pp0_iter8_reg);

assign sub_ln703_511_fu_3790_p2 = (sub_ln703_489_fu_3670_p2 - data_30_V_read31_reg_4250_pp0_iter8_reg);

assign sub_ln703_512_fu_3804_p2 = (sub_ln703_493_fu_3684_p2 - data_30_V_read31_reg_4250_pp0_iter8_reg);

assign sub_ln703_513_fu_3809_p2 = (sub_ln703_494_fu_3689_p2 - data_30_V_read31_reg_4250_pp0_iter8_reg);

assign sub_ln703_514_fu_3814_p2 = (sub_ln703_495_fu_3694_p2 - data_30_V_read31_reg_4250_pp0_iter8_reg);

assign sub_ln703_515_fu_3819_p2 = (sub_ln703_496_fu_3699_p2 - data_30_V_read31_reg_4250_pp0_iter8_reg);

assign sub_ln703_516_fu_3824_p2 = (add_ln703_501_fu_3708_p2 - data_30_V_read31_reg_4250_pp0_iter8_reg);

assign sub_ln703_517_fu_3829_p2 = (add_ln703_502_fu_3713_p2 - data_30_V_read31_reg_4250_pp0_iter8_reg);

assign sub_ln703_518_fu_3834_p2 = (sub_ln703_499_fu_3723_p2 - data_30_V_read31_reg_4250_pp0_iter8_reg);

assign sub_ln703_519_fu_3839_p2 = (sub_ln703_500_reg_6259 - data_30_V_read31_reg_4250_pp0_iter8_reg);

assign sub_ln703_73_fu_286_p2 = (data_0_V_read_int_reg - data_1_V_read_int_reg);

assign sub_ln703_74_fu_292_p2 = (sub_ln703_reg_5046 - data_2_V_read_9_reg_5035);

assign sub_ln703_75_fu_296_p2 = (add_ln703_reg_5052 - data_2_V_read_9_reg_5035);

assign sub_ln703_76_fu_300_p2 = (sub_ln703_73_reg_5059 - data_2_V_read_9_reg_5035);

assign sub_ln703_77_fu_308_p2 = (data_2_V_read_9_reg_5035 - add_ln703_reg_5052);

assign sub_ln703_78_fu_361_p2 = (sub_ln703_76_reg_5071_pp0_iter2_reg - data_3_V_read_9_reg_5019_pp0_iter2_reg);

assign sub_ln703_79_fu_337_p2 = (sub_ln703_77_reg_5084 - data_3_V_read_9_reg_5019_pp0_iter1_reg);

assign sub_ln703_80_fu_365_p2 = (add_ln703_201_reg_5090_pp0_iter2_reg - data_3_V_read_9_reg_5019_pp0_iter2_reg);

assign sub_ln703_81_fu_369_p2 = (add_ln703_202_reg_5096_pp0_iter2_reg - data_3_V_read_9_reg_5019_pp0_iter2_reg);

assign sub_ln703_82_fu_373_p2 = (data_3_V_read_9_reg_5019_pp0_iter2_reg - add_ln703_200_reg_5077_pp0_iter2_reg);

assign sub_ln703_83_fu_377_p2 = (add_ln703_200_reg_5077_pp0_iter2_reg - data_3_V_read_9_reg_5019_pp0_iter2_reg);

assign sub_ln703_84_fu_381_p2 = (sub_ln703_74_reg_5065_pp0_iter2_reg - data_3_V_read_9_reg_5019_pp0_iter2_reg);

assign sub_ln703_85_fu_385_p2 = (add_ln703_203_reg_5113 - data_4_V_read_9_reg_4998_pp0_iter2_reg);

assign sub_ln703_86_fu_389_p2 = (add_ln703_204_reg_5101_pp0_iter2_reg - data_4_V_read_9_reg_4998_pp0_iter2_reg);

assign sub_ln703_87_fu_393_p2 = (sub_ln703_78_fu_361_p2 - data_4_V_read_9_reg_4998_pp0_iter2_reg);

assign sub_ln703_88_fu_398_p2 = (data_4_V_read_9_reg_4998_pp0_iter2_reg - add_ln703_205_reg_5119);

assign sub_ln703_89_fu_402_p2 = (sub_ln703_79_reg_5125 - data_4_V_read_9_reg_4998_pp0_iter2_reg);

assign sub_ln703_90_fu_406_p2 = (sub_ln703_80_fu_365_p2 - data_4_V_read_9_reg_4998_pp0_iter2_reg);

assign sub_ln703_91_fu_411_p2 = (sub_ln703_81_fu_369_p2 - data_4_V_read_9_reg_4998_pp0_iter2_reg);

assign sub_ln703_92_fu_437_p2 = (sub_ln703_84_fu_381_p2 - data_4_V_read_9_reg_4998_pp0_iter2_reg);

assign sub_ln703_93_fu_442_p2 = (add_ln703_206_reg_5131 - data_4_V_read_9_reg_4998_pp0_iter2_reg);

assign sub_ln703_94_fu_446_p2 = (sub_ln703_86_fu_389_p2 - data_5_V_read_8_reg_4969_pp0_iter2_reg);

assign sub_ln703_95_fu_451_p2 = (sub_ln703_87_fu_393_p2 - data_5_V_read_8_reg_4969_pp0_iter2_reg);

assign sub_ln703_96_fu_456_p2 = (sub_ln703_88_fu_398_p2 - data_5_V_read_8_reg_4969_pp0_iter2_reg);

assign sub_ln703_97_fu_609_p2 = (sub_ln703_91_reg_5172 - data_5_V_read_8_reg_4969_pp0_iter3_reg);

assign sub_ln703_98_fu_466_p2 = (add_ln703_208_reg_5137 - data_5_V_read_8_reg_4969_pp0_iter2_reg);

assign sub_ln703_99_fu_613_p2 = (data_5_V_read_8_reg_4969_pp0_iter3_reg - add_ln703_209_reg_5178);

assign sub_ln703_fu_274_p2 = (data_1_V_read_int_reg - data_0_V_read_int_reg);

endmodule //dense_latency_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_0_2
